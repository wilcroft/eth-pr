// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:35:04 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
m8E0QLr+EPq6eNpFfaWFC0GdBC0pHK232QtwoZonQPBC/IESlARfm8XsZcLfKjmf
pFy41rXZj4kr3QtaV2j4mBz2M1V18obwZgT6wvSVCNoDlDhX1DlpXSZh0UKBP4uR
ktEc+vlXKA2U/f7gnAdhh7bObzkqd5OG5ULsjdYWax0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5568)
3WykMyKIvWpc+HmJlfGCtFA+pj/lpnCL2YZtMVzXyrlY7s7hpULveWPSPaSDb5v1
hvhE1Ur9rVVXaQZcSh1h3vinO+LipgDX5u23V65dim8D1d1d2K9rKM8qZtRczuy5
QIVSpRO0FXHXIE0TUyMept5Gdl8H+v7UCF+5CxqYFx51rQHs4FGG6ba5u8sKSk3k
4Xys23NlNvdCmBK/HwRLSCJXVKmFfZF++KegLhvj+9+g+Kg09SlzBzjLZS9lDGiC
yvKXCLtjhaQSGnD36PutzxidtFRMS0oeOtr15k8P87MMilVS5Y52FFwfG5BVCHc1
1gaHIHEM3CLhah/einbK5itTL4FSnNk3DYuJq+HyPBPWJJoLdnXayh2pKXCHylAN
8CBxs/wt33JxF8CIHaMoq38/v6atahemQ+OIMGXySw1wVS1MrZfGNSDIwlhHFzAd
IRUsD3HvuCeXUEIVkRq5Rfvk+3YPXInxzeQkN/RI+IywTjIicT2vZRuBbkAyjvaV
ZKiGunN/7k1I9ODJBaQ3PoJyKGN3ZWYqi1loi0w2HPIxQMyP5Ody3ZSMiGtF6uDb
VvsgM+ymbgbnbHopy9lR4Tl9XATLeawz4Am2ElIH7MmzuyWAreW1sxDQPT5h64M7
ekM2z9+yTEJILrpcBXvOSVecs1g1bL9E4Q+obexa45pPtMxA37GFmJ3rEg4fWL1D
B6ikJJM9J4HTqvDwLMegLRB3CircMTcrHNgp2U+3C2w97VnPqmNbdM974u3quIBU
TE5nJp7sbCN8Kihsop0PvkKQA3aZzXNzh81fn8I3fO6bJDs0Q/CtDKjX5fNcWOBs
0JyCJ6twTRdBtLA8kU0nIQfy+Z7hklkC1SmzitT83AXZ1zQiykL+rg4GUde4nq92
sXKUUujwlmRE5hZQKrZzHEaakdG2wMMe8sSgCHfHFjq13hWKIsV2PnSAnlS8Lr0r
/iDe8yi9AlneOXuTDX6hZhDEDBJNsx1WVcMI5nWOs2s3dUHw2+KpL724w/6Y9zeh
0rVsNBAdrrc6TMj+e54LfvkB1JxrVN+pFcbSv2Kc9xemYe1/5oWjAwpfZX/Tgol+
9p7qcxnJjKHP/fK94p8BY00Msjzd07aHQPxl+Eno2lO26co4U5wIDTdHlWqXUvUr
FJwSMfh7jPb9JBIsEiaPeWG0tI+BL1yWAybFLgptoHre4gp9h98ca59h5FdBGR2o
pNxZMyuEH+xyDw478vEkxApV4LaDBZPkKndqCr98c12dkdxjL4qnbzC57eWw9pjg
BBwnF143y6ptj/LKRAbmswbN6lGCGd7DfTrX9C5P13ql0W/EeZAFXzsCQF6+2thW
jOpyiEHld/4SJDRTnZ4fSC2T5OvYoYzMsIu/H31GtJwxaLFS5K9P/G87hDhXxE3L
ZkJdpELP+QwRVkpcWZAaNlwvmFyNPE8nyGvnSkFUBLBMxxWGarRvBgAz3TVc+4Gl
80K7p6tajyxkvluPUSn5gAeR5omBgC/UqBUhOFaPUS+QRt19+krmgt5AQyfDT1S/
awP4dsqYvtbyY6yE1EE/OyP+Zs+xitgVkUDn8hW8tgkLsGRrmYY6vR+hbIx8kwPi
aKztfKy7uJ65wQP2BpIT7dwWkkAIj7nYGgBqqyV6wDj4/cpYO5T5EziDkiJEvMGF
HAfBBlXhSGCn98x9UdJ0cp2fAANLMyGJ+VN89y6wnqDltOQPTXEVJEeTUx7ylSuA
DWk2K1YIzN2jE/g4oslBcUDvDvB42GRvxDTsE5lnoMOu2HpvzZYhY1U72Xb3VCsP
gWw6ijK00oTJVNpf9D/ejAuUeA+n101ogY0okULajMPbjl4ZB5zevpSO3vcszYIg
LH0WpAIMg9uynk8WrpVgKjcvfEyK5GgkUlS5IxM5h7XeyOJfO3fkw1IhNbzAOqEn
o59BiyS2gooMmlt7K4ygwL+gqjBXZWfHP1g9jw9ErFukge9U1FSQ9OHCKRmgEkde
iHdvPjEvYtZy9y2SN5jJROnOWhJd9gNxNRTzDFIw4j+Wli+N8mV7FeuW12ljuXKV
DJdRT0OzfXXXZQUfccfJFM6v7goi1LzDpTtCBy65/IY2HTnRg+6oqjx8gCQ0CYT5
HSK1kqhUxU/uDyT3yxRfg89KdCHv+RtULapa8bjKgtx7zIWw5HNiBwPBG+xisKsw
nDPIQpuBWT1aC21GDnTMLGGvDNjNZioZ0cjj2mkgz/NELo2ZzlDP6YCYC53BhPdO
ZEKJc3vASGYqil7fjGizPvdr4rPrMlblN/e2+zbAO4U2ucuPuL+xsnB0n0Tq8/f7
udXlA/Ng60VhRGfEgkj8fyGP9ZZdpzNFtUogeiXArq9Ye6TXXp+6BpeYydwUPaDS
zS4hYG5prk0RaakES6NybwG5/vmnryCN5c2/E1h1MvxVJNMKAngkl5uyXurHU6Qs
7XQ9Sgoq3ypoqK3FwHR5HXZGhE1j+qq8qoocjLZH/oOX78yplBoG8KIgfC5y2y4G
IBPLwi+BbdxNeLecyAMnLVJOv88aHK5C6S5s21aeKuIkXI07aElrHJRo+ronhDJh
h8B6BImD59Aay8iBprfz00DGaMMx/NYMjHKEsBgDNQsNn/9giUT62/vTAwcT42p7
0Q/N6k0Q2MTOobsJtXBbEhVzFiYniGY0rj40YomumDyFyYFzZvbrdJjJV+/bd8iS
YFk3TJ2ea5QX7coevRPHPXkj3eUAt2RKTnMOu2k8nZ2Gn+e20Lrpatl9XMqopq89
ayO1H8fj8btjF8jMg2TRICCzeKvbg0wIgQh/EIThfSHuCZDHT+VXUGh7LSYVSj2D
bmwmL/HpZ1ab3uDP6hjJXczNHuG37OfUq4VjfRup/3+zqe2ZyLrwjdghaOhBUo97
UBPSnYlKS0SBn7jGInG8C5CE+DCbVFRuMWL30qVLd7/2AjgDheqblcfz5Xg9CzqW
fU5RU3kkR10de9d8GoUOn/lSG3pP+8iAVr+oR/cjPoXwrrbY2kHMEm9U8zziqm9B
hu40mYCJEmcv/5AihPDaT7bmmn8CH3+AbB0NC+OAIQRXzhkADK4odsRYEIkK0964
WgbG+QWWAr3BK7kD6woxd/3F2FWjNWIQLhMIbSevUleqhKMztwn2aDuO3M6Xs7Yv
bjKHl9ns1jM6iPX+EX0iKBvFo20FZ/7YWJngp2QhBpYrzVaLFjvsK0q8iXaTIiBK
4cQIm+E6PhRlT3zkNGZEsjnbnd11EmLPdTDeRg0aifU2HiVrhcy6vjuhiw53Buth
6AVkaZXE5ajSwCMZCSLAQMrX3+LEEJ+4m7yJiHIHO01I53iz5rv55ow91o/HQhJ0
LsoJDvqikbUj5lLDslRHiAn42m797WrdcsSwLT4r8bOYuWAj7JSz2H7MCM0IQghI
VtIFSb1To+ivZ+zX3MSRh/PcoZs8eYAqgnMKU4rwmVIErB9bOZAMJLTvK1OLCSDT
+HSNA7ZfkhWsz+9aVdKpVktJNNgMlbFEC5IpS7lPgbQNEiI4CTD5A8f98Bqi28No
Qhf/ooG4yCjwvpiCTNiukzXCClxH3aISYBV4qO92LwLXWzLGbHOI2VDB8rJ0mvms
8H4LHqiY5zWvT6ajNJaysqBOgW7AbftZOCpGCGE+gxFggprd6eHO10Td+5YGIg3r
Ipr4YuuqxPS4AR/hKxLnbz6M0VizTk2bzZFcXWaR0kRndyZDoJm8nxKtwOzjCV7d
7ENwoVkdpAO8gOn1D4Bl+yfFXeQhn9ZeS+yfOMsb96EZAg/NAIgQJDuuVa1gmNLX
QnNl+gc9AgicLtGtutjkuDSyEBTEJg3ExZ63FK3uGIVLr1tFgwpwWmdNPdq0G08M
L1hfceYS+nIkmE/6894IPSIWjHxTW/hYfBqZAEolt+GzkQyBFAyynFIFadkK/VoD
Ad/JUfZPQRCWVF+YQ0LBolhX8Z4rt3lCONzb1xcIJ0MXokjtXfQLOiGjHfIgOf8/
b5V6bii54nLfFtA/wSIN0H6IE3B8BOmqCksdIUto2Kjax13dMOUkaHqzYoV3y0jK
6Ej5pC4AmyiXBTtPfl7bGwbzQHFNpPoBZJ/H0EQMhtMTMOHrd7oKr8bxJz+TSr/Y
wcEL8ioh/cpDREUmdH+30GBTa2sQh+xVFTyBYxgsg/lwM/B4uOudqAq9oESQMfqS
bzIJpf2jWqhKKjzs+9ysXGOlWTn9E0/2ycpRk1RpKtV+Z8/hbILUm3M5MijH7KJx
z+qV8f0g3a1fVL9cgtWvmx9M3f59f9ZoOoGxT5a3tZMZd0l4A4UVVeYI0lg+wv4e
UjoNkaHsH4R5y/VWgRGy6QbqPzMZTcLjdtOr3NCVXXCxJWKJktHnU79Vc/pI6X1J
5QT9xs2caI6XvUtB+cok3iBE8/KBwWYd02UWGhHlChYinHVjCB4b5AKVinefDEmS
VPvHfKq2cmHnwccFSxDJ6/DMYX0q/EcOM+MIZIyL07+auJPvRSnAOg+/p4/dANtu
L4Vk75saFTtWn5cE11UYx1lNnSsJ4PjiScTcikJU/A4xl0QNqyrQWejgFN/d3KCb
iEwc0M2M1JUyBcg3g3nOVgPHt4vlM3GyrU9lRPLMMj1qJN2gcaK9ruQ+yheyVrOm
3Lfi2AC1PviCck+9dGUrOclSmF0wBFT7m5eeDCSBFOM5gc8Y3GkwOLgVNDv52DDF
L6+lqOnYr68TrC41pBQccvsaXhIAFHwAUcESGtBOBi7HMZY6EVjy5qntwSQXnK3D
1WKWdNlEE+r4J0ZNFFrKJE1aVAf43WPHnNoxxWqTs64npftX2WteCJHAGnovki1B
NvqvoNIkjmYWeAQ1gRibB++QvjiZpJHdMUgTgFACBprXk/SUlMSFFpdU/Gw3luNe
oYAScalpskyw50YxbQ7q82HzxF1YNCiUmo+37CFIoFPq7kgpl0lpgbHnoBgjflNp
deDnfqGmEzBvs7bkkL64ZYm4G6j6gV3sXeb7YWlwpPrVKCKUxtvcNkDgXSt5uGdr
oeApgTLXUFqiLOk0lQqG5S64s5rYDSRE22eWrF7MBCvkeJgj3C7PZIFHo1KNOH2d
L/S9tQC+itvFv0wvQqYJ5qPOwUYqFN6iGpJ4vyk1f+/G9hXi08dGY3G0u40NqPpc
tyq4VCdyiC1l4tuv4sb93D3jsEzWQ20TUT5zQ0JHMAxbovImURDP24ILSmd5gxvA
ISgPdne2sSKXr5B9ZvGgwPoTHRsKaf83Ahwh/GQO/w4R8R/tjHdi1JSkdQEaQwgn
mrrsGGAK3OjzDvmYywxV88m+tWgq4KwTSgRR/qycO38gQTFgNCXPscvkR7dYA41A
Kbmw36rIz2zKEtueQcRMcNxM+1QV3SpT0wpR7pdTVJ8ZhgIodO1Q9SS1ugDM9MU6
QVa+g2n2qJMo7C0QexKQbqbmL4flWNwVPQ62tto+oiHpqTF6bc4uubIIem/Ng6ai
NqXXARJHXQbBq9ccYRKu0aGo0CllB/0SujniwQwVqaa/ZRfs4xA4CYrUzjGN51AW
IlG3UAyaAxGUoruTaf9+PjrZzfvfq+UKbmt1tSVtWtmnmDZCwo1EbPgX+fQzU2n7
SIMYiBaErxIVQteBB4KV9uubXRlqvLioH/oKW2YV1sL02d9P4P0jnjVTQp1uhhiq
+t8S3Sgewb25byyJ/E38DlrTU1bk0IyvEiHY7MZnTR8WBkE+Y7PXRjpCs5sY2tIw
30F6P5gdlY/DiAR9UU3buWY/IT2d/RDn6kL89h9YR9+gjxZ8uS6nVc22atGxYAuG
qs4TthD9xKhZU6Dbl0wJ4KN2b8AOPZA5EQjj1UPeVWVt+zzONkWEVB1GR1NZXdZu
957G1brsuVzLgHaw4PTlVhMu+QAzxT4GVc5jfuQInd6mqYd82TQkUCHBRTehAZHn
faKBv3ZRvnZsJrN6BlGIUkNDKfe61Tw4LIQixFpNz0+OZjt9XwQFJ5WdwoUAPfzn
5rV6Ts6i3qYHdQOT3F4lM7pMMrd8jmtvRFDJdLTrivamGXParGUaYJA0/b4qHJrt
Mi0EdaPTo59ZjT23fnbVuR5HTqD6rBfjcXk67ShKp6b4IL1mj2sqanocsT4I/MLH
nyIByAPD3+4otnxjkLAyqkX0iyoxsVTk+AsfHH3shoMmXTFQ644hpvenK0nB+mH0
UyfIOEA+GE5UvgV2gMkX5Xlv4WCOyhAPFqgxpgo9BpuySY5FH4nQIjVj9rGRwz8A
+vCzBEebWBkn5Gwc2fKR3j1rYYyXDSZqmVJcqp3lFf2+6jKgd+k5FZAH9O3Q5Av3
nYa2WBCuX6RZQoHqfN74nzKTG/qcuAFrveXi5YZDTPOLTNiha9QPKAWkwOq6KclJ
ndum7Wyr7WnNgdkJuubQvkigOGpsRKtn8vGEiSkOvtMStyMuKzF85HbtqwDSHnmm
DYxFLZxXplLm0zM8GynYMQfoA3CHbY3vzot53yJ4SmydwOAajksZOzRzU4vNrM0L
qcDeRnWA42aJzBqyKbYfEj4eMBV59pueryz1KVjFyPxTvA2PeinS0gvFvqLZTgco
miavKnh/VvhHV9dAV+rGCY0XsbpzgV2sAedCYCJipJj+ZsjmTcoYeHYJI7GE6lNj
ZmA6b1unGm10nfAUmDfSRLkjdqQt4UepIyH3pLS2CWz8EKOR630utFh3pi3xeznD
F9UlpQaHgVOKJLtwdUmMMOW5plAlx0PMao2JqSMar6IINnWZCMNRSEbyl2ztYd/D
WFHaRpq3tVoH3Awx5Bn+z9SSSEdfuVRXV18f6SNIRLnMYRMftGr8BiBt+IFo77k4
ISmqAzAZuLRIR90GHL0OCZjw2IwLsYXR8DFXx03KgPCoM25x2iLtX8AR2+jdWD91
Eye55zrasYKkyd8g+U4D0ebPIK4+bR7cPUbTSvEKFHY4opicSecGHMjAAMchR3gV
xcWtXV+1MnAk9URY4uO6aQieefNk+5G6sKWfABjRwSaUGEw5DEHISuVIu/gu80tU
VMmv1ou/4KB39MOrNAJbX5lVa5wABvHeOlkEdAA9CalwtwS7ETMdbnEtttIHnENc
KVtvJ8x758do5aAUnObxWCwiqH/AYOM24EH+QUPrI+FEM6z3yBl3TO6Wk0b0Rypv
XkaYdbci1jOQoUOeNxHcC1rbRkV3Rx3DzEmSZRKVk8iIQU3edhI5adEOCU2rYLpl
i/hLvvbhmDE4ETfGvCzd2FRfBdps50iUTmJyUGdEp+8yCBWm1OLJxwLgBEWNv0yt
XnuZOv//1bh94tfoxSnvFHEAjoUfcljmjJqLJeddNR4EWzxNyviBICCDX+fom73m
IXBjndVzjQXgh9bfe2L6VzU2RWELr8g9dum2W9i7vtHMcUaTwCXyVMTR92tN28Rf
2cmgccO7oRstsiCKfG+SBhf6/JlIDlwOMoAHZhV9Qm/9u1rYDxZrviO0HVKSsqEs
`pragma protect end_protected
