// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:05 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pDL9IVE3ELM2J6J5W2N5fZ0bTSOE7C8zfUz/LqExb15EsQoKwP2a8jqaabLKfFIb
a7Lo3A9Z8cv3MTwYpNdkcNR85AYUMoH3htH0XvGtQG8Z9zWRIvI3MJZV/Zx/U1lJ
AI9Y1SQ1BSEnEBJzOGqeUvGrnXjBFx4xgCGX1ahSDEQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 35376)
7S5/JDmTjuu6yiu2iX9pAWbusUGx1tNUml5NNXzho3Akb0VSScI1tdDMJahNzb/A
SY+lpNhEigPLgC0ptaTLats8oD9GCPfep+MV7ArpcsGUrhY2Lm6h7oArO1zSKTdc
UqsWWLQl/eB0XusrvMrZEbTqFyRdzdz/dTkJFmTf0MveKgJGT5dDeZUU1PifcvJk
rBsum5eVa6s+WkGZrp7JVuY3hpCLgwJva5vXVGDGirkI3t1UJRYF2tnJpVNHkLlo
8aPXgWTZKBs7Qt/5+o5U3Y+pszFnZTOlY2G9Iq5fPkhu9Rl4XWh9WPu18zuMz9c1
od4dC19GzNtNE7HCx1ob7ASKiHSICKTPSDHkz5Wt0WDNMzuTq0YfLQj7jmYMaCQS
oQp8R8TAYEv38QxFxRCQgHmsrc0GIm0R5cYVNH2sPgechip5V+V+maXzeeSSFfmZ
O/tBe1WmI/G0ckPoE+1F4QOHI7+IEq8+xlqA4hYAwDMIcwXOyAkk6AWbaOONIM1a
z1CiASOuYb5I8HBTdVpPoqIKILBAiDLBGY+uq5bC2y8W2HMp8mcqLsJINts+zh0U
AX2785gd0yv3rsTyEx3ipwe1xQRsvY5hOk5MZFHJJzl2vIL24PX6mmNnGzUspBwi
bu2NcIanF0n2+k1zICdBVvf4+PqCJz+o8vFmp9kmDMVMHoUt7uKodw7tobwesjJv
/EC4A4nUYfFipsFH8RxcoY46ELDYqYbuZI14hQugLNw+WzDzo8dufhWyvB/ujApe
WACWJHjbJpX8rmDdXnvN6do1figajm+RntF4WOhiV4OXA4QhXeFfD7hXvDx3jKoB
Kigv2w6X8IOqxpU6e9Tg9TM+N/z/mJVYFwZjARsFnEfelLTZgqReEouRGSECHVgp
oMi17p5vOU90XaE7o/rRXvFAHLWA7/bZPXc4xSQIwvEmSplfuHFIsaYp19T+VBBj
SgyteVsGX9A/CS2mKYiqFF4iPjWApczWwqwhzDQdUnzzlag8xJcl0kAWylA34piM
yASOeL3IOgJDs0/J05HPG/fiBKHg44+qjalAJ4h5xpNqPeM3QO0wx0N19hJxuDrR
rSkl5SEbSHV4JAs0fCw5XanVtDyD5EKA6jUHWSpRHKMTW1XxqrsYNaPhHClBNjLN
Z8IzgMU+4vOqaC7cmSo+BzsjaXi7FBICLLTctMm6cIiFg63VUyf53l2oDgLxI53u
b2K3NCjwxOlMAfTjvA+BOE/+l9LGgtSpYTdev1ybygp9Lb8bQh63j8++omijQwcs
jGJQsuNJlZ8/VwnHADKIDUXoOfVgkEiqp6+5G7q3T5adlz6VeYC7RU8Vqu76OTht
FtobSnYDdlAcAgJhjLIycU6U47Tm1F/507hwZH1yZ2HO8hvSkAHtrq8YA7AhEPfP
jAdWIb98ETegA1HFxtx5OdWGAXyjqCehIpRqWabFKeN2wjaHaNxCVU5aeKUGWVFS
GGtFpxxSu+P6rNKqbRCIbqwqysY/Y02ycXEkYlMGQWLvYRNxc7WfRLVCDCKBVPy0
7APy6UyCwxSp+MvMIms6KzhpIRyWH/Qo0eBXYRMqnfC0oI51LUfhwenIcaGfaKn/
IXk7ElcpeGZa8uYotFep5SuIGpXVqE7DYgIU02ex9Idw4BbupF2YcgshsyvwAEvj
sb+rN6RK/2mvmxD9ytVRHToq2P9+qawg3h2OinSAbT5QrHDdyn01P+FRZzPJSXDW
u8NfW0uRZsdxq3JOTnbmTQ1uMqixnyxTT8LaGLftcmKWyMLC0zEukPrHeWneEP4c
eo54ROybo+sFfrjzp5mumMLi84DDPb4Duj6EZayioYGCJCc92OWQvbmJSRzXFHci
9z02ZRxzwly3/aaSlHEc/ZK0LpLsdLTrgWsaJsdmes92aAbkYHJ05kS94+fUeAEb
ZABk7Q4z9uA5tJ0u8zrppSTXCGUmJDg3890bbMqu6U4RK1pvYd3NpN3iyizgIr0s
yv/2PIA9UT8EkNyYhf+gWema7IB5cXg50CQ6PZN78ehpo3Z8SK43ek8bS/6e5yd8
QSyyQ7MRLObDkDFZFyK7M7wuP5laSWqMA5dNau1CGThPinYDSp3AiW/IhkV3MyhN
+QH4Cj8vhppbOs/VDhcgGtwCdaBak2RPcaQxZfejxV5H4ydKFGaiATRtKEy2oXc1
7CD4D3/r67FpLsPyNWVZ8cHGj7V+PfJvJ45ViYOrzdXVgm+P4KVbeRbPG7093rnN
zPyntogkSY27hrKpLY3UQE5twSb7DlpHjgvuC+iTJWQ53Oc1y/mdrOSmJ3RbhG/K
KhyE09rA91Z5qK31yYmURNB3VU4Isk5+GcXcgCJaV0k5VeLOU+smkfMkSjn9J5nB
0fFTvI5AF9LBD+2+oKoFgatbhJKM3ER2VxpZ74YW4ANsr56qFgNfPdS9PwUTuoA3
kaoDIpfOAF8s+pY7eAJjkpPNUjjpWXLe+B0/SNv6sFY1ku8SsEKhvjm931t2R/eM
82iUlrDiynV3pfBN1uxratJrh6Nt6t4CiZL+U3rr4dTWtj1yUf8EYdywHP65YIpC
xdCBnLsIxWXWFJXkEW9mQbo/uPLy3ejNXedqYsl6VhDBrV64+6vHH9oDj7IMiY+S
IHZ9ZphBLwJQ6UkKK5ZPhse/hAcQuepVDvkr8LraR/YoeV7CwfuJDtaP8/vLNDA8
BRIMKdl/wxzmp0EsE4PbHzeOV+hP+nLMW1Yop4KrhCnhLqnLsA5JPBWy+haGv9Q/
oQT1deaRwkQV71bCtfL3cZORO9LxDQn7SnLrnFpVzUXgoB/57d3QPsosjiGbvXMi
Bw6OIQfFomhakmIWTCJZd/XJG42bKdcyRA2zAtTSEHAu1WBLPTAMb1aHKVJKPdWg
Ev+jlKfL5aZNdJGUh0BjrBTTPajh0nZz0jjCMbJTHR6DjXIPTCmLT8VIUcFu+qfe
9TIM3uvgHldell9XIpoePZHecHBeDlh2mArUWLu+4zZjK+1Qi14037HdmbndFvN/
vGxGyBTHZehNAPENH8Pv+RhRU8wt3PSm2PR7M3jmcDXPTHrf+9fY8rhq6hBwj49/
ajkoNv1wKes8Ee2WvyP+SHy/IIgmUejrO2IxmnMLAEQAIUU8zisnMEOifdv6kay8
OjWxE+oS57Y7B6FzYBPbWU83qpw8MQbwPd5PVk0TIRYiGTO7WoJp4Osa2l+6djq8
7kf02tkvtAweifGOqQDo5FPeRqrSgfPwN4oF8Sq9MT0ssDh98AEPALExFlmDFhW5
zGp1hhVqF1HUbjj0LhVmrWkwO5znJPMgL3FXxFptEqaiVHb+8YEQ42qgA67BEaUR
iATPYGeCirQ7WfdMTaKTW259lyTL26a3p/9B4fc2rHFfh3zgKNLPRaqy647Um2ZQ
99p/b9WQuErwxT4ZekC6lh6yM9EctzRy7nFV0oqNQqvYeGhXlUaRzK538C77vzUs
5usr3EVMJPgtubRS9xIRHZBpmwUymuvxH1PKOsTpVYkxbF03UWkQAzXlXq42g8UR
uZWkBry44348xT/SdKX12tjja0hg5keth1xFPgFqg8/PJftiFt+H43XFeUXE5QgH
Ilm4jUz2MCAa+/ASq6WtMXrmorJFyQykYzdCGRYmHlCHMVGWMZ/f52kxeMiWiqF9
QE9Kt72OPXtkfB/GeppKGmSkeUaCRcUR2xWa47Vs9wiM+KFXw6LAI0A1ZLT13NwU
nXTmuwRS9pwRXp7TrBq8Rg4SPiVGV21oCJQ3aHF7fLoaBsI44TnCMmYaXKQVMG4B
G478VZDwHaoEWcssscKmzUTQDt7lbVShKGORtQTYE/jJiaNE9QbJN0cMww0WuOsC
H/rrrnHxfeWiKnYgAbkRBafTM7QjyAfFgxjTcP1HAB1xZgGiRIOGcOFwEDe0N68f
ZsafhxyZqK79tDUjeraKywAwEh2wTcgleMhuM/PkFTMIYKe/9PJRUSu1RWYgZs28
5clCBrDsWANIc9htOHdrDGubeGqHtsZHCrmfF9sSiG0ocswvA7ye+SEE1BrqhEIA
XYVhG9ZTEern5GX1cdwPzMPWnAnC/jBHctcUXny9glRmZ8AAUadawwzl18mDKbQc
RAC2E1Qu2DA6Tv19zBVhNlikthTw2WzKJRqw3HpgO2o44s2LTVNyOFbvkcvA3ios
zqtY/xPjscFajscn2yjH4REyufqCaL9DAZu0nNrk6XpHCA4HLcO5M9Gehzu2fxaZ
Ud3ZgCbc1DvFcqomJKe9GUovik1ysLdq6bUWljS3etsdtIVdOZcjXCWb8LQUSoEE
l2FdLida+OU/c3y9Ww0+X+C6sCRfNFjrHCXvQT2ghNr9PdRk1+waNvaSXNuc8j6P
ypkND6B/eoJREvRt7LmexC6ZbUyy5GFMYTuEMx5jJzS5Nc1ujJ+UrpReMXuocya6
O5WhAiZxSIj0VDhkDAuJfwwMFnepUY/mJ3TwsGKea3dNQVB0R7NbNfVLtDqCyYIE
FLIHULl/HHKsVOY2UNJsw+wWddczbcfkva1c34Ku/Ny65uY392W008Y+pNCchZ36
DOjr39acXSSyImaEYOUYIa6tvXZr/vCJ2YDvLBjcFQCCw59v6EZWmfevv/0NIFUB
EU4bpyGKrzRubBclN4WgImAhvwzoP9S/mUt2oPOuYH+QnyhGVtM0k2NedCgfagAN
Vytt6pZ7bjHt2AB8z9bgvpZT1vL1r/TYOoERXQtVx/5HfXyfDEiCgXAsRZLVeYTf
KvAfquCDwMK8LomTvdMKQM1gcpunHCt0QWZul4I+gvlrDX+/1TToCRVjU/n8msfp
FO2j9QhkDA6MQpW1xiLwM1r6UhmEUq6wuYYJ/4HW0AjqKPJcfn4LXorfnRmj+BQJ
p61hyyDIKQuAIWqhUsgpfkqk0pCPvyE9zs7jfA1va4S0af651kMNderUdb9neN+m
vJ0caW9LwvuJC8M6Dq/CiNbBnCpW0OB3FdOJCS0WCzr485cZ7BbVow8peG9/B2B7
Gzhk/vLDoYZ5J2F+CZB4aoDNPyrrXP0Aw3nZVtH3nYStBa7MtCDig992sdNkE+O+
bZ3l2XCTy0zxG7LpTO8w3jh8W+pkUVFLtQ/4/njvBzTQKgw2FmGFadvWlYI1RG85
pjwU6JnyQoBZY1ozWXE5QcO2V9Gl8lWERErtr0W6EB7OcpbJgE1DtykE/6ypa45V
ED5RafbaVfGFuru1cS2SjJRGSkKkjM3mqf02hDUN53scnAc307X6vq0Vee5I8m7O
6aKw/IWcP7oauuuAlz6oHgAijYjVSxlxOPGEJEGgtqJyxWoZIjtbyA6m6IBcnNtK
WPmg5E5eZlrdqUOzcaDerOBZxd/Ls/89ZBsoxmeNMPwD5tqSlGB8/M3L8laa22+Z
PweTir9gVIK+IZOtvQNQ6arWS/hMT0OA1BgtEXaJQuPl6GpA8hUiFRHBrVgY8L1w
L4T85IwcrrrUlCsJo0vbkc2D4wKcR//afrR1ODcCbOVl09Gy7r7hDwD/9H0LYnpF
rGo6yYjt0F/iJaARLtOuR0kNCJNZh204Gkg/iqbH7JZ/BK8BLNspH5LmAbSaGbRj
+VFD/LOZKumkgMu7CR8XitniC8oHdab5wh9MAKm8uCxji4La2OZt9tO27x+lCTJI
+2ucqSgFz5cmPFHAeLFNGo1d0xmsBJ3xWRqglV4bcL/Ry5HF1QGi6ETdsHwJXakW
7mncBBryWXjPPHnJOUAgcSWpdiul6HcKr41L8+b/ZPaEMIhkhL16XYV3QAUtMCC1
Q3T7CuIhPoCkroc+v5USg1Ae0Z1OKNNvrzIJxC15AIUJTkXXNXMlo1uSi9Wx2l0d
KoN1G+PF0MYC1BK7PCX5Z7O2cmi25PPkC80JpPVGOos76FnJJX6STot/JcJM2y37
TKxGrbYpoZVpQp0kOP6tyCfMpkVfQYTB7c7gEahwMidfKnI29v5DYy0t1QoMUdAr
1lWOmNF53rFKXCV3fQDF0GjTH4EeYc4Kz3rYAvs6X88xq31A0/NMXKgDsJKdxTy0
YyfSzjC9Aj+v0UVzY/Z+7PH3FE+dYn0252nWo79FdisAySoZxYzEInkHKxUBC06H
0ZWEYMF/+y08GMPtY9GTcsCv1+YPJ7DHOaP/fcFORoIcS9eTMNteDYSnooL5AY9A
9MJQEIhL7rl4MT4hIkSRq+y9HbH8y+G/TeDqyWaDBNBHHJw6MCH5GvPeyzDZrj70
FB17pkXbJ1PZUtdXUXwybMdChMUf7Gw+yUg8TOBeWMukvJOUOsShUxcWlqh+VXXg
W7q0DAdDVZihB6tWwc9P5uyh48Yat7kHlLotOH3euX/sBagHFEImlMvR7Xc/2IZW
tGk8QdFO6g6EDIIn2ZaXKCgwNIfhBWG0afVPH7Uc2dgPjk2iHXwT9LBwIGYkQ28w
KtfiQ6YBblI9roUHj5J2E18oD8LtaY3Zi4YxbTNBtMUPXBEIwPlzSqr4vsamDag/
OvVdE5lD6jWwellxOiWIYXcAVdvUWD0L0ICeM6Ah41jsWdBfxBBBMTsZBNQDPVCn
kqZ7SIi3qQZ7ru42/PdC68d3ZF2se9O7uOsmfPe8mCvnyNdWBn51CRNjSH1/xrIU
UCyCbjBp+TReUZPjJotICZ8nVoZDA5PNQRYH4qVUbIOl0rPxTBznE1JnolpjDQQz
9/xmZGF6KCS10hlCVZkZ7eKOqHbTkWjvlLgw2YSUXLJmEzGrakbUAWAWLTK7d8fh
c6sH3scekO8Kv9OWf52Pup8v4o/vTpbEdj0nEeOnw9/2KPL+nTEKJWHXNe6jQVMb
Ksb9CAwBvcTL3aq8D9VsBX4D7eybBab1CuKfCzxP+q0VbQIe8Fy3pyKiBZ05Y0tC
qEP+JdABih6UWHpfebRJEmyGRbOepDW049Xg8WYFGPsSv4Z9zEljnXJV0KPx+P25
LK4cUSaW4Raa35EqK7kUZRQ1xI1Oa+sdcmkuyd3CQKdfLkq2L6llhyMJXg2xHZ0T
KxVUXL7y2QO/nFYKAXLEHMxNyhOnbOQi++/zQAkPZKzT+sRP14fGby5mywcNgsAE
G5GhKnRfO541652vuN2vHjsOuH7hS5VVxVN9P5Y3J4PbkAAfj/LUe+agXst4RVRF
99W3SuYwbBjMmBguwFPt/rTnrEaqqKX4BrEUQpXVm5Gs97rCHxIDAdbAVpRdX5Uo
HzXjUc2T0z8GCOaVWJLXChklsKs/NAbIaSl9mbHlE58Hwn97bpC3BEAK7CDllu6X
dKCNBBBeYj0es/YSXdl+1SI3T5Bm9tRCEvmFozdX7d8095rinWAWGUJmJ1bBxAIV
yyDRYT7cApBYXEy1gByqmJNlzSKdo1R8ILCkh0BTzyuugdL5k8O3HCp/f3wKkVZV
C/ie3r4UN4MAkc0iyNx6o9VZHQcY7y4RQlzCWmgbdz2kcmKjPIhRZ8Np4jO/KFIt
FTEkAZEnNbe6t+MSniiKwQPu1uNBW0cPW18X+JbGBosKUEH1QKHwoIxZM1XsxK95
O5n2TQRIY01VEFcJAEe4PJ7tmj7CDFHlKunC6hKdLJdbum9WoxIWf5cSMtxkjsfS
BaLJirp0BWDkUnDvmVvYZK7esG2iqmQ65GWj3pp7p3+mW96VJLv/lek5c5A9sn1J
XkJz02su+9hQz05qCQime8ezk8XAJyN9BKVFfBjZFz3pzg6oT1IosLPLtuBTP9Hd
4VGox8Z2nzV/bt9+u6qMljjz1zdJ9qzX4bFu8SojNvaUOiDP1yq5nkBJADOnqfK0
fLkfDMRpA8NTCrLG/YGjGx8DVfbDeN1hLduYar6s4IzG8ZaoUa0BA/iDe0zHG4sJ
2H4m7c3jWhvkt6q6P+UjOowBAs1+Ye7w6cP4R3lel6uoCw6qeU+DIpnW8IAu1Rz4
03qNjDf1U9mlzvjnEZFw4WKpYJtzfvrie2Z9zPogTGxDbl3Y0H9gvvbr7EXgkv8a
Pw7MYtHO8Re8yzgbj7SstE4yc1tfhOERc4sqOQc2sFIhYTnmwXPiTur6VXtiQTqN
CANIpkj3eabaZWRnqV/h8NE618v4Mo3rsO0ZpyJBk1UDQznhIbbCQQYucPv9W/G1
ZTLzhEmlSTpwQIZm5KBE/GFgsu4pYWqWFI9SXQPOSyzsL1FIaJ8S6bHeAU9rbjiX
KQMD5AEcZtOhLzvLCYLKBgh6oeA0pfmU5q7plvRIhMegqXdt4LAzffhkmsx0KEXn
J3L7wVkXoqslXellk9/nCn7XCjD44j6M0b6u8oxmZjLW/ZyoR4sa55NokUgJfpMZ
pmWpsFFQjmi8whN+0CXTxxubLS6LjYPzpkU5HvF43Wab4YqeLqhfNbyaPlKBtMns
ie3LxxQHK3lMM08IRknRsINPgRGKP0k6Q7vu0hdJSY4/SiU/qUVmhuqhlFigtqcq
VVU6JjULaSnsg5q07SClwE9JUMRQWkPeTVHNRinwRRvN5fOnwIsjpRJDRH9LoYdd
eNOMhMKniSVjQXmfel12uTbQpEjpQUOizBWaiq0iVUro3cWMvu2ZYkwYm0KZLtKs
VQpJxO4HSbEdAmbaAr/a6Siy1rCDNsrkevivAiTx30LZnutQoERZiYeypDTVqH96
L7cFtvKKqyvfCUDbJm5hGNSQFscHUbMaxjqBO00+Ae3AmLJidh2pF8PZucynkt+u
oZ99jlVHcs5CcaBj8Eh7YRshfK+xrecZPOfD4PQ+P/mSzm4nuSiwd6OJ3ub0NV7V
cSPen6lIUbfJG+Y0tuNofsNug+lo/wg5dDOoJ2y0+d0fcqx5M342Ni57JSWyRRVC
qm7PF6zIunWzhvv72beK5eSdemm5pRka7ky+OekNsE/C3jo9JRa68pxK5CY/EkAN
ZecCwrvmEwiMKdoG8FaB9a+vTHHOQA5+itzQmR+S04rfDVEeqsbdmMewYBl6X8L6
6TGocaylbcZcATNAhCgfCHx+77E8uEJFPgi3Ukb/GhVLv9Qlxlz24atY/37ewGl6
Podw6sWUepYSY+P+uuROwRwyMYQXRwZE4rFrLtqfh40ljV3W2A0Oj0c8jebolkY+
aJmeBfjyOPJc8B5vKGWxi04vvA4xT+yQqnH70P0LrBjNAA1quGtZ4h5EG21c95Hi
2EjGB4p6Vv4S2lnTex9yfc7lbpDnGNEN8BMW/qhvgxl7crnw2X8QBpClB2MO3+OE
ny9HJnSEde6srYk9j37HL4C0/rbxhoIXdFTNJ+n4LM+IMqHs8ys3W5qBcelV3K/o
/Ww2rHcOfigUW+1lGSwCmJhCg5um6WxGwplhO29Tl8pLVsfX2UYjN7dQIa0FpY7l
PjBR1n06xt9OJwtBgooEBstFdIisyEEz+872M9HEXEnVI694FmpuHWeGLNBHilGi
1Et47KiL3CzsRxgtRJdNGqeLcpswkywzRkPHtipPA2Zzez+RWo+xOCeUOb4wQpDu
RoIWMPXRokCI47of3RqRwu0bxbzsrUhDtGnK+GpVB9g9dIVU7x2SF1+YPOKti02j
Thgpdo7j5opRT+CPM77hVIwgg8FhO59O246Rq5NGz4j2xsih7Kg5pn1grrCijXd1
9vnQS2OjLNHTJWItvCPMD/TkHs8IynT44kg7+jRErr9bos5RUaKy+5FTl8tZvo31
xX6tqL9pzO1RioO1Y4gpCW5p47Nnz7QkWSD6SlNr49dkOrCHnPSijqegyKgQOaWz
HY2Fk0HNFepDpTQF2PnLe56HX3lZnAqNBgj0DZTfk//V7H10x2NOkcxjUXncsx5l
ErW8Ff1qgse9ZHuMQ6wPxN+FJwUcGig3oHZn190Fg08AVfhULZqmOZvI76tPJZ+/
mBOrlhnMWsaeISWlKy9qs9/sorxW4jSyqM1Hm+KQhIggrVasKCU6JnXXRWU470Mu
nASdU9gFSyPXwlwt2tFQYjoq0gQDrkNRRjqzKyclq+VG20v/mmdwXZD/37Bu4ZRX
0/xShSG1DiQgNKectzd4pq1bQ2yNFFcbC/B+XQuMjlQUFPKbua34bxDOBBU+GdBk
IMmBvhLDhhdDCgB8Q3M187bxdkq+qdlF/ZjExGstqAz0Gkxy5QZXsb5/314hNpk9
bjuwgtnruIWqYPaj7u67elu7bFY0wTuUcnumRbOeUxouxx2gxnI8UwyS9GOPZ4JK
VmHf2xJ48NSIKuTm5RU6a27T1jS4N4fTe1VeCyioXZojLra96lQzcV64F5H8iBi4
0Xab47nZpfMrb0jtMKNh7NVfEH1B/F24f6UGYAlAqD1RnqwGvQhKwEDlqHNEbaBx
PE94WHrSSSxPzhyJckwPE0zeqg0lHBqpk6y+tJuLGhy/wIXqMnq9Di8SL9w1YyTH
41eZ/yozftQQr9bl/BfaLK5QA0S+HLPVnyO+Ub7tgot6OtkPn+oVOMOWm8Fqgq3j
aPrETPsJlMT9MwzBXawpVxYyeyNGJeoY2KXtfSs+4mG2LRMdPQI351s/sGPW+ciK
DKo6p1VFN57R3Y+OH08KKdd5ai7JZAA9u8g8ummqeC5W/1nrRCrXOdTqxcZ5fOfz
CCw1fvJAwcwpX3QWDGUgv/gUqfEOWXFwGEr0iYRQEdMOuLMjFs3ehZ6a8VXo7dau
cwaxln87UwcoknJCIKNgeNJ6VpoKXgbUb8inBPzc2HbKct1ciFtRNI/R78rNRIum
sROTX8B/KU/rcQ5/lv0/utPRmtWMEu7GIKdhQihsrf1cvV1eqjaUlU142SZ61roz
HKZjXke9m+LtecmvfdyOd5xojSqfQlE6jf4ZzxBCFu37xBaftnKe1s/dP/mkb+YI
yubr+Jo2FP6rZOWH7PK2K420aw3ZLU6ogeYLbbrLhkyEfA1Ne6zH4M8PHsGsdzNh
/kyLhb+OigsPDlXCekrngUSINSYSaZH/wtOlsNMd5wt4l8kMC5pIlOD2xGprWprb
28+q6BH76KW6qXwxrI6ffhvLTtuZDm3KyS90CYCjUniq1aeT0JIqeoxB+qH17aNb
IgWS7mVuDV3aiXZr1sdSSiRBa4rWlLLxREnfoLgfTSXWktJGQAYhULa/+mLQQ1Tg
keCyOJJfSg2u2GybFrxqgNUSPw7855Ob3fQmINsCSwcaiGLwBICbwdb44iTkgDaP
dTI5arZXyGK0Ys892Llffo8PR0GThFsX87FcKJqkdqLN+8END4v3kgcmhGdNEx8b
d3V3EG89igsEay8gFdnQ6sg1QWBA3JnkCJnDy62Zwgqj1mzBkWV/ipz+tNC0VxK6
QU92vLeZEIKUeboXegZwCGzoPOL9Dg4l/4hsSwQfQWw446LDWmzgjbXfmA/f99af
MjlQD0duEcv3HPKOIKocesiRCKNZPFPHUHxp/U6LAtW5ObaHB75t4Uxg8aQikfGP
Tm7ESuZccJ74ea+m88YU6tcnyXq/lM6EBTAwnKEpbVSdsAxuHy4s1XRZSpAL7Nmr
tBCnxU+w3Kotz2ArlNJgz4ywI9U0wZl2sT87wnCCmkoQPBja40iZ2kS9GGenqptV
IqR2hW4V0SjIzNO2T3LO4n+Er0dljMIxwCr3gqDwOl92spM+YoSoPWWV0ZLT9H68
Q7MaMjQNHmIgRh+sF782R/Bvd0z4bf8KXNadNPLGAbvYRYHy0WSmQ+WfxgYh0Il+
tZ4H6UOpmm6LF9kKd0WG+Ni/xlhYoD7DvmhyZIpCkVblPP9y/tr1T7JDyrVVSuAx
TSU/EluLOZAmhTSQGzK6yX3F23NJZoslPMzJ+HMToCTXvRYggCqP9nlLohkM0o+Q
7CCw4ooMDZ0pmpKDlcvX737Oh4ZJCFKdCN3q/mEekgCqnIaOT4lGO/M5KFql1ne5
XIB/0B1tP2/QUNNk8BbIspX2ZjYZSWbdyN7BUH8kx+uElTOAeEbrnPUEzQ3qhAnO
c2DFPzEe1fFbZBQt3MH8uKWxT0bnm0LIVzUehdPGPmeBXjfLl+rkuhJ70QrU/pys
D1T5crsYTPEXMO9Ho14m+MR4HxB+M8l1KvZCVfuTm7V4v994XjfmpKprkDLddKac
GLdXwZxsfIzqSSG7GJ77nwhUKcLkyrUm8kKDdyPNOn87GaAJfuXIMaJKjc7qz9+e
5Ss82wvHyVPPvbXVAFVKUMr8+MUqEg+lmMO76mOAuWmdYfdq+1ystLz2x6MyGJyc
5G++ghgXhE1mqV2J4BSt+oL2FBGWPYgmlBqFRyeB4Djn+IrNBe2HDBkgHCXt1xkr
CKqAe+EiVhAw3tm2uqRp0T1+ahRAGIhMk473hIz0eNj5Psz4P+9cpDC8u2Ez0Jjb
lxw7URD6EPm98e2Sx0UhvXpzNN4vKoNLz1+Zrl+d3+JnwyRuEJU1/9UJMBhv34q4
Lqjw9Dxy+4QipKpgEYYaBkYSiWXe5wKyfoKyYwnrhP+rt6B8z26hC0T9diHroZnu
2pj4ZoB8q3CcLHQKgfha7CnkjItxZqAOWOyD1GmurV7a4fEvRSD9nLT0tiWhZtgv
QNPGCDmoR/H0FkrHvJDd98zHpfwm9a6hCjMfZNS885N85Z5uJfSxjdtrtFbEZxbc
ricACBNwVI4p6ATbNQ08bkiPgjTlzJQVUFhmI/Baf0R3Uwvy7DrkEqm9AGfpzzyN
J0AkIayGZSCHuEJQVHmgNNghFcxrN3NkKc8rXi5suBCBKPUu8sKHxNV7gYhEg1/f
GWcTZf3x8OSOVjZFhUR2Hbh/yr1owaDrRizLyH24VJKSKdexSMUFDZrmx0BEuytj
zfrvChg/ZIq5sGn31n+heprASH5+9Z+iqJr6wTMW0tIedPNrbcyzMsjr19n04HGX
8MwExlH0OuJCO9OL2VBeEEWKoFGkETKeXHcCtkqpVg0ibZbvSEag6jOrs+ti4+zs
mhAwtW0pX0gCar98IdVUaTfxEbgEuDUmySxYPgzY5j7LesZjsyYWChlfmnY5yf03
uLCYxeOHZ0jGVJ7QwpwaHjTZnAuPxzAxx9brmyNh8hFYD22x2mWHJMHvn0iVg5ml
OxQHphisXZCS/I1FjumTkpB8YOyfqWVfAbbrtGY4rmVGkZOfr6vOyGDEt24vRK9b
0nchhr1qREsP+eOuqSwRngp46Fhw949PgQoJO6kvPLDtep2O7yyQzT8nOD9Jrc9x
GkPnkLfbpa7cZBtFLphdAaqN+LVlKUwSAp5QOsB+8yLw27EG+YbSnP1mH168fgol
OUSNw/mSky2bGJR7DQBzeZm0p+5pbtjgvfBx5kpUJkQEfXbAb5FJk22c+ygMOH9b
LL4yqKPILGtwYAyeuim4wxgBQQxfEa8aRzTu2zkgQlBoYaF+TF0V2RiS477YPoPD
sWJzM87eQ9bdlipByOjtjnXbJNAcC55i92TLGo9Et1gJCmvLRMTVaBvnXhdQRy1m
sTd77dOZZR4evdat2g0jzZzJMW0Dz7EPFPCraPtSIc3udlsrnX1W8sUUmZEu89al
U03qAaLQSVPuIfRxb9/rTvMcYdCDwQgI/3WGhfhgNBbfr8MHwN1Kxj7Pnh/klPG+
PJI13SbZCQtG7fpEwNUkRMMcvsFCCQp+FgIq38rmbH6u3ugKHGK7D3kRVyCs8psh
KpnNeLq+yaGQbScGXItCDhN9MuaWmyAHy3j4xM8sVGBjckQ1zz1jfpFPf7ojENsW
nsCHAaBeNIKcc6DOVRhlZrJNdqiSRiqbCMShxdGGalR1PdyW4uxbzCYgFrsEYdla
vwah+P1BpDLgraz5zK93nTJJwWpMwtj71/9L9eVq/yw6I6W4QlIgDEPSlfLrZU1N
qPm2FHIS2to6VmVMuuQtCNZYse9KG3j8e1J4upRrSGSwuJEzNfh7Lunw0Xi5Qvim
lJ7RvaB/LeI2igugjXV1xVlHkQmLKfj3X51/nOh5xlHmosd8BnONSEfTLKyg2atn
hQ974xWgDbnppVIUGxKXgmV7s7B6hysQJJU7icXPmx1IzdBCjI18a47bXxV2BjvL
ab6Ar4+qUkHOTjGm/NeALAfFSL2v7AlrKUbf+qlYCDFclul855VBqyS+JkuN4w9f
rMwMz/c7ZM46usDMkyZg4tGu8dzcrugv65HdhaAj+0Z7qbt1Ja+YJjtmKIn1ZLUy
fTdS+ZqNxCEIDNGtj9tnr0IrfxjIxqPly1GuQ/9XasnhEnuoXAxSiURZxgXq928f
nT6gaodBN6JIAAUlU09DtMHKJl7elplJDPyA1OdSxZIsMsS1bxoKS9Xm+r1J3xVJ
lV7Wfn5u4ge3Y0E0w733DOPXnFfEcSyWpIKAK2asfLrah3MC+Nau/qFjNXZbm9XP
e665k/8MevFYTzhlV6ec4m82ld9RYsT4bV04gMT45tGotUo1CG3zV65+ZMWOVXyP
jjgrg8geeBccVDW+fbcKu/tyq2Zsw7JgmxZeXepveXA+ftiJ/jviHEAD0I+SLXSz
gqH6/aCZ2Bxyra0Wb1Z/pREvtIX60RjW4NmYm/SVNKKiQbWVxv3pju8OiVySckTU
aWkh8a0ZMjGoZAHU0xleRl1NGnXmQoNyNeNqldWWyCqJXlVkSY3lecg9GrsvgPJr
2c+GoZPlcqIBBlALYtG60v0g4gmpZ+ypaC1UaTRm2ViwoNS9hWv6O9Gwnpd3wBp6
iTC4u0D3OprEuPoE9wm8+fvrRW/kh63IZ3yMhnQpCZ6XTUf/01x8tKagehAMxevE
lBQshYj/07PqQARfd5o/RqA6AsGEjzpra+LqPc5XESrzF8UFcIf27saDluWHzbHU
amJk5teD29Q7tKz+yM7sh34OJQBANGj1X9UKc9Ytf5q013fID2izXhdbGdStxT3R
dwRzjR2VEuGZOwWWWBpsns6U/x8Mdn5OPLswWsR1VCpB5Y8IV4tSESP91DvBCIsq
0w00mG4EdeVTdPeOKsMtf10V6WCebLsqhyyE4efbs+bivi91zUBXA+canfIagWrB
lvfJKB6QDWb1RR+uwXgZD/5H4A2uMNZ0yHevT797Y/6o3NZLaipBrB5ShFP8rJZJ
kutqhjqDAhwD7v+s9m7riXJQnJ6x4Q4nqQc2tSD73JhCJHy0qlsrIJNCumqZtrmD
nyaz6MOuQoZWv7iHYekAMKsQRcSHk52HEUb3JFT/11O17AZcSQH6zt45kWj+lQew
nQGvbwMdbxbns8v0N9UqEeIeOn3gsocupFWqsLCT0kMAxk2ln3ixyTWUSt8/dXHy
r2hOBEsPStMlWbUNlNz0PRwMpoXzmqWkeZiDUEUJwVa4JzgGBvLmIofy6oeGfPFp
xMZaxWf185dBD7VDvloVQkUbe4ezVDCZyAxkiOVWbnaalzQCUdbevNhmRWrTrVju
OGeM9gKwT2GCaQgUj/DM28YtMJMLABOWToSi5fdL7RgnJ+Eoag6Y8i+dj2PtKLJq
y5UqW3Bj1JGJ7j8MQC5GBZvQWTEfzMM5mQjtWgsNccWB2OnusLFu+1hqsbNvIBbc
ahFeuN4VCew3Ty+H9KEhCBeaUhuqHRfTOa7XTE7Exb6xUvSIfJi/mGbx6+MRJFLR
l6fQRk5Kl4jeeWVir0hTTXAWIalklPhEcF3DiyuKvqoVuUvyVJXr7zdHWvW5A6HP
A/P1PaFSwix5DNABb8FCIn44Nhv88vsvGrzaGY2zgVH4mQOD0l6f+QOKuBRHaDxA
8r4c9liaCVQQwby/IJBi855huJC7cXAueAfbo0ajWrQo0gP5g2hmiLTYBX2G8sls
WKvtKbW7K4ogOJC0xY3dg8GXEbl7YT5fPPNpHwqp+Qd9vzKS33RhhRFlr2oGryTl
xEHZBs6d5h88JB+Jl6jlnN7I4OBJ2TXktG1HVoIbTLG/N3jTD4MSi2+PdxQbIqK7
3D0KUtXmYuHXphrCNsmdVYExAHTPo/pEzqvg3xMBLJOtadcEJ4NmTNbPxoRZO5No
wbSGGNOGPJR1HjimBu0NtTWrNjWsBMgDqAIqaEkWF6FHiVcKxEeiUdn8YxHem/Qw
SSV9+xlDG53y1t1urJDR84ltNtHy0fEBrueAtyb1lRmknKt1zNnH8IQAjCGxyYVk
SK5VgKqh1c+S2VTxqEq3DGdbnabwbfKMvAAn58cndArktgmRY3T3V0MXELcINvdm
U4NEiMwl2wvScbBUA11kD1x2CO/NA2Glzqy2rwPL7JUllCf3Zxo2xWTAoGI1zbth
h8BV4xZwnqyuRIQXOxdEaTTeXKGl04FINgB4U9aW4OLOcmOAJZciHp+jgBF3WT3g
e3M61/Y7i6ERSpahmajExrqSUpRNTGojg8K1RerMuwB/wNggrWJDTonE2PbK9sBa
JneX2S9kpErXfs6JYGfPFelwvDlOWv7Zi7H5BcXu5l86qqY8UYFRINL9ImNL88No
EQBraFXuYpBq8VaZQycCrxAkqZ89kO752xzrJD4eTaLH/+by1BsW+8dSe/gt9g5/
qxh4O7+E3R+JoGl/bQ0gmo9OiG3beCTCMYS44eiqP7rHNsUhChw6MnKwMohBZscl
Bc3QCMOiTPxWxvzj4cL3gtpdUQmHv8/pi64I5aV5scWYvNMud0WVNQJhj8rmKiA7
4oZ2QqpksDf9gp7/aC+ISfhUkZ4iAtdzO6omU3UwOifm1Ty7ATv4WEngRgfc2f+0
zK38w6cn///uyz1btInuLgwaA3Ke91y9aQVjNtwVJUzNcT1QkVLz0UCqGM6GvtEn
VcppF45uJMuE856FMQHDrmYzSHFFZ+EhNL3nIAZInZQuJYnl6H2815EhJmjSp4Cs
oujYaWSd8CNWq+0zfBzHinS6oHdM4CZVmd1E/+J66rWuBUg3bL3TgTLea82pAXDW
QFRJmrzn/g0209ktuX6A1bG+X2PqeUeL8bbcA7pld7fjBQlP1W9RH/sUxtzsgqMH
olYyYvUGKKRA+yOMuyKb3wsfvQ9M+aqrXa4KzzcqcvntJ6v2ZyneQAtrMgJCNi8j
Sz3L5Bx7LFd2XFr+iPMjCUf92PUruJnR3eCRngu37P1lio8Dizg/5hglHmP1qIV5
U+Gfe+/+8G/+D3A3xn2Gx7+RrTIwF3aVJdaR8hYN4FhcL+OhjL183fcUyjaNP0pR
lDhqL9FKKMEPTzWobLONk6BIhbHJKP2MXmwd8euD/Nc1gfzznuAY+PzonKG17XOk
C1GS4S9i6wC9uNCfI3YmKC62gBZFRK3Ry6dDtJGwYjzeN6D/Z2JHGYv0DrAIk1kt
UwtTERrSCdSqYCQtU7H4xBIWbUZkxxodBMAT9g+3YbypaJjlteC/IRatj/Yu7FU7
S8snPgH5R0gG3/Ljd/yWx7HkkaMttiE1iPadX3kNso+rQt7vqKxMAYZUdKUYqi1z
cfDxBq5a7NMcIE8UpaW/nY1uCFE+2RhVcvghemLVGXKLZYoV6IU2IYIa4eUIUkdR
kuvBGsZB2m/esr6Jx+U/7j9nLF0KmYLXVgWWcQ2eEodpNAU+6wA0/TQB/msiem4v
dwxJ7cwNxXEAJQz8lv9NlRz+VmHDaovHJGx85PH1vJvv4AaieTvaDHzNq1Vs+9dm
g78hUq2/gSpSPcngi4v8vZSZ1mpYQjVWOuJGi8HCdeCtgozyi5ENkqs19NOdaqZO
1u7Ij6kDn6qIMZLpKvCMb/zLtaozUIlrZISO+36ARzxYggATFmHctZkMWM0DCH2S
okk6vRn/i17m5lP5xG2+BQ/SkMefHxmRWHHATvMg408qZNrhWSO+dda+HvhM3s0v
+gHMUtcn11bBIDmzsuQuMFnUra+6mGFTR3lYyL1N1nj2hNrlAOVQKtOHI8J/6Is9
rRN2Fg/ZihVD4Yj2VLPSHv0G1Mw2IziXReBmG516LV4VRXZdi2+er/gY8uV79/Vw
KF7d+RVRh9NQpkl8BO77w/xdp54zTI06WVQk6dhmdjGniIC822C7KX18jHh/HP+A
fnJY9pJUx/0I0MXaEXXSxFTbEnt9SrcpEqLFDkQsiji71Sp981xw11GqgKY4aOxV
EFuEr62KzIsRT+pdUSISj6T7WUhpJx7fDMLdo0QAW389Fn72zrn4QeTdjiKAQ6ZN
vWlAWx+xvrxNllCKt3MHuK/opRFiBj+tEwdZX5Pwnsb28Qt58f1HY7GcRjIDN/25
HfFmSNKZ2lj6ajixU8Btbk7fbDE98Cd7nhX8Y8CY2OWn6van9+O/cPJhDmOwZQat
kUUH61SJipib/bY+puFHcX+kzW6cqpLmTcafr2CaXbjKZO5eeBo+QD/b/7xSyEPv
JHhH3gpQRx6V8Bgfqsl51mYizRw7sM9EqHxhS2N9pUa2bjiWTvSrE7rbVEdckXPP
PQKmzaz3q8M2j9Kq0Crh/WlUNlbQ2+WFSIPcky70gAijr0MBxqGtAYuz5UmQfVDQ
Ur21GKOOFv6SV1/eiYm5SQ6SotNrfLDv3/t5fOAGQ4CCuemS4KwnPb/neyiuvaZc
Rg1f7In7LNDqz02co1xnoPPwfJOlPEH/KFpqvcVsPUgD2blBaaexXcTtGQX8lWXZ
2MK0sorkzNMnj5A+uymTuC2Th7R9QOWRA3J4HC8hhoPJjeAoII5WE3T9NtQbG4fw
vlAT8UTOmgKjtIne/PbmSgvdTBkjKCP4gJz0Jclkk2cWTCqbNhFAaBUqUsXD0yvW
fRoVzVHkDMlZr3NXPDsh8AgToH5a6VexZxpdpuLY942N3GNKj1Ramm6z5bHfPOau
cgBCochkxXtBeUwvg8xK58e5NCHtAH7luP6xNAOfX++ohYChgo7AGINBlcMZJDnE
A9Qym9/h+JdR1C+EfVFuxKAKegQ81X7M06mw0N7He76buM9l/gJuD2e7nyCDrEi7
67cQpEbbQDGMN7ItqXIgf2FzoUs2d63K7x69JojolhroWwUJTn9fOMcF7v6Z/9vN
EOKrHsdTQGKeqWpYkZ6aDVl825jeC0SLUD78Sjw7110ZTJXRdbQTDrw80OKi9o1p
2qPHpYMUiaNz60XUlDjnJ0Q0DPECIFvBPsmnjpHxvKjc5bHRYHnrEDG/0en8QwHy
YDuVMgi/5zUoDl7sSUB0xn52TSRYnuGizCLM0+0mF+lUVy/UBHterO/SLb/6LyrP
aaOe9FbaS9ijE1zQdzDITlsT8wIanvX0Tqke34stcOm1y3jNVuxelCDm4h9pHfKv
/620dmVS0SBlVeT4aOmWwo2xAZ2XyNJP8asnHmJPZhbGJAUbGUz9mAuiulfEh3Z7
VYwjCgReZ+I2zzJUlpu+ilpSi17PhlKsX7FuAlxwXF80V94EQ8Ip/mG1xFhYy0wE
jnZKxdip12gxZrJe5wxDkokjUw4pem1Za6LwSBH6DEsZDnrjon3MPl8U9SvkKF7n
7SXgHqZia9S2lgiFPUt9zRh1g48Kr3CUFl1NWOcU1OlrMv2FtrFAf8K0O15Pbh0m
7CwtWY9Soqy0dWe9Ag9EmcP9sKFmtsbcp93IftSbXwfA/Ih6hLlS9+bl0/cvnwiz
QhqJT3wq7nQG6aqYddHWh63N/1S907mdrcSD87Zs3xD4+4Q0FsfOzpBIhi1mKvXg
phCQTDjuYDFYKAOnwKxCNbZvXweDU/qOzNYswpBPPVAdJJ3hdqB3g9b/1DoQ1cDL
SvO4xzSUZvEp4gJUWk7YjPCquOg5ACZa49R/rF4K6rOahApZsLF0ho6WRwfZhz2S
V22M0/sUO3q18YcGSQVU5/qqfp+JV/QsmLgBOjXBlzrczCAMiPop05ioQRJfgfwE
8e9t+pZYSmWLxUKoFvZ/nh9V0FasCcp6F7RGtM3xe7XmPixQRGTSN1UtjGE1WL8T
RRy1w1TS2ud9SEFkxL7Aq6NxAFgOwr5lBV5n2l2xpXg2HNTajstbNaUqFarzdho/
yOP6YxX68R/ntzuOh410GIv4ihV1ELZwnfO3/y4qhJ/L5YTsrdLvQx1+cANOUfI3
Jzn3GFL+qTbdRYFKCX5f6X3ITEdQPKBUZKWXD43zbVZbU+0AfYtS9L5PfbM4CRoX
COYfwLKuAl7oqT19t5YXJlH0yX2nQjVZI+7RDIWaWhE9FqVduXLYe8OUqwt9rMrV
iiRMITpsPXXGTeERP1/N9eRG61ykB+bVUf/R67NWO6/o8ggvJj6uhfeaUxuQiEl+
kRlPWky8fmAaEAXhQd4qNjrVTHL7tuh3/vS+xgAGFgcGNMlR42jSWrD5tzXH32qo
dseb7r877YyJv+4I2xdtLudocn1A+I0Bbs9C/zc9QFT7pp8II86KR08i0z6Lxr7p
R7IdWgPKQDGPDxnSYwS2i8wg8H9mTJ50NAaYtj4EoWW2GbgUt7+vzXW3LbZtevrY
TE2NKtsV6BzHhfa8adFvaP5EUFRmkMsU3kGGVrKcTfXHcilJ89ALm/fzJ4gEjFEe
aLEfzQm8TQniz8bgUu0F0ayKbElvQK8k5DdGMmQSEomOrSp2yLGF0tf3ctPdg2Kl
WZSSvdPvFGeQEz8u0F3Iw5S5PQWZ8O7/U7po+gke+s09Dc/YYEuwZeDZ6G3JBKhO
CStWHBSEMiwdebDOmXDF316dOvMLecEPeK+PqO9Tqh6dvXKEryCvBEDcy6bVj4w4
PRChnyVT1pMzQDEyJ6H7sVi8YiW5h6A9lIRIpXzr4ZOtVBGeTMfO6NOVyC8alhjw
4a7fbFibWNFuUyIWWhc5iLHs+Hu0/V71ij0BIs+Ox/9ERIYNSUJwCI9quCrkU37X
eY3TrbkVhQpG9DaXzIoK/haL7WzihulwQwA6z+R9Jmnn/7HEoG0ve0Wrqsrv/eHY
xu6gePWX1GDAMPjPPNp33YfGQbQA6F/rKbpQskO3dkDydTaWzhOF/Jwmfy+7kbA3
U9z2fmb9CkXm9AtU/ANBQpQWn7ccNauOZ4fnawD+izEXjQM5ALgQMv5YRzprL3kR
z+2BW1bCWT0UMujV20qr4ZCcY00P/AzLQbYr9m5cPowsUEFxKyp8kXX2StgjJOot
faDsPLzDpEsXk8a6DpsfEuKFfrRxJbicW4KOWU2jCGJdlJvmI6DA24+xU9XVZzIB
flgbow8grIU7U+cPdcoYsP3k6lueBMEIs6Mx1BFUtup8YSannp89mdh7V1k5L/V7
DGQQPkL71uY5K8WKVNtlBZcOP2BwAh4zE1OOLsMen4O2OUDFHogbqb1oljf1A3bK
ua/VfNrrDp+jgfJ8cV9YtAwv/5r3PiKjT0pFPMMUsAC91xoDdjvHLQ7VY/01oo0q
ZvluECSCAMQaIf/8jqGeXtBPLIYseo5ds5V8MXBPdkSGouf2y08Y8NEcy1s18gv5
Gvsl6It07CC4jenYfQny4T/re+t7MT/LyKISnkzKazgbX4xcbDBTaryn3jUvyKQg
3FJ9UhVdqYhZTW9D3kKAUMuSCwopvlRStqGrTgAMOIzio69keNQ8NlN8jQaIEEvJ
CzSFseonfA3oyJrCDrDgVMds5T00FdE/zZGNSye/mEhTTVPqFLb2uNnJzK9odXzr
CZeAhHSFDm9DCSH+e89Pn8DCE+w/dTXWaPusTYe9Dz29CFpE6i669AvjD4uY7kG7
LVzHWgHsunl1Ck4PeykjszdLXeAAnY9GZUWDraPtBUs915hJ9YQ453qjkJ8k/PSz
pQ9Vxc9yQV/7+xn8dAaHiO3kBavuUn1i76FugEW1xTDg+0QKzjQR3/nWPusvjonD
Y3R7stVLlGgVuGnT5DGefo3PLENzdU6wU76dXH4J4pSRNm4XGFJxxjySn/0xUOiE
jrXKbc2ZtHo7AIYsUBc5XUdrPSW9DULmNR/We3crA3yq/zMaTjVn5abUABwNBaYw
RxKwq0qZzCiX7AcFpFkKcmjJ3e+6S9Jtp+m52ojR71za5Bw5K1Y1nVL1Y5EHlcUt
0B75kEzNO9Kxl42CZgVPYdzQlYXGJk9oJ4J2H+bv3xnY+DkRuYdUwN1tLuQU/DG0
hlZBNvw25QKD1ZFf3GP16LmmMzzFV3K7O2Wqu4BNwi7O7oR4W/n5vZljFeZBW4z8
ZvTMzIU7jyEl5RuVcdmgd+g91AlIMwvp9HwHphLGXF9GJNjsjh8ARZMEHQqx7/Gp
voSy11vlVmBozzwJ4uBL+cauUxDNK8X2d4g9G6nQE2yoMhrfFCNPVMTbjgVoHUgV
3X3tdgdCoqJ2oDsQzAcb6hwjl0APPCpYqJUO5OV3QxLqGIpDRC1wbv3Stn68w5tv
m48I/lefx5eieq2VS8BH1uyLGymS3sJDN2l0KDG1P7+8hWM4W2GNyez0lmtQ9S+j
++LgWB7FoPCgoQzAPmf+6rrnz0ALDFazE1gGDKUok/Iy4SHCHnMRW4x0rp1VZmm5
NRDmdW92WIQoUDBaYa8VF8uG8rbxQsSnnOD9EnjzfNelr+U0Wx6B8vWcHAKBcu4w
hfrwbDz/D9zsSQ2ft3JfMH1BlV4wL5I5c8PzGS8UnCkZk7yNfBCHAqPowpBv8uyH
hZr9ANQfG/pELFP8Yp04Xc/Jval15mU8bjJIRxhomZNAoVX4Hr7NqvhEJnvDIa9M
FVjFApArkAi7EsBvlUrxiW0JLXMjV76huYpxvsVeeTJQ8yB2C/bWB4TtuS2ZQk3v
7DPCHuIyjdJfQezkI8qwNzuNtsNxueLOPmWQM/mhp72ivLlvVN1UcNelDyWGYKux
jD2y0mDVBAhwo03IoRg4FHKO9U1/j7BprXZeocDtpA3QgLAhb36wbcKxefQPJJrN
VRFVWTtQH5Ty3811D0yH+NbCSwhAZWR/keImsD1H7EzkACGHjJDGsGQBs/ia11uC
Sr4YudNZZyMa2sXiKmWCQ6U3EeY1mdCKcryQYfoFoNXVpXCqJuHw70eO0m6q08s8
3cJhWWfQ6dC7uyTH9O2r0iJ8kMKQZrRAPHLiZ3fTLoKi+Pq4IW64DjH4kQeJvpMo
+YnLHPi+U3FIHTvsNXlbxxF+HrNhRr2YIeYAZf+GMrxs0x6lFYC/Q2Ss7QPr0aCp
b/FEIdKCwdu62Qlp8x0dwnP0pAAWYYmFUFHSbLlPsoVoS6aLlvjj6S28jC32cv2h
A75ySt7SjwgSl/P8RFABRhW4i47EUu6inBMo0lqxGzzDhTTxHbbwE0ZV6OxlJsgh
rAda2kpPFyZ+PKgtw8ofW3dkEcTgbbRyN5qY99iKeTFrvoIcbNRA3ZuWn7mShOgL
FVgtyI/MjbmM29k5rf8O36CNLLheLkWu4HDOyHL0Mq52rAlZdGouQzjHLZAhpXe9
Qo1xbWa/9qEViOBZmmlC5Glc4H6ydbNCQFBiKyh8bUpcKFM8br4MN2+8kRsKZfHZ
AIX4gl0ih2WxxsKym0ZNWd9EZS5Dv3r795jetD9AiDG+0qS3g1kVovgQFeggaoNr
l6Yywjw92IAlmiTdNo40wvJU7OCBO72qzFAnWshG0ICVsc2KhAs+nODclHRcPEe8
jSqTOTw6/Nl9v9XOP9I1hatpP8Od7k+lo+u++SSS2qXjYLRt5AXRgyzf6eKuJ/+x
RPLcE8vUHl6Gp4CMp8xp9D6E0sE6La0TFiTsStOAPO5Qlqcl2VO8Z6yQ9d1xgL6Q
ly3NrRoXHTGfD4J/f5GcJB/gOCPiwhEv5S2AL/00mGSiF5qA1Ot6GV3dkXiV/wXd
prUJvOie52asHCyzJ3qwg8UGScosKw4XMN1R5caBfWJF/EHbLbqMmirUCNBcpkGu
9fJoCYiIXbI/xKfBYjgKp1uDsXPlm4SN9i2gs71ce52jI4AHsD+SoJ+j47MM0DFL
+CVHzEdGUVg/weggnORa6YWVpXWTCEuxSBZ6MrnSz4krB8PQMpMTwD0sHAsAE37/
GQnsJ/tSJiOeHTYuAbMSqWYvBTdCY3wWPvNERvdBFC/TmRzbpaiFpo4NJgFC7ZWi
33QmmKLYMKeTZV8ILhiFvE3wq6m7hwwE4S6taHN12ksK9amw6nZ6DEo7Aqbwvz20
fs7/ScfIVs9oEUUswwncc9IEApIQexb3LMrf7KQIWDktprs6J0r5CUMZ9blCNrmH
AT+5v5w9fIGmbLMkLRWkoNt9H4DIkBrdewnv+Zv9vhv/UIgFB6pPCHJLAH2urjmh
873sP/tRKCFHJnCgFOM57sVNexCa4rFFA0mi1xxv3QOBtliNZuNqUk0ROCYqnYhx
qU4umj6H5y4+nubjTXzqUXaBczjvJPF6sj/WWIbjHca8z9M4cVhXUr70zM1HG0VN
2caNZegROQa2tl9va+aIEaFzOvVBtLkDZ02E+tQY7cf+kHH8MBP5onRPjaf4I1Zi
FcCA5BxByyhENFxTcRS3ilPweHrQuGKt3DkzQeVH2tTKXutxJjmjtGU2qns8CPi9
5Wu17P/j8JarTSVZI9P6tySxCNKfcfMojL8/QLaapm48++Fc+yYOzAcfUFufvPh8
p7rOKJsQWipZ9IiI2hFO92DxUBRHEkQ8wNNHbkilExuQeq7YASalPnD/s7AY/FHb
MXXYAFmb6KaPv7gwpN07aB8+kHc4rRsyk1+yRCdY8aWWZOYeyuuIhbOrD8T1GGsR
xCEyASnmr7+5a2qV4cpt6saPWN/XQkiq4d+95De40YZQyrbD6cFfWBy2ysg1R45Y
Uy5QiiePrIwTWf/DYy2UfowtsPBMEig7ctYnPb36PiogNSZ3bHl5aWvi+wLqFRE0
ikbi6N/qLUoK5MpkAmAG+xSr55C56Ts1Xx2pFrWNvdRU4HdmiG3Si0aGwS+kNoY7
jBH3zUyoKUNDtKoPJbRfJRiP/Cait8og9LCWNIh5AyDpWYGwtOjRp96aB26ySS/2
WtQ7m+JqHAnRsrbKt/H84UZhAluyrPL+iSjv9gWVR6Gs+5sfazvU1zCpQlZjVqB+
PGMZUMkjKGsnbmJ2Skoy2HCpAm0PJXzlJjv42hwzabBlJhw7BOes1Z08CvosO1/g
hKutg+GD63UA+7PckuVb+xuxVeRCEyUyOuIb5y6JF9afKpscwcMe/vpn7JOSapjH
nRlriCsoTVjwveIgHJspu5XgUWoDteXqd8q9gfSbe4DbvJTs2LwOP3ocSkrwKZng
L3JUivBeK/vUmi6mnGrwqU7EfMfUfXKZWRlW+LbLPY+GyF+OqL2RXdfK8GsTtuLG
0hnYBdmkhaXTg+8SS83Im3kdorXgc4PID/ELDnxNBX8lJvkTc6T6DCXcA8Ir5oMd
iWE+qqMeeaWa4vb6GVIBSNHokkckjiX4DussnYIpykyGrU9U87V6NpphXKfrkjFi
hmjxneVV4HgHkAcc6p7/lUjc/oTy5Slm8uMXXHfAn1JEAGlr2++B+qQYpmgx12s0
XpiDn8BCgvsCmNeQ5aILPoTwAOF05MW1ko84u38lu9jdjd9mn9Crol8hrKikbr0b
CCdYKh2DJeOJ58eZd/9mZ5Ukkm8zG0x4km30vbLve7hBI3gOrYLjlyz2qyKJmZ4f
0PGrIIejmldBlRLSGZv7N9XDBCoxxvhJTjmGdVYEV+BL8oK6n69yBancHEZLgjGX
i3MTCreZ9LW0Y5ZLIZpON3kxvquXcAsm/q7dpTBcOTXhn3uZJWC4aNpOiSfCoHB3
hZv5ujP6XzUL3ezGuBN3AreZKtFje/dwikjWkCo91I1+zzNeKoESZ0h55du2bzSN
6csuFNv3u9rBYibHiDyDz0QsT2KPFqMB6KAP4ShQF14pxzIqvAVviAs2vl7wk98Y
/g+YPl24nOIwGm4dX+PNu4lHKE2KHpaPYXBf0jWNIeyu9KhEw55IGTTKNb+L9HBl
yrqzrfueU8Xa0ZCvZ1luPzjT8j64haDh7TLnQ6UKGKL/o7VTx0SAr6ZdMTqevOsx
/ACeetocyyBAN+caKH7GJqAwNbKkqR7Uek8X3R6tVIUUbTkqKv3aS/69DVvyfOMr
/Jw2JxetbWnlX8xqjBCPAjfbwCmzjncCOSjlcYKb6nzRqXpPS93F8GmbOo7/yWLm
coS2C17glh5PwUIbiRFOQjaqZ0mv2qXgE+x1d7wozMhjcxWFEbLk6mVRmbHAgzU1
U9TGFK4HdKvaau9xXloPPCMkCCie8Jz1Qv8bour1QPjFLJ7Sdqb7AIxHiVH8Ro9H
GcU9zqRuYKwhDWC4OfPYyd1ZlSPVzyfI99/taILB5nTGFoNgCV31L+y0zTIrFXuV
RzbeM++rz2M4gdf7kfzG/qmABkfxOYBJut+rJFNZyC0G64LeUg8LzErr+RfC3i8w
SeCtGHaQJm+XMxhWUU6t43YCcyaHjZoSzRbiLu+E1b+nhS+Z8n6YOhIovYNkDEYA
oKFlWoYSZ6xYxYBv3EpzpB6Kk2gFMwOldsj1/v3dwC47FRwYifPmJl7fP4uFGdm9
45KO3yqNbb1xQL8hVOCEXeWadBlZIfrCcdu2CzkzfTtZFIB0rvMtiPpQPK0B4byU
Z8ohQ3dTxK3ciODVHcFlDhDwKTpcRml5cBLouIh26Z4XK1xSePuG5tnaYoa/EpJv
JlYP4hQuSliFQkLg8Wfc+5o0O9YACbTY35yC7sZ3rrLDQu5N0STIdCS9kjZg6cW+
XCMNJMFdYtxY5zz1MZ8jz1aDrHzvT7SNvl0cXgetZ7FHFc8s9gn7FqeQnWldhkrK
/Ly1pzO+QK9itu4JbWvfJIv+w2qBUlMIeoe6ML5XtlqQgNPc8HSQlSPUH8vMvFgl
CSMAThLuA8/kJcNfnd2lgLuG/YoRtJs4pDJqmM3zLn7hFsZeGM+N2jSCcwxLUxDI
xKCgE6XPlePUqhia/v5XHyLa0SPh0hrk7KdgP1UQT55C9BTWbmKJDWgvZKjmmULh
XiJlFHX1vwTMncHeVtgx40X0Rta3C5Z4qASbctcwmuqdFg23NDwnTO7/fK6mespa
/pq6/TJPZcAa2ox+oY+3J9s2Vb50H2iWAaT+mOGObt+1CvYkgmERv6E8ooFHsjv4
jf1Ea9pf4ITpZNZ6qyRHxRb4sORgBYJnY2JEFcu7HOPI9yBXBu8JfZTuf9EeESwm
m6TAR1+IAx5t+W/OGYhy9HRCdAnTSOFXEmI7DqaMVv3XzeT4VYeC0/Fo8kjlVvxJ
bMFgEeigCISIBdvvLdDw9aY709WRqjhZAlL2Hqjdjl+nF2oeUrojY736PymPM237
5LW4QZgZnNPpKsw+JrjVsNH0ruZOeMYykPwGmef3Mz4ovuzescU/FwwdtkCRCTCa
5rCTkthpbFrRUmcawd+eB1cXWbAnfddCWXCLH/T8IbPQ5xhv7AhBCgeNv42+E8fm
SJASd8beg8jP6czrippvwgI8v3BhgWuSI4DA6tcVtchrEKVTPRkQIxUMgV6wMDKQ
zMpTylCkJtKz8uquibqRSET0lIeZcMKbVOLlHD9tsF9OeInJXqyFgdmGLt2lHy2X
7u30JpnyryjW3eLAECHwGQeZhZzo1UC27gJ7ABEtdBcFlB6MhJm5LDlKUPD47+hk
teb30xzgbD+qqkNkb4PsEF3E2OjlatVEZZ7hPgc/XGioOxl5e9OH/Q8gpR6zgT8o
nxpEqpgnfZrS6UrRawHGEMhtol81OrNN0Z3D64EI0pHdQsIvQEK+bFoIRt8FXaAM
RxK3O5yYLdlp8kxS6IAdfgkfc0awynxFMkC/b3nlVafziDuJit2hshHHG6IaI8HB
ed7MnJpX0qV8HJwAdKy2a9+xFHC+Fn4dQAPIwg2fWAfJvYB++Dvay8HK7VddfiTj
8pD7J8/iyueyysbGkyd0wMhKgu1Q90IB1HJYa1RK2hIVX6jQIG2e03cNsY22LN0S
zr8RsEkbXCVGHg2Me1Tiy8u/h7bWyhFP0urAqLny9tZe9iiQp+jJT9Fkpw5NjkCL
uTqvbSPBnX6yW1yCH6oj6W2dnWAE45Bal/t3nXsiC7X9wZpsv+M3FFvVMeBNK63L
gw6df6tGql5553uCTawH2rUS+nl8HsbccoDXWCTK7QgUvRxSTUn/0RnwbjmYwIiY
lTtzCnoXYJTxh5gpoI9hBFwIxG5f6dfKrMgrQWLbLJonNl4XbXGXsj/VY4jPGzns
thAHVQ8gyyRE+GHy48qn+Bf1DWxjgga+hB9A8haM0MN4VnZtrjGAo0HaByOhMX8W
YxxkhR/OmfCVDKYXoB/wBag23it/RkaQ3FOtL5OtRI6ihQS99PEBLmjw2tvnPqiP
+xWQ6VzD82qiMv1RsgWww4Y1zEGP7CcRY0aOislUucthYqFSnC4bV2T3qQP5xjPR
5igpLkmWWdcqItWyZF89IsYxYgQOca9Al+sPmwuQixzIRunZiR7IPSn6d3Vzmwzi
EfHqjtHluEQ7fnJnidJ7o71NERRifHgYimOmu50fNrRmksVOn1YdztzyeEFoB9/2
ZNuPJgtdC/hlsBtdfIleVyi5UiMeUhmoqjA4njuyJ6CVGwsj5pP2PtzZduMwdu2E
4W6GaEhCCPkAIxo6vUwE9UYSHRQH/w40pEXncNeU6D6BcwU0xjFoLcmyTtK7GuxR
2oZaK8zOs41N6fXNXyDl7VEzc2NP8/xCajcNgPzjy3hXNsTiVH21kLViaMROQHZV
hChZJgiCHQ5N6cYgj7n2WyuHM5+pakpfjs65zngtcCi7l4qEOrYzSb/m5AUwfhFp
ukW1R6sTDRQJSjTyDJjb+am7D606KAEwmQWvI4ZJuZGBTtb7L6ujTMe/g9O8saa0
ZbiTNJAmJRq2FakaiwHf7EF2Al/0dV8dxsGsBf7jN9H15ZyBaHLf7N7EYYK97V2e
TqKnp3nwWqOfE19nMG6r/uN+rfGt7laSzU2W04nTF+O2Y7DO1R/7lnQzjtX2BwS9
pIYQLt5Cs4AJOHCleLeZEiYwCtsh8Byh3xW6/Gf7fkFpjI03NfSN307tVMokwKf/
x2OdULXWp7GSxv4vQ6g6R8kDQksE6CvYDKjFJSJ2XANiXBwQUfaeHM1ikltoLGsN
lve0lXa/PTv6I0ziaLwbQLEij10f5O1ARde/uXlGVfFUPVfeciVPKWjCREKWC82Q
DtlNpBwnQixA4wKpCDublPVQjNi7A5KJYWuW27NGonvkmwDOiEjefGnMMtle+F84
ikgvX6ndCQaUWC4heQAr11503XhePTpB5852TNhYWTEIvza7xB9s2fO/4BGSFY/e
jpZhA0lcjjf94W6OguPwxgR783D2SYjAPIpbm6IF4KGBhKzhwqElZRXL72/WddQC
ReNbX3HOr+Z2Ef9GXxs76ng0CVL5c7eP1Y4c4U6LkhBKwWwVp5GdTdh2XwEKOvIv
PrM8ZGb+aaPGIltjsZ5lknrz8ZpRc+2RPSe5ptOvsUWcOpsZZ9MnIkkpc3a0vRF7
tyYtbp2Vhf0W/ugDHnsus8U15jebSngJPujIz/oOTPL0f1OJvTKr3xlcrW1VVeNe
rG6fJyf40aQ0jacjdHDLlaM4U14ksjN8X+uVoyIw6yCsB8yI+SrQbLVnYUIfRV5/
PqC06n7iL0kCMdIZNyCX8UmmGhv9ig/vsNIQe1U7ZtT8GsSnX8YbIF7WOmbQSxDR
KLOFNqxB25b8MthRAk2KU9MNwQ9yYCceqJJmMWPqP/VpYXiD0R//wPLEWdZtxzwl
Ag+CAtsUBoonF5xbhO7lcC5TGv4HfQcn/nIrygE5BMrMtGqpVruxfOHBBSQWhn8A
xZGNVUivIGTu5sXXWSM6Qzj6pgP8q3A34mR2ukyavF1n+Lt/MM03Qwt4Q6EF7T6Z
+MJro6Pj/exEkzPt6G6IFAg/nHMrCctmxoqYPoKAn0Bk6FQkF7IYH0AArUjXi4D3
XWoDhXjmAMAGA77RG8cMuquHBGSs+7MCp1GPqLfypkODrxdQx7+fzVtQA//9XbDZ
ebAkYZiWQfTV0TDcvyal3RJFsoOrkWxfgXMz2YXXoDOX3W+AmPusmENZZtFctgat
axcqkNSP9RgWpXwkKulAC/H3qt5eMYgygVZngOARxq8eQ1PoxL/u49nCYePHFfKW
W5QVrjZBTrWZj1aivfBFLufjAyxYneRj5n2ngKpRr/K6OgWlnoOKMe4R/q0nIuYl
n2JJR8Holw+sQ0fYea1ixfIxDPcOOekA+KpmJxorYzndJQs5U4owFRAa7gMgJJsL
S4NtrasduB+zKrOEjiEPM+Xsu7UPhj2hvLLne/tFBoQ2hnrfIpEXyeLqaJxowP8C
zUefxF/D+n1qhaa7qnfv5Efsdb0zOYMKQnmDUaVKO6nYa49Igi0I9YnRUW54cdmT
Y8Agxp+s/yRTZeNAMdE7aw2EXZ4pW+DHEzxBs6/INZrTZb93i4rgMDr/BOH7Ng1h
M5ubWdyI9BncScKZt7RDbt2rYzc6vkCLO3XDlfMqdF/rrtuxMnuD/ozu4DI/uCdZ
v2VCIsJrb0uAIyXThQ+zUEgwqU607GqVNgeNTL9xDr7RvphBv9SdRIUs5sHbuRjG
a7u2JfXsGv5qQqdX2xg6EQfSay5q51FDViPFu98/2hMS1Ki+UTHAHmm/HapsV/pK
CV9zNmu0WGtkNuW29ZEISmm+08dIrX9UPorS+rcqkYx15lTdnCWJFdMzTJIrefcK
NYwDTR9L7Zr1kpq1hjhp79rJuQEJOLSPLo+merPxSF5wF9Oc0LRnBvfwXGco00wQ
6V8J0YXjMJb8dIqdkOkrpciKIJmoPODvPtN2nyVUbR33AFqXGjHE2T44sVtN9/GF
RJcZx3OVpQa4iP8XybGN6CLXED1pdq7UP/a6ujkHCJ5rWSJ1oZuEprIbq7oiL9UY
+lYAtehRIKHKf92KuEIuwX/xoIYJfVMWfyHRso+cfNnQ3tBCq3WPc+PhTcUKQIgD
cNVUCZ4R/hBYL+ieV0XYsgaig3vl5ajgzxLOY0DIGlq0tFGDT5dlI1HPDXWa5h5X
PsgpVjuI9WkfkpUYQsf+5TqT/tpVixh1kpRhIQbC8TdgP7pj6bUtcQ6m/OWsV9iC
M28bIjZ+mabvd+/bQNzR2G5wWd4SF5B4D/TR/xwJM3gtzbh7LXcxFOaWhyO3tltH
PfVJpSFqKBqjvQnYLTX+hpm5xvOmZqyLlmDWdFKZH4ju72oWpP2Ugh0KrF5zPjUt
Yo5q+KTtepvwbpGu6JV5dxOXIzmEXHwM1Ud1CH0m67Wv81W0ynjbJKsFazDb/9bq
6LWUOovpdJ/+FFMUTd7BlaIbw1wrNkbcaRylkE75uv8JdLQRd9vUceDsViUNFlKa
BrC4mZZsjmLgP2+zBRhjomf1ILVvcmz/fl+0rh9/F9eTOIngGKzDuoyDrHkWiECx
PH/iLm7RXmCCuJHcNnVOBJBNrNgIasvym3hLmt1dM5NtYt2nCHEFmiHZRjhj03F/
oTmbKaWJ62XmiX8bYIKvfWZPn1n4ZKqd3hjgzP1XvYOFkQ2HtTxw/pP9gMDIFUI+
1vJC5WtSyFn0XZEq0MZR6nLkkEvktbCQ4g6b6xyYkSlvhhIYr+Ze7hhX++DAtrl3
5fewe8vcMFpciEIof+wvK3NekTtMa1QwPeTSKeSAdItoYy1FoSeYUETs9eRJAE9C
P5OP55wNIaqP7YTEsTLmI3/f41ipZu32ptGs0NHkKgaJ2oJ3z/Vi1adwc14qacBr
fkGhDjhHwGXMX3kQv89HNYBhswMLtK6J36ySPaAbQrJ1onNarXNPN5KuknYn2xp4
X6oRgQQIH3X+Y80y4PBscROACWw8uOcm0298dZGVpUcNfLVhhCvqXLgDMAWjSfYO
kxsXwm6NypePPo9JVgFPtSxqQWsTTK9DqUeC5KXDMIjO1B3KAYUDmf5VRnkCxmPX
T0e81HkepO81xBdaM07pVuxLjugdp3CtYR1LQ11gKcm/w89wJwI/D59vvz/E5DCf
MBfBf2880dXpj58Fao+4n3NRXAK4ksSwCK7Fa1g9srQHiP25M3iRSZprSu3QNY8i
fga+N0RvhxgIEXVNttmz+W+9nKzu/uXVbrRGk6QFsEv0VAZXcsX9nhfbJ8ZdIWGO
FYZJzn2Ej4a2xnBuFU4HrUHJxdVQjt9kMTOyTqTn8X7ebOzHpaHFH58hX7vnt/yI
56rpb7/Y5JBFcqbJdrbVOvlUDbPLvhztpvUfzrj9ecUfRjZmLvlAivVrOP+HB9O4
F4WV9EymphMBuazOYFEFwbGSsAidFihtrGloRNKlV1xjvcOeVR5+0Cs97UVb/BA9
xXZwxPn5hfwCLSb1C6kof0vjzXsgcmqz6iwL6BacdCLd6qKVJ+PmtyfKSX908JGD
jiDx5/remNHvUgaFBXIMx5PrPvCojgYTzJ2kjtLy4Zf1pPYsDlO1zotoCy2xWOSW
cM0gKjW5Ae+1ltag+Q6g7KuDSLHF9AhhSsWgsu+GpKOLLLiiMTPzEjiuHkky1b4M
FvCiHgLr4yOL/KKQQEvssgRhIyw7iDNySobdSUKu4R6+7ZXCyBE9uJqljvZGVBXt
qlNDqUAY+UFgchqyYLkCrbkBIToY8FZWCvT2MtT6gg87wB/9H9Mt7ab0Dzb2Q2I8
ZqBoLzYVVF/Wiq3UJKzDUI9Vt0g92XCsJjmiOLBWL6Dci27CNT2QeCEJsXQAdJr8
Q3qyuGoRFDE2n0XkfCAaDYvmlqyCeuHY2iWHFjRTSlZh5FlhykXKA6gzuXxmWzog
5S3odY9WpXJdCeLlLppU2BibawNmj37aZ3rcmdr3dvn/xzVTE9PIzo8OdA14vDEA
GaeZlyEINoGOUSu7nijJHDxRpmxCYfTGAd1BOwvFxjEystP74wXEzHHvRFV5fZS5
j1ohwExaPbKfJA9ZdadXM6nr4+AJZCFHzg7GnXK9RiL+HHY9PYll+ljQLaa6T7DW
6rnWBeGVKW76J0hVs9k798gqR2tk+cqu1WTLLEzlE9O9Ox1Adwp4sZvVBdzgkXNq
GSEWlEArspJFDXZ1Thz/qVzW7tV2Snn7MXs8kiBS5nlAloH4Z2/B2Q7Nr3rc8uqC
TaQoHIwIL8vZ4NPKBt+WmxTb66vT69Ur+GIAapMzt5sfk6MKmq1wY7BMx+LJ001j
VURlqV6ovQA5H36FpfBbezYPDkQpgSCf1Bxxe/82rNSn/HIEjlBI5L+1M7f4syn2
fMnSnivILAd/701vT45lLd0iog6j9jJsGu096/BE4/70PfKd3+20p0YVMobhGGp/
JWshoOaPPonkRBBWf+NP6tx6Dtl11VR1wASwWxsHvKqz2Q2WemuSTd+wUF36w8mW
2u0h7pU207QexJ9FqQXPOMuy5syDbMjuJVVMAOOGLSpGbpmD9uJwnL/oRNecoMM5
70jcLzLXgZfI4/hR9sz6059g87RCD29HrtGDrLsnF4YXPC8sp5jQP66ihKrNl5HK
slwvHVp2hCMKvA7gb9MUf+igOGhvodM1KGq+VfPNF/+5DXAFouvTRSKHlGZ3OXU+
jSpQCLAL0zgWhHh5kZL/MaETy8GJgBoZop2G13NtLALrpPpLxEEarivxXwPh6Aoq
bg8sx9fiWucfllm7kQl/fUsQzoZq3O4aUIzfO0lKV+74MVRiIIb8RdJrhUPPFeUn
o4v8cVZuEep4E4aZ6SHEYzw3yWNP5FaTZVEsE4GmvMMFe+JIp8XdU+GefkPZ/ZtE
Jh6d+nNftwCDZfoVHQ7OiGH0XG98Bho1FIAWUdhM7cVciRHcxkkGLtqKtQm70ITT
5OVkL8MYoGct3m6oQ1fW0lN0vnjfl1OrPRQaq+td2Pamf8ONd06XVYQzeUGr+aki
fxD0s9YrmKUjOebh6i6ISHyV8kejc1xiWbH6WoqYJUO0pmRuuuKKzZ8ujEVnYo5a
BZGAYr9mYJNc4LL8K7yJoIxpfSXiS1ul5M+HXYduZs9RVSXfobZFrxBrgv13iqfB
5ZHih8+/Lf3ToSkjXG0r21WlsyIVfyx2g2YmHG0fbo1ED/7J6sIOGeAiMWLs6eAS
reyP5uw2kFX5UdB7RSMwri28pOZQPcpaEA/ZOC6KJB2mjl6RePdfn0wCG+lLbPFJ
UcmDYoIAzJUWnO+2uNaZyG44uhiSM0BLUCXoYFr/DA/Gw/lkgYiOILi48vm4uT52
85uqlzURnyb/EJ+8qAZvOauBZjMQO7XIlJFwFVPNmkNyVsrI/BzMdySBnMMlqlh6
lEo62wZ7KcI8twQU+F12ihQlL1MYgHwpGXwwcwLs8M0pB2PJXB4v8A8LW4cFwDYl
767/ZXB7K42P86BuY7tH/9P0xHrnwH68mqpRAFTn6Ployo2YfhK6syUOR1uvHzNq
+gaSQ7BT+WQ/V1MPeiwe6hhauDrkQtZ7KdIqIJNa8BpjsF4aMZo39CV5TEo3C4bT
2IPBPOL6UlREPziJ2I2m4Rab0I3IjtQDD/7phuEQXWHKYfqK8zIxyBDRFnzM079C
owyITPHJ/c6nA/lV/5T7jMTOG7lQd9rNCyb+YLhUFCOEJZG2H0SIH5V+r20jFO0D
pdNYZ0ZLU1cD+wSQdvipkVevvRSo54wG7xHoBdCbSgpOrl2xehxdW75V2sKxVBEN
iGVo93ENZv+LfrN8bQgFiMiD3tqFHTXAlFbaJFuhn36kNv5mBKDzR62o5MKFzR4H
HiyQFu+z0HBLSLFamwWT41spxO9jqfW7mX5c1Lxtoouvy8LvCmCZ/T0xM0R/OqXt
2RqH29ia5baTuwh5B1u7OuJHzFfjqLmCnHw2v7QDO3CEsBKnczQa97SDNv/QxeML
hQH3qEeM2Pqf4yWeVoRjIc9bb0oNNjHMzljpNtzquj/gMaFSCE9+PIcqwZ4RcsMX
cX7cJPC1UsWFX8GtKzRTQkZCu3T9scBb51onKzidsJRQvzG5BfITDt0CulMcO+uY
lK9WBi1WWBIWeHPhroyMEZszX6IrQP0+1ngZKC3Ihp+rdbp/3X5dHYQGHN8fE2qz
uNwdJj0AeEwjNn3TAiJI8DolwUJtEoop3FwOE6xob7YeaJtT9+AS6SU2eKgSV+HW
1F4V8aB6bP6A6sB2Sgc1OarDUZtiij0Ax3BOFc6T7jiWlsZnaoLbr6eykzD2uf5t
ixPdYUfcCO4EOciftnG/hx70IiRDC6pHg/cO3xXKOcPiOxiE7hqfIuanXurGg5QP
pgG0E5mv5HWPzi7DD590FQ0Yq+34VQq+m87AFcOyRk2wg9EPIIJKUTkvRzauLBf/
FfoqHr8XpHs5VTUjcEAQ0eJ8kyvBO7Lfdv+bNtmJZTJE3zYE/mNFZhCLj6khR7B6
D8LG4A3TH4w0Mb9uSl2woB6SRY/QSOp5ypWAg1FVPf9bdMbIYTNmOyrjafzyidz2
yh4xrEdKzrz0fjFiCEV+CFdxtaaJIF36SoPm+f1G1Ql+uXrzQIPX7U3iQ82WoZ0Y
QW4dP8ODIdkuDsyTaKvGGYvxuZzMOG8YKKVTdn0d0KdaWIuueEfNRk0XZcLissnh
EwCyixAT/qClf8vHpnnsQdZj07CAcVh5RuT36y5KXgT0CriI0Tp6c459RcysTmAH
yYapvPTDJCV1BEdjAho/KfYOCnbHxfRByNWDyVnF7iRnY1mRU1vDZbLlcQ5mPkLn
M52C4uJqwpz8m+FZruBzOP+jQbDeW6GOBz6SHsHoNxclfNNLhWqdb+TwuIsuW6iS
+Eeu1YldoayIfj1Gy0UQW/iRG+D672Eh7mCIsuOUyExwBjXV5BqhnuHqn+NE1vEG
KJ/glclUhH9gW/8IVvMuE/51Vj0nndzYJi27PmtzbyvKDG9cpHTlyoMJsy1NUuLR
IqOVCllxsqcR9OzR9A94dU0tksjQZkOHLTIdbQx8D8uyeejdAw4r8QdaSIw0HIP+
oIqiBVfT5/5tAkrS/TdtPKK+vH7VGOTJZyNQvK4Mz33DlsQIufIF4Av+H2BytJbn
AqpxeYOOxr706OfXl8mzG2mPTU5L2bvSv3g/m3Xen2nmVE86rr888m3jAIQSVc8I
I/z+Acn6qK0cx94lTpvMjjV5uCAnYAdpgq9cikO/Y43qgufNsafxh9yceun947J+
pSc4hl36+qwjxpuzhVGexlMsyedInOm1gBRuJdov/XDqxEhXKD7Y9BTQk+SKuy5H
sWkcflFzHy7FfptJuvBAGlei2pD8kzCr8Kqkukksb/opcdkiIACdh7EHLNNswSg4
qGaRa/ys11TOhxt9xtfcZnNktEMQV9f/9Yi9Q7xCtnBWQT1STQWR8uIUENx1pyNF
9uiGDCjIozyOryV27vTN8JrXqxYP2Wj0K4wyKqO+qh22boHg91uy8hyovdi+uJhE
rsna/E7cNW8ymVZlqt7ZofuiCVLO8K+6H3AFdVg4Yg9o41osT6+VOsrPx2Wtl9s1
D+MlLKTMf+bHDjq0AnLmYNSWzUal+zCdZBcqTK9l0nYrmQFnx4w67ywOxj8Q+zoS
LdDDllJb6Zfa8LkBa4twNei2OJiNfOmf2H7QsDGvyQctV0838TCBsKpi2tDvTrIH
sHagJQKyH4T/N5RsukmJG1IOkkGAtxGTqHBpAU4gMMLQOEfneRXVuRZxdB5zzWJ1
0LHvd5Z/EWNflW1z/MwbI5iKCse0GCT+C7fIp476SxgMPyzKOJFsXuBQIXYInCKE
ZtxxutKegAjMbRle9z/3HhikTAK/d0PtQ9Gp2crdvhsXtDJAVcIgQHpHpi3VlzPu
+i9tB0VVI/jXLBf28dHPv0vhxzNPm5jHfT6JuZofHzEoOjv/UIaWTrygN8ox0ypY
oqgIMWYy7whpeNZBATRmDtzoyCvjsmDgOIKJzgpuHtMyMhD25tZ7q0ECaRkWXIvR
hXyUN2dZWU/f+Mh9ey8gRd5EJYifWeGse4s0OsCchukFur/nlS2RFAgyp4D2WnuS
IIKs/6JEHUPIt9WN98JAkAfKee0qBACj/RNG3d75qYdqHOGcsAIrRdcWc9M80PUW
Dor8EIyWrW36gDg6gd5q4djie7dki5UPM1zoN/7rydrGaNZbUQtK4XggqkCooQWC
QA8g1v0Tsgv/7KsO2Q7sAst+SBASjrTkfRXV0mTml0trZeKbJkYqvK0AIF9YSctk
YjKVL1A3+gwUf8iMs/BxYzIXdOwd84KRCjrR2Dh4TKAOMVT4YbLHMVEhGmkLTOYq
+LmEWGOjd7SW0F0/5Gis2ElkzacgVTFbhT0Ad6Lx4EarvWQiNrU49jlwuRrV3XW/
+EuI+pqxWcsccVnZDIjhsRbFA957IQsnw+dmypckTLBnmfpamOQpAnWYvM0we5qk
+cZcFzrZHc7ez0X7/XY1ymhTK/F1ApibYYNfaPn0Qrw9+9AFkev31wgf35IEp/Xl
2rg+riCpKGbLaWB5yU1styqmK3yovf4D3J//ZNj/H+11Dyw4KaTD7FRQpSdG4hfg
Ip0awXkdF/Uft5Q7oFLIqeq1Nry8uT0ksoA3NBoPMJLpfzGO8o4UeMX7Z11GLQsM
em7qfmsUgFa88n5oyHvhczVJsyH8Tjy841dyLBaVx/cnxRFjr8Io1X4mTkoxFdEi
Zvh+dI5JisSJDEdhNVVZNxCCF8wteOP889ze71gLoqfMDcoJ2w01iGZfWCg52E9A
Ius3Pkz6RzDlkWpmeXHU3lA++ZiACeKH5thNt8fBJA7zTkRgGWjNC/Op1ELcTO9a
HaktsroKiVD0F2MTYNhmoeSRh1j/uKeWXh41k49y2lAEs8bsskwgM/SV1g3wRyu9
gk+5oNuz9UdQ28iF+deNH2rJs8OqJiBZ9xmi9pSWGI3ueHh5i+7IOCm9xIbwIJ0K
C0pdWLlzWjPAPuG9Q/CQsMj+/L37kml3u9Eck/0hC2xPRBrp/yGDLx4/RAOy8slt
0e27AYWKZ8pYBVPy/QRs8U2VjhGDsMpALyzJhzyQ7LXZDd7C0jDN2y1gOX6KPwjz
orshiOWfhseSX3jps48uAn2lV8G1OGK38tiqrkgqYuycXr+S86qc2JgonpS9LIhJ
OOFg3OrOz6y/GGCrimp+kMyCqI2+CyRXyLXGY3sSbOLcNfoCEYRnmfZAaKSjqWJp
i4chM2iNd41TuXJsXhxGQWlZpJUSziHeAXxAS2RxTAzOd7g1O8aiR6mIaW3Qdahu
mKpSLPTNAiUacyaJau+aYB0v631YY5dE/wk5znFQT86dCxFoAye2bIoUlnonehz3
AhryeMiWSsycHKO3QL8sBFm40AXSGgwm1Gpos2fNTL4lNatm0lMXT0EXFp2/UGdN
VNtD04Y9Q27fUfdHLvE8cLqbxoHJiuA3yIqfcw+Ixm/8LWmOcW2WoRyr2jfn78It
ePZ9r4Kpw/vDV/FHmT7Tw5QoVBys7+wneI/NBJH/ds4zwE02qms693tk3J0mE3lR
3o1/d+oz05A05o9GvHGGgdXTgaNXnHZ6tr/FO4sX4Spmc5d7fEsl3Arbkhvm47eR
YhzLz27f4NoxwcBo1d1mnnwCwS5WpECwonBHDRIaTHWyRjAZkgx8kh5hZ3yw9R+X
lFg5T5LNQVd2dir8WH5b5ARn/DC7d0VjVlh9gqCsQLNY6gSaLNeQgaRGYYLd+Yiv
kIrV00Eq/u5yP5TfXNX9b9HxJ3kT2BZLT+rXbCgwe9Qk+3Ga3lybR3zaxNtj0gNE
8FUh62oshVGbHuyxlGIK2BQEQ91DFisBijH753r8OZ/WFka057M2pm3oQgDUCGMP
oTY8jHDOpjLey5M8KhJc1VNNml1K7pyfbZdpG9P7/nwuDkg/bNl1p815UfuCKKWK
dhm7BvRTE3uhqI8aUvy+MB7AE8Hs5yeHPT0dBmwI8Unb/dWSpFUIiZ//HAIyCD/K
PgTMUkGcU6XSCdEe+vcgum/DPWDlCAbsFUPIfRZozxx0608hGGRkZqptHzH/GMTz
tWwv0DXZ+FT0nyPmGlsr1tAQDkJLYH7m9oxjLSPelZCdJBhm5BuOTx6bz0w9EC1T
jg/9vKX+mwS86pWz4eMNHBz1+Ql9GB1SVgoeSIYjzHNXSvhs8h29OlaTjckGN67u
m66zp4vXbhFZwavPPadRc+JhOjP8sTiqkF1Bx2QwPKj3TcBrXF5kaqrZtH71uM7v
VLfAL5sHRl0u/4IuKD9PZlsX7K9/VpnaP5BcB7YtWZ/DOUqdyb2fZyNfNRijIQZX
MDqsM22urAywXRxr04YGAG8rInl243FlMIVEqV6wj8wSR5G5+k5GdzxTbhfCWZH4
A6r+aCfnPtT9y5AYh/Crs2/mRmo0a3s8Z4cCP69OLYEGUCULMVWb/Ne7zd8GBPIp
AQ2E8pkWi8OLelo9uCtrBXTKweTLeO2p/LNzMu3Q+A9CoogFCuiWGt3ItIpOu6xx
tzyM53VVbrVf9J9JgZUlgE3nXnrWhkq7Fu+rj1GIMCH+iahVviU3N9SzamQPaKES
sczt+jR6sJbXt8MsZa2JM4klWBMjSuIrKwymacfBtjyNSOu1nhr80MGA8H8X5yiR
cyHxLqo5zyQhzaPIXUkKY4xIopCBUGzWk6ilS1A9hYGBfnMVK/n178nWwj2hpquv
mS8brpZPX0c6ys/6pIcqkLLocWs9UeHuYhUVL3pyKt1ZRPzuF6FoQyltw4RnSoby
LukPwyFw25smo0Q8dHyF/bGZXwtFkzmC4OBjZtLGKLcXMu9qrfkzLTHCDU1MIV07
dVF0EYAQTAGeYCFQAFUKvsrvpfTOglbVRFToJGyIOTq477eUW8zQZnrliUvHQQeR
nch5Em5BVeNxS6UtM/ly7ma9FoIkBrp+rFPl4hibvgb2tYjl8Ahn1wZD+mlXriyu
YkorJ9ErFrXoFAvGnPTUZeo/mArwZZidAgpqUw77Yen9SH1SrqUAXfmj7QtFs4SE
/yTWNTBVOZxOBho9bqTrtnZHp7vtsyc2YbgPYxz+vJsn+VbKe6MKLdTksH3kkjCS
tzOGfOsl4afmCq2kPlUSX7Tp1ex7nEcL/6wFUpI045upxaUIVX1mr0yYXki6Izbq
6TuKOM0OxZrfNSgQLBWjcFEgOmG0XsLHLhd5jH8MC8Lj8UgdxvRnHMGg08rca+Bk
0HDCUvvln8AP+DKhcDsL6/UEcsFxH/kvSmiSwxx0liOcRSx1z39ZAj9dN2+OONHi
LmJTIeIUPG1BrmQpWDYUY6Y71bLkEuroRVmyzFFQoBWeb3bULUGVuIYGLcGuO3yE
jhm53hDatzQQDNvcfqMuvD3RZuXkd1WB9H7PyRAuxKayWVCdlXcdlnZrxMNZGbjG
FG3qQ9eLYSswPgPF4TIJVmOeo/GRAoE2Xajk24N5z95clsT+R+oQz9DiPCol/G4k
d5fwZ1TwHUtfLsoxHAgfXcnW+HI4fAY6gj5WXSXPekY3mtgSd5Z8yH0xRy4IcR/W
X/yWkLr9QTk6HSywHvSD36VJN+SJpoNc9M8csYiJTLoQVFZBAnmBwHQR2W0grrYp
DMhsUijw6VaZs8FtMYxUH0gv4qripZ3LIBGsxdjtlYKVjMRjZNJ8aoD1RdO/z2XD
0RleJbsLE0bRL8epLZSuEQ/SaVssTNiLOA3fn0cdD48PPq67NQ2LNZSAKiDmiRcW
UxErOqaBBA0xiLjbmoG4s+LJ7NLRptghjPmTwuQFZe3GHEz68co7c67MQUv4Dhsl
Iu6o8CKl8+F0mtrNSd9jc+o6kseirPIyGupZGa086pk9eGjQJim0ZEoILmdz+oZj
xfWWUhEDCYYfJZeDgjG0knumXB93vQthjCeaqlanr31JAV6kfsZN9vY/w8t660vD
adFZlwWcpCw+5HHXw7CI19s04tk/6BLySFOrSWhPbdefRM29uoL6InPfVS9v8UYa
khl8wiSH8H+cl8lAeOPmqtmkYqdj36T18orK3/u8vO0UmJKIGKKaGQoREXDlJfKR
88jkauZa/iQOqKpKDGyvnTVRXSZtslgrQM9iX3hTkaqMI/sJp66f9B9XdvMkfUI/
4tRBLRkCYqSQVAvy2/6YDxE9zjyE1I2NJ/NIMN3bWtEEHSfdyYKXjubmvBt6lnsV
YF/8PBXoNHdWbOBqIApIWNfn5MAVu072JAU1O+hMpOJFxzgTXKfPZdOW1KdRhyzo
O34q9neNnOLmxPlzTAb6xiqIQZ0/ebvbtQdg/FDLEvoXZwZXGym5j797H8/yAikd
5A1BtPK3xRUEYNZAnGeOgY8I+y7kDBe7xpV47XUrW+9MA/RTvIsE2AZCU8InsVw6
Npvmf/23YL2IzOL+W1z4q+D1Umrdilb3VQURV3Uw56F7E3QSESoiXA3BEtN9qTmq
yS+O13FmZySMhpKVmVhSByoGy9KEt1um/de2Amkskxfa0v4duzkiUk0lD86VqMRN
W7RHDmbiGl8gbJf6RgqpH49/Z6RaPXHhlHc2Rx0vdS5ApREtHcqQU3Pgm4CSoXwv
XCFacmFIn2s13WZpGug/gQk90ThYwSzSUD4+D9yI+Cr60I7hsbcthWP/Fep/qqLP
wNzyWDMv//Qu97FZja4RU+h4LOGqx2zS54hIfLYybjAeTjlTkgpSHAE+jABY7xUH
tedG08nnLWKGYHoUI8gX/otKU5sqGTC/sGuUwvwsdoZQKuvl0qPtLIkj3BjJx2Lz
/UxJUr3Jd6RXL48SsDU7JYZcPzMqwIlBX/bw+MXsZ+hPUe796d48obO9THgV1X8/
JJygM4ue05zUI1+PXClTLUs1WlC0VpuPHgahnLpPovAooy0RcnTCyBb1JMf2u6mM
x69RI4M3NwclWq8sRXFjl9XcbFsAnDUCjyGD9LvrKrL9ZyssOlCQkACY4xScsR9v
vUVC5ScQKLEktjLA3Tqf9EA6XWhzHK4U3CJAMV8NJBgEpfw5zKrDaC12cwXK8hfG
iSW/MATrc1/j5746HZefUB1gfkr6WnILB2wm3STmCSTcp036tmJeeOTQXi4rCEvn
ca9XXS7pTOWeiRtXbjVuK5+QH08+742a1LnWTzcTzhU68Wxh9tJkJXOMYjEaICtg
j6MujE0ax/3fp9iRYUZW67fGschAzT4gQawnkTx/V7vvnDZUUyjsgWddD8GOk6Se
wm30tJ3b/8DP6+fcflhzfTcQuhgHAacvI7zKaWIKvcnzClM+CnIHluuEr5H/FFcv
JwnTMIGzBpFQ01nR+PzSdO5EZqFzK5uO9h7/CpeDeY7adio5I0bwHxfbBT1J/vDp
+apD42wjbjmU2HwANsYlkZH4G56ZEaLzg2jYmuUmRYIoCCJV3E06OLTGPVW0JqEV
0Gk1DUYQfzU9YujkI/m3obJ8AmPZGZbFhfNFMIIEIiuHu6wvQIQpAZC8Yvgeic1l
2rsZzHJn4nk2/ei/Z7OHqGhwV6zVLAm6mx9v0oNBpx+kitjPWhhkPnwgydUEQr5Z
vOES1kRdvLIZtX0QXti+J4AQ3b8bEsZdeUB3LbxrGI+Mip2LhNCa26VepKeRVJf2
+t/XiwmqaxeCLoCRsYlG8yABcj71o/kW/ODWyTz1Ff5pukMja0x2MaEdmBd8xZiN
ACOUGKR8FhgmcP/gdKkho4qHAgvmYOpjxvWTafwHlk1OE8ev0cWgqU+tBXSpSYD+
EHxbskxQG5iKKABxMMRbdCpcFhggExEN7DOInTn7T63nYL4aiZPlLaFX7lL9rCzQ
nw+R7ubu5j5Lp2QEgps3IQcuzgvDJ+2U1T6o2G8SJnQGl7DUvBWFWfB/k4RAegLr
ClHWfO5W4+h/+O5Os1TLI3S3e8Z1xiox31v0ZzQvuFH1OAVZGxGUnZiCDyQrcR5E
4QuxYXh3MmobfHcsQH86IFyBpKqqDGAJxbOuKYmAVK7JCz+URAi+R1ABUSQJ1qgp
UFVLxtBxukuD6fvZ7WTnz5XA9WcuiCYXrPAONfGSi+Jdz5cL240oHgyucGVNQPAL
L2Fbn0GMk39J624ESGjwXuAsiVsXgdYdHAJSVv6oYcqq8bxMdPhEUJZAWElmYZRm
kWWOfjaiANCIT7IicV+jKrw60NT4TdfQwW/4tJU46RaoK82SOSF0Gjtfhk2fBf76
PX0tkBAJReJQz2KqsRP735cktMTpaSAMSaEPjnGL1MhcCPfhf1BhRz5IxeKVC00q
UurBbMcAfjDMV0k9v+ARGU3ZXSkpHdRXqhfhhsQem/hBkBv1ehmrvcTjUYqsn+0v
9MjGNNDImKFWC/QLCCqpdO0NTRJlmViL+F2hv8waX5860YtP2fZQW4yaiA3Sjm0d
6vYwTek0C0YNaOwPYgDC6EFKB2X9rge0GKPa+rrZyo9zdE42sViwfGIj6D0RmgAc
z3LPlsHvJlBg0ONwqDcTJRDnHPgXxkOwGwul/k+nduV5dbGfC2+5vzU/yECDJyC3
3yNV3Yx4z2SsCyN+r8gMT9npFC9mHO2G7p0EcN8NQTuFPxcrDw6Kn9uoX881mfOI
VWl9TcuoBXSOntVKopbjlOQ2FaAim13hqK2C9Pir8NMaTlT3iIWwCLCShYJY4mdl
GyCAKzGR9Y5//IgE+Qa7gJ2XisUvYiBS/jSBGC75HqBbbMvR771RlgWZnKtOLX+B
QJjP3dAXZ/sPhA/RF8pKFgk6OacKKDUsZPGcntRt+feMFodgOxGlquYKBXDMe79L
Z5r1cMMxHJJaT1BUBlLx0kgDEIY0EwbGWhP27fGJffrnt5wtnAtXdVFeuNTfl34b
jXhdILI74S+l33sq2GOfH8R6O/XpD2SIVEtCOCQEBR4fRmU8b1QnYjtU0jgChu7o
pwVTFd/4lLR1ElL4/KZrDEf+oaMtlkHOB+FlI1WqI7knRrk4UAFHyh6bofbd5w1m
FZSqrDYON3wn3ek0BzNVJQ00uVlJRyvCwmN3GCFeO8tdE7Az37ksyGUYl3fy3rnw
iubE6TNnCryyITnODAH5KAd0ZP8R8cvJ6/dlST2l+aLxcpOPonEXeEygFgPaBYHj
BWFJ6ANZTckUhv7spHhxJBwwVtJQfUhXiu6Mx18P065MMUQgFdAqgkZVewsiosKV
JXqLNPLL8RS5q1NL8v0pKaltJAxppuzrl0+pOnxN7rjal3iLwCwyWOBlN8uBXqxL
eatdKyXukRnhgMfA99Zy/WFEBNlJL0LuDIuIu6NFIO+KC4nVjWQCH+m72JSOFbik
gzrjGtu3egVvVv46FDK+pwiCSraUHlBnyVrGglhWAZoq1IYc2wd/y9eh3VDOwRCK
5HPSwTIdBErOcASrCBoeitcC8I6TWAEhcEGIqdhBtjxk6Yaw68HNxpLD9HTSb4AQ
9z8bgphek5Ks+UR4wrp169oW4gsGjuQLzfleitrldCOOgOoI/LVv28LhDEqF/k69
uAVq7/Qi96EMpvLO2kVSzLwK9/HijILV4VRRRqo//tusiVu/QmDEL63b3k228WbB
qyWSwtsOFymBPpou5c63MhyUbrfvODUDhlVP6IeHsT5sI06vTniMzSPNC93ZpeL+
lhKsp7qRA+ou7lN/M1ph/u8AucxENJcDPdxAw181o6Cqi+PR2uDXw2GilfKgfqMe
MuykqCxEDL6FQ4owYaKz1Y2my6MxJgQmTxBU1Fsnhhh5bP0k3idaVcaLYNf2AIRW
rjaJ1uPw8S38F3kuk/OkPZSeTHGWrBQGqAtg6v98N+nhUb44cyTw+gwJxZ7jVqzz
Uu3atPlzlaP8beRWznkoT7yrt7XSTLUKzRL1PjqnIUV8dJmgeEnaZ8u5c5kEmnil
0gKAlrop1IDcmyUBGbeBh5fFAZcXuJohLnA+EqpBJClxQL2mqHvFUQD8Or405X3Y
uwAcQ8KqcAb1gPrDUhL5fyuSwNu/qsBGaPM5pgTJ2orYW8/jD17tQh08A1GSx6Rr
TnDdP+nFtorkGcUKb5QMPEVGlmY7rbzP2h/fnj1RWlgPfCt5JmRTalYpwg4G1HGo
NAVRmVBzkjmP8LHY2adSxM9syFt9xNiz44c4jYv7ixARHwAbg3pNUA9XcTY+IC9R
GlFqA4SZ1Mw/TsU7eoigP+2BnzWDQb7/mQ1G5VCuJTaVkoh2gxdd+SakBgaZDmWh
3B/UFzI4h8lX1FtexWLbTbxII/S8aLEcPiR3x+FNnnEE5NK4juMPjXXO4pwMRdHV
rmlBcokMCkF/WbicoztT8EGjii9ByHdfqVjC3LytYoRZyYn2bB0OhC41oQqCnnQU
TBWeA7bdF+q7WuLjFnzGMHRXctdGa4uLb6XJvNheshQo3yI6IHUPDTzeRb5Tfgfp
SKYdPjtbgJwsl3PlorU0kTCya6umie9PtqBo++y0cGaJ5rE/N2NSbFYp2fGkh6Mm
Ovz8zzOyoCC6PIkgBlrh+RlOnmSy5Cjgw1Y/mJ7DVmg5rkYMvrWNBC2QA0qInwJk
I/vGdijijDQL8jCMwN3Ik8GO27MFqbyNrd/pUBnLvhKkePD1V+p0cG+MqCYNo1Om
bdlmjgxTZqLwLIZL9iOdTmmAlIrAUBZquE90pkfeBbjmxxmYF4lIYPBuW7qyNpM6
HvNFxVicSI6uMlTfM0+lrG6ZnbrWHpyFHp4Y/oMFj0lg5UuK1LP+BoPrx6uYjuRu
4y+9EG8GMp3GsVzKE5EGcvLyUoBSWMEZ7vwWsolV7RAMcGZwFPoKoaFKGOQI3r5o
fHz6YNRn2WFzCR26b56DquRnt7JI/YifRoDe2Yx8UdfmTfa4Pu7h4LAbpPXNWGif
EQP009j7ivX4cCpdg8nFBlwwDv6gdhXu978NmB540dfv+mxVBn5moaUuJsIVp9cf
W3IZPCMBGlX1vDCyz0kSV9rAP8sdk/lqYjpqs0jupnmXs8Cy9jJ/hHenM6ncpKHi
8g7XJbIqOCopSNQI4u2DXxXG+VvameDc4/xnrJf8vnBM3dztDVIoPUxitCpK5C48
2+DJktTr3q/C5+Rx08yxSvGf67hPW1JwE/Yv9KMPM4kclfF8qigxRhwh6G4HDjBw
ecvFG04LeBiUiFLdYrAUhyntllJjiXo/RHHYYz14uZpgqxJzXQlzR1b8YXDyrEUA
KwItNeGX2mVRai+e+Jryts/RZttbtjsWvxixqVmUzJcSaxRs+D3M6CTLv3BxUlAU
vgPA/UaAeD1ryXDokn7Kx6Hvgmmw0Ug5dmHVDDEuGx6IDZGR9OKQ/OxhhBEFlxei
fYhSO0/iQ4iXWlUC/rdomLkB5muAd/6SqtY9X6OM4UL7K2TvbQcgun4nVRcCClE6
zW8Jxm/2DgLb6uz91gWXa8bzIKehzxSt30utp92FeuEJkL5iB8oeFw9Ak7ESByAA
bSCP55ZRowIn89rJ9m70wHS/Jl28a1zZ/pfeVHzIqTmC3pRFj/KUI52V1h648ihk
O6U+u4kNl2u1a7F6CEBGg08qYZx+JkKwgua/Lc4FSGt8xp7w2mP7d4acSTs/skAf
rCkqFNT6cCQkz/qQQPaD+DkGH2g42v3f1P02ycXf/IHXbqJq06zoCwTfa71t/Jov
NyVqDMBEzFUhDYuEuS3UlW3j666fOuV+u1KzsrxL2zmR2pEahFEkWgordtSHA7k5
Zc8IzeAolkRGjj8YDdSq2Ixal/mqA1Prr6Csw/rbValqqTWpRRW0Qe4k/BVPTFy+
fG/oXzxydbQDeq6gWM+N0qkf4NddNS8Pi2XENX6O9HJp9USIRG+QJljx1iAUydfZ
F9gvLMhsQCNctGT+CZJgtHZO8JMSryFevtxjllJHt4E3X54+dJ3NoZ9TciWWt7Xi
qHVfXecUrcYgXaC4/pr7lxb25Goa7EO49wahIcIrmBRv0mxG/Vuk3iebYtb6W9QF
T8mL22QzaiNVyUsAxynXKWvri5RuFzlk1fvyHcoy5nBj6QfujYXkiMlk09m7WehB
yGJbvBzcb0fSA7FjQvMIXPJJ9s5R6nr8OVavvvG5GHr13Rw2AvQDvm2yUpAYPZa1
5vx5Uo7phjTbW/9ru16+p7N0cgdPFj79nmhyCYaUJJIgJWXglsX0rA75z7m+qKcP
bilDet3aiVi9iliZUYBs66UL7voPtgX8oPsGBVesQ17wshJdLn4DO2SaJGEcS+RP
avzRpxTUAgDUPrAuhIMw7lKnEYsr3Cjs4Zsdeeh0x4lj40vqWvquqGzxEYNfyQ/L
uR+bHD0+RzHlNeSuWWGR4sEyIVPF88NbE7954SJA+FlJnx4UCPoDsNfAK3YwKqJq
MG0vE7wsVcO0TT2FL/0zjx8ncFk9XfFZftiQCtbPFfaFLkwhbZMRDfvxs+XGTSPP
70Fk5YyUchtE3O/PXfwlF/UEpy8qZmcDBSvOQBam5Li5Wa2yLoncHnx2JneywCFt
A09xPKR6oXJK8qkxOCvedlQCdB8dckojZZ0wcTlFLvxZkA8TbXY/aMD4N05YNPy4
m0kCBhdX52ra5H71GdTGdurj3d0xgFP/iZg0BOC6Ey/UD49Vfygnem0OnLREhxUX
4xcTbbu2RBKUx14mz5bBkviDx+OVwSJx/PaJ+Sf3883wZAeRNc/oNjb9n+8c8RIL
drKvX7uVbWROiTewikXl1R9aQJ4sfKwGoHd507ljN/pneImlGkMTmRS2P4Udc+4d
46wDgn2wo0xk9JaVf9nsBjHYuXMWZDJrw9KoEh6QiD59v7EZDe3Usx0C/j/URcVr
+7KXqrumf6UOxwovlD+WaysgNAv/4iI99rOXMgA2dHJ3Zcp7+FF7S2tmT5r0KanE
`pragma protect end_protected
