// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:35:06 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EDQAg9Kh0KVbOv3rz5pbQwrQYcXRc8jJnrBuKO8wEF1Zh4klxb31iXrhRLopo7sj
qwTI+zdYkOqWgrkJaXnsG9WcrOWxXDl6x+tjruxuQDWtf+2EB5TOwOE28qKEXD/M
42IbCm+Of9BZx9CeYmQaGeH9JytcUHhajIAROdXQqEk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22672)
RtxgsvdBeCcIZdHYwEHnHTTSKGndih1D4p9X1t1kAo/G5/nNoDkqgRYePCHhZYrl
kuBCEz/VUIOOKho7uFlN+rO6oW2jA/bKO63AhJpJqSJew/INuQ/rrdDIrNyNYovn
pwMXNx5gWkRPdjHyJjsLotvoT651LMAtuaxYCnzAdiAFV5qL4A6Hki1YgMaEsjuk
VqCKBGwCunRjtxgxXWERv43egiSPZJb+40qgAYHbnne9rWxOUa4U2+FSIe1b58IL
WO6xb/XdvbKWIXx1EqwjBo3N9xB50itX/1BNAZ+HH5NpkBK5UOqL/LGuKBlvMN2B
B+wdsXZM6cMu3A60j9rW6T7v0cDZcuS/nkKooVLa7CdWcdxS1ObvcEjaB8A1rghU
2bFKiRibW6o5tbGv3fCauBmck6c8YFmpmXVKrSaf9UD2XDI4hhuBvwk7gA1aGxsI
fYImVHVTJgqsXdiravdDMq8XIEOhjTGKYnYcWG7UttahbwNsozXCAF0mXhOYsxgl
wYQtb9Lpps/4zOxV6BOpWZjJwAuInOVAcwciTI2FRzd0XJ/xtvp2VPmAfSyFRmCc
niBBJci0j9QU9BaIbyR1F+4ujrkhhwwwIkDahT/q0bJSAwrP4PL5AiCy+cdVgvmi
xOW8+2GEiBQjkoxUD2ll7yosn5ux640OJ83VyPUv4PDfwUHMcmHQIiYHWBubFCn6
4mVxmkd1h1R1R8bRjQ7OzSyLgN83kgKdXrWWeCxk+UqHc5fPZMuO9mSunMPgawSH
Dmb1bDQVsiJKeuML+lFXISc1xAeDSDlEX57DL5SJJsoAjyFssuzDq7TmzRIktMx9
eBnKAkuZP23303PpoMWGjjMUbU3/xX8wDfNG9PXQ1TAlSLLCM1ikWA39znHnTFOr
2hnD5MD9vGje5gWXy5NXZzsKwp7ZO5n4OjboWycglEasYdNxqF7t12kfJVsssaRJ
vpJBBHUcKLSYxgMjtpPV9Dq/OSq9UdFbpQaZXGS3zEHccZjaAn9Q26babliKGRc3
yE9MPcW6z6F95WSoDFMulqiwj4zFcg6oKlScmruYD4/ADzs6RJ7RgQYTXVAXnMwM
Zu7uEGDQSbz3XZNaXQYYMNOCXOCT31K1HWS+q4+1inTTx6ZIn0XyNU5v0SO8Ugi1
Y5jF8pR5jDVQ4WV1Bnny8JVShRht4uUMSAmDRWuSLwDEn0qLJXeXF5iWu+67WLgh
26Bo9sLCTRXDaFOpL5lnmkqPNHAljswy73XyUsIfZomcA2HTaGFklzcaHu+Vglka
ZwDZNnZDYbMw/9C4WvkvEPkTFfKCAqEW8INJrncnlHQpM8LQb80N5wcgnLzo0Av5
fFgnucTaVXiHxKhaeu8bnzdh0SwIHtgI7eFWEO6+MxAx10vUIO6ZYSs3fF4grVNj
KlEpb4eT4ZLdKNMd7M3t2rQHaxKcgiIeU57vuwAAqAStQe1XKv8IqvO81g/UDibk
2jXhaPXxzdSqLyqANQbkX6lUF5z/unks0Gsz7eSIZc1peFWFSiEeau6Z7MC6eiJ0
GVclkXJZ68cNB6pLgqRu3MtoeXS83qFFWt5cjY6MCoqSo7YQaKYuknlZUiQvZqAU
xWXm6UeXLt0AqANETSlutxjsYDjGudwQBo2og+4wh5dvL3q+adZLayoyGVFFgIf7
53P6COwlpyyPTXrZzquNkwHMZ6p7j1F3EcLkes+8GrBPL9iOeUvAbFz661ILOzoj
a9BaXuzVxK0V1t9GczUcetzraacruLJKtegh8Y5S+pDnIhwvbbj1qZyGm40mzUV1
pBum5F3dbT7nGsnKHW2BP3sbCKHuKpj/V4HyIxNPqWp6gK9HZIVKd68pTBNSVyEf
M7pF52AWu/2TL5Q08ynJXTFm52IAhPDB7htks12jnOgZJ3xKetM7MjyEazBzJwuS
bC3D3WEguA6YCOFmuQgM8y/Bk4RR2GmRMG7Ando5MPed2RN8P/vWmCsEotq4Lcsi
L0KWMjndcKISrjh/KmLplRQoLmzOVahhtwVzks6pw2o6VKJmms+U7ery74w20tLa
qmqA4j54GFmNG1vMCiHp2rSkKBO0IrImlBDsy0MDu9UTXNILpwz3EobmfmtssVBe
S9Q9ix+4o+rU+bgI+o2qrGU/pxQ/TX8Rb8JN+SPbsN8LsSmTLHU6NrKNS05LpjVA
o/yZu5FNpu0IhTXONb8zSjjD6Dr613WU00HS6yZ2BDloXDpa6jiK2658f39a78cG
6Gixw6DFzybblFaitJu5vlC8hdZl2/WA41uJTasu6l/jQ4c65TrtWRGO2+FDVk8C
vciElQoEBeIOQhFgV93QRpyFCgaQNYElIZ4cHCb2hH4rO2+/j3y3/wYFmP/U7gaV
l5t9oo4pO8X6+jjP6ThEGZujzTB7zoQ6OY7UvIN8vmkxjjAbN7cc7PN3MvxGzEYp
7C37Yro2PlBihE16a6oQ3J0A1LPs25gYLIXu/QkmbNCZL6Ct1uCw6zeLzDeZK/1a
hw4gfI1DR9ZkoGj33+VbqOhItWFkeKyP5uqrJZevNeMToCZkJkvAiv+uTWzevKzI
aPZKDw+S3AIsjgmv+35sBJt0IMbkbAqzwkoI7qgk1az2Uus/46JlGd21tLPok/p9
NCWjV1SabuNQjrS/H48fvDSYhOFTmuU2CA2mP9O+PGyxzjLEnHSwVnjNN6hRtAyn
vkIhpUO5FL94a3i+kpK2T71WAdsZ4z4GvFZxPxEFQwK6gmvQNJFVfZJcaGsZ+wCd
WjXmXqiRNq87t/XGdbQ4LrjhMT6+F96ZBUxpVZ9JaUOFmdMhO49zXzcxkleh2UmG
vDuAAsH+kxJanOP/1bmVBjv7Japjahy1kBPK2Q5PB1is5ZowXP2sSGCP5pEm2swz
Oce5GDB1Pm3Lzccg1R9nQ1c7g9c/08c2oN6fYvh80vh0wqkxfXGKvTcdJl3MdIUN
Cpxj2pEyaqdMPcbwaJy9yuj8Pkjj1pKMC5WhmSSL0apLNXF6HNOul+7mZnqaVUu1
3RBVEj3rIHt34euz1tgcmFcULLnigMH8V+CYyfu9FsLH/H8NincQa/eXyJy6XGm8
g+ujlxOhZFrsXEb4TXVsRHAn0jDpeyppksTQAqAvpFLDlI6YUlcy7DcoC5uoW8+V
/Jiz6CtzgJLtcwJ5JaOd8xGwjzOTYu37S5QfqBZMDx3hZNnXESYLulYzSxaO8PwO
YQEBR2ckdKmaXxrinGa9zSaoxp93di44KjKhJETo6eIq/H2esWGIbJLKHTfzPSUR
1wHujWg81xkA6KacVhCIXL3eQzWgbWEMEUecH6VYbbGUgEZ7BaIteogWtaO9Ihal
Zmnx2Zp/V6E4VsxHDPu+ec6DGw9+aB+0KNixknD1Q4jACjiBdZjtM5K5rSsrNiAD
LBDHccTFKr9BtGnjiQ8FHuIx6E1ym5++HRpDS3+bX96N+zO0PFM8jSPWukS4Pcdd
IQjYE6LV6qc/p95IUNec+e28SOryGNgClTt9ktfhAFBLrd6lPoNHBLZif47NIxld
VtXHuCAveB8yFW1zwoIoAQU+Cn6wsXqPrIZKrgO6rmJQAilxDVx6K4pWtMdeEhaJ
MXl7MRRgT9etnpkHTAy6wErQqBdTOftdKOuRNuNK8fg3AKJutLOatzsHzDnMivyE
D85vPLOCjZ5Xowgc8wP0dOYPSRYECutBJAycyspnS70tretzrTAvnL4C7mF54Qj+
uc5h3eAcuwUXszPse83e6iMnZmaKU1fD+Zt+WrjVvA5UKWdP5fzX4+FIx4rNXTe0
hBqNFReoJHFNt2gctbxE5rArVRtbw0+Hj/i68hOp2GhbQ26DspYs7HwO4W9zpStI
u8BzeLJ9bchGMoPXv17jXmM3PJm+e6CiCwZnCvAjyMf/8ZjVgifUq6g6K89KHKZ9
eIJhrugCZp3N1WYG9CFrX3dWpLQKCXOFY30N+8w7hq4pI0sxeOXfrLmkzsWwsjK1
wd1hmActDrMlfxjRMUx2Vf8vFrs3DZ6CrdQuSgV9K/k3DouhbT0S5gPcGTcXSO8H
P+cxm3VJ9R17nOWP+eVL7HfQ+YRJ7ZxWDX8a0AZmbBomVR1FH9Ft3YNuebzCcFLR
t52HRP0As2bCZMmk/Gl877D0FFgTjCXpffMHwHwRoWP/lNQriwIX8SGLfQe+1gHk
sJ9VkMm284C8cZRJvcH0wQ3K/Cx1oujUwdoB4NH8Gj6+z/WUu7U8m4CjcBqa25Z+
X7XJo08oPD9E6vBJNQXqojbT8AWwCVgly5BHZysMemsWm6D88StWlwskOAdh+G6e
RRxQq0VMM+nX0254BBRUWX63eMqOXEogI1nkhS0pC+BQWrnHEvov0/gumrUxLoQn
5OvVDCw97wve151YIPnlMofFyTBF5N9t4cDn/EHx0g3MhM4fXY0bKCkC9V1VV8/f
mQjNlmlh7s4QZOZPICZDlR+kbwt63zXbensS+fP2eQFAudfmoDzO0LkUhxfEcuu7
mdRpMXLbWr+H8w2AuINrLkPzZCRKo4HPt8jySuVwX5ikA83jvOMS023jOmpS6Lhp
6UfR9q3fb7LSYlkyPh0FC77FlCKH8Z9owL02S549al90qmV7kAA0WUhVZNlqJWDu
3gXWRjGD5WF58xmzHS9puyWd3CfF/sd/lgKDahapvtyNJyb4xbALQCHdaCe0SPll
9baLZ51twNWF+/rT7RuNfA1E2Pxgl/0GJuaj9OCfFyZhf0M2tMTMp1DVOsDkf/UG
LmJdbqBAhy68ydpAhkbBzTNtC87mavotJVScDI5/eDImhHpeWuOhjxxNPpVfz3iL
erswcbV8EoDzIJrFBpvNz5gqnr7+GG4R5dZX4Qt49RWvVvs1B5OM+jepfgQQlcYy
jBO0pe6QtPeR4AXglQRNfEuxeEU/kr9J4eQqBZc8nZB1nTs4vKQsqs+T28tvR2n3
TzjfSe4SWJIasGLlgd1/ADF+UxP9dIh+YfhUQs0pJ6SvPIcvh7FQakopAUF7SKLy
gxtyU+ntn8693ABzlXEbqinXsAXQ2NJnR5AqaFKakxmFT/MjSwd7k7PGnbZT0O7E
9HgUAROw0wJQpr9jerkBTXa3Nnpw35qB0qxRTtQV0Y3YsZ9lHIo0YhokwodWSy/Z
y5483IUfzbPW78GB6u8DBSDvJasxGorSEAmsVN7ccxJewzPSZI1A4oDNpiAT4qnu
H+GXRTvdH+cjv1BNGJ0ZuGYZVYJVOIvy2tHpFI99Sd2T4KndtYgO6yhes0e5l14Q
T322kxZYpg0Cjpgp52um1C99ASI4r+06EXM3XGtCt4XCx9E7DgXkHg/EI3hlC896
WZ7pDaL4owY4ZYbbBIqsqLBCa2t2/nqynbwpQ28DpAzx0PFyMIPR00A9Ewrrqze/
ZHTsJYTK5A9BP2W2xN/eSwNJh8iOnnrLmkSJUl3x8za9ZmzZLNwO3YirdnqdHtmC
AgSLoSWNgbyOnA5Leke4f/6F6ofheYBYdzFpMAWZBRQ9GxUAOR1F+o5pJgo48LGH
/+LAiI8M3vnqwY3nCC8FhggYatv/cpjDxXt4/DJnL1kbkFjL9Bm+o9OTNMMAGK+X
Cb8OtOs49adOduNoifqbU+19Skv+R2PwkcuZGH0MWic2VHROA+wNaWImCSK9WSi0
J9VFUyyz+DpKCI0emRn2Biwu+ZITJxpLfWHhQVZDb1bEjSAgEUUmKEWg+qoGTvaB
If+YxUZCGIcporwZSdXSe/KdwsBUzluNGAB+TTvBxEkYbOXfF7TyjpAv7XVOlGMm
pxvzs3AohtrVZKGwzgiMF+QwK7wtCk2ylrFGGGPAljnt7SEsl7j8wMuHc50eS4QU
2wzouoVXhwmzK9GUHlQATYmiaRrSIma6sfROSdcu+eJm2W5aX5xnLz5P7JT9YQOC
T/OsU+EQzMD7qXtNaiQMUjoKlKphrYdTfAZgBdwOQE61CwhWXK8PeS+Ffoqwwb2/
yeoZukr+wippOWc90ExIvHdzb/VsrkuT2OZ64gWBLhQ9y3PoZ1369HXEPdyv4QKE
xl7rvbHpXTdM+8xxbd7pT3wOn82nAh5SrxPSrw1dKkGnQ1i6mNIY21mOuXHtFljz
ypHXEB+KobSBexEYK20FJVN7l4JPnALCm89wlBUtk5KKylmejcStKP6c6oLKMJUA
b5ArYguUeYS7tqaUfMilx+OICWsBXGjzrMeJsJajiu/jEUbEgLIgTIBjlgN3N6n0
jfVdX6YtI7UAKBSXOWMwFbAC/3U951MrcAVgfI0aFriItT8r0ZaGgECB9xjpJD52
DgHzTg8FF6k4qOfOs9Cx/CiWX+HquRej/tOD7p2jCcETml30t4RRekKLGiR0LTy5
Of7yNuXU6URObrwCycRby9fS87MVgwP+D1w3EQaVnXCnZol9aPYpDF+mSQobCvTg
d46tm+szaAzS0VaUxVwsOddz+xjzWD4WbbIDHRlnbqD8IubmzoEU+cKhjjx/9ejb
wewbnf8dYZ6ZJJxiCNFDrbg5+a1XZEu5sySxkbg8tXJ3gUYPlehr9zn/gqE8bwcH
8BPLket6g/7VjJ16gxoE2+p3Fng2Bveg2vsOZIDw5RUwDp33dtozSeYzoAyI17aX
O9Oh4NlFHAKiZeyiQTdnp2RF32zs7kqCyXsEwpSATvqeFd6mBRI9NEaRS3CECzvy
ezrorDW9+upgFLMHcO6ltmOFjWAWynpxLzA/kUOJhYcsDE0mBS1sLZtRtySaW6eO
QoU1GQehfvjThkYM2Nd2X+OcbSDuj9lcDwnzJa2K8Slu3TVlARyQeSvV19mjfe+/
0t7YPuDqqICDJZF/uTS4s3Tj73MvHht4axNiMltErFsr4rD70LD7lwpy60g5zVw/
1gL+yaFfDmAB6jcTQNUH3PbaAdzXOZJaik73SI8NE3aDlegO8TtesCZeFHaRC9J1
B7v9avjoECAP2bklFovbFLa3TGmg9dXttM+YnHzBoPayE7B2n4nMzAPzfvHdUh7F
ZLLMYhlF7UMPD4uKaDcr4u9Pcvj1zN2LM6O49BBfGpqoQUn8ipbpoJD1mlvDBdPN
DWkDjCOGaAouF8/EXy665427OTnuzrMp2w8AtSozM9iVWlhAcXqJwMTuQfhKdA0F
B08a5emo8I1oQ1gSmg1e8U6/mLpalYOhJkyGI6Bl8IF8wG95FYwrBpBrqxTd8IZz
0IRpxzQiCJzpyPBXEO61D/u8S4zA3lJDzR/jIFIC3Lgu6uIXCOO1a3CjtKUHPCpf
ksTuMQmdwDwBkEn4DBd4Rr1ZgYdzd8vmfhHplzFwWSTPonMzpAsBC1VAdHqN/T9z
FQ/PURWyWqAot3/1Ynb2MWpWBlQ5K8Tugm1aE00N8b5NkmfPadmORXcxa8hhlagF
2/tqNg5pfiAaSJ6K8r2SMdOb+pTBcI4a01dIjcRMWDPWGdztjntszyt747O2epV4
GcaZJXA/oTGcBlu/KeZAQ4NHfrb1D2LOIWCOoZykWJn1BxwKdNrOQIB2JUjNQHnq
kTN8obug4KxK1bBeJrHqbsY3oTwNiX2B/9MM8hFAj4zGuEdljJh+bMCj6+Np4w5Z
4H2z45a1HaymLswRorU6OYE/bUSguVwD1vaPCoRx2aJN3m9DeUic3n+rH83jK5+B
W3d466katE648NSZACf8S2LUYZD4o9ub37VHWd44tp3Q6IQWrLid1h9cTJm3K3s+
02GRR+n0Gt8M8KhodGeSEf9z7ZWmTN1PcDD2mXAn6SH6eYS1/UNV7Muaq+lM9x6/
06FV5G6N0hGLzvadV+Bo6BWG5j3o4NZiJE4/3Pfw8BN3SSv/dsIizTYNfwUU6o3F
UzjtRnG0g+gbkrQV3CaQs+Gjm7jXF+BUSjt9Mrm66Wb+npiz+6nOBwZef5/isQm9
GMEYJpLv9Dv7+3TepbCc3c69/SYDxOOHLnSJJgh+9s2i/7YM4PD9bQGXR/CRm2H3
l7EN9WMgkIQwPECIrYgW2fUlgEqVFnTjbtKMpzWQ2EZXz2CDrbIcLv9zFb/+fUy7
cf5JT9Q1k52GS8lfaS+facTvLNDv/QbTCAAapAAjd+0ON5NXQ4l11v0cKySQeVsH
8pXNRQ0CYTJ+DJz2Ngh2SrB9S10Ftg2cl0+K2cAzTbj4lcA0NvHr8EiW2kguHvMX
9xMXR0HgxXDR8gIxyMnGuSWmNu+TI/O7cZbmwh+/XJhfSTbwQUMN9WPiURu6DZPK
Adv4rS9gWi2ElfhWyx1hxN3RrGd9d1A5uaLsoAttENGGFfh7wG+KQ8KknpyXfRTy
sxvPHIwqBjOIcRTF0/Mk7r3V7KLh+uk+VYpqOZf1/J2LjKGyPdgCd1GTEUbE50J0
99hacdo1sW0MVcfSsbcvqKtGWkF/0prTNK1MYflyu1l5rhq9S/CjYXxDlwG7nopm
65242rzf0XmaKpujHkcCYtsFMvyM3OF7DHdQ5ZaQ71J9nrQh0aAq+0dV1O2sTWkl
QXakPp+I3J98Rx0sNqF+6eDpC7OpOfT9qSpbZtu+/V7hdM/jwwCJ87j0lIggHf6t
FXNbn/TEPFFgyw8VD9itCs2oDX7w9izOYtX2rBUkv0605NyaEipIojh6SHZd4l9N
8W0EfM99/4n0uTKFuO9HgFqoJhDaNAErOAiWswMEyJXIQukZ+Ggd35o8Gk2owZ+x
nQ7AM7BhX6lBWhMSjPUUuJLc3SZg9BPfQqXeFhRZJOuaISWzSkrHYh4sTU+hyJ7g
FsHtq43niarZTpzI1sVF13P4JC0iNuqEKXteXt+QedRQu+yHR2G8yOP28qi2/dzi
bwE8CVhT0i/iaSmtrpU32c1jm6qdzmMyx50ZO/dQemcbtHm9ZVWGvGIPftCf7Gau
IS1g2zWvb17nQj7qCICEy548jaPU4dOygHDQut41QE8p8qNfNac+l7gLoXX2Xh4w
NXF6qGar3LjHUk9YYMd74Mxu5jONoIqhAtUsYNrWEIO+G2vTbjlQkxy+xhxrtMNe
uynjK/u8xK0MVwl9/wAuntCdxRZW8ICFJuErEMRK9seCn6ExAVrdQfeHJjDlnM6A
U1qvPnTb5Er3A9LX7JKvesvTGaob0pyxsURH8qFKAvVqQMEnNiDXzxdo4KHokiBI
oxszXBHnhdu2ZhAbUYVHCE00ANMDPfi1jHyWY3N4EouLa2X96WWujAGlDwmqCHTy
C2QuEBQp0JOf5af/IruBgi0znFF5zaOjgjFz1lR9h1kg37o6PDEfERVPzIoj8A+P
flU5i5IYbA29EmLVW8tDDaCqDrohuG4HxLPFrctVOGA2k4TObuAnhFXPJm9cTbVk
uHe/9c6IY4TThSx2CAWkXFirIDb+z+pR6RPmndjKkVajEdDF16rR8gfvlBBU06qA
7p5pDfoI0ZdeArls4WUN/HYX4MgUcnXw2nNrXP/rYJ91i5l++0r43m6McpbmEzb8
powLNIeEbN3bISvU/j6aqy8w+5o9Wr/kXp8V4iEmbvUbd5TAsoJPE89j32c9JpWq
zJ2qjzt4tLsK4MHUSHTLBdU2kl/+y8gGZTmyC9HQVKYNVjNhcFndTv1de0qyCTUC
suowAFTgNT3BpUjS0YCGdNBNCSEvVmG7VfFjFoDZQ01bV+EBSj8qs+Dda+PV4H/A
D32VSdSTOmGT50UK8dajwVP49GdHFB5cPVBw4HH4b6kMjcsS13W/POGBB9gHxTPo
KJdf44Fb+ZGZqFX6vWz3oZJmGlV0K1hTXJd08y+uKyx+QAT/aE7ulfqMJM2wJSDQ
NLb9qh/mMZd3pt4hkaV6Qcep/5bPWkDZUNbt+o8Md5lVYbBnWP/k25AoTKCict9/
vLbOF5TkWV2aWgdm87SU5P6nVOYeXp+cm8rmIZBtc36IDRnZbrwASXKrZ2cqqZ60
0gkwcz9WGt0knjVgedf73GM5IiO0ZrWFljpk0/LyCL5EixymE8PSDf4bWEM877X6
hdqsWaA/Iy99VSIk1CKb7XBrQyp+P9vBXl5KxHxpmdO0lJhhWGv3hiGeqpwJzVut
V1KHWA2z8d4o5HBgElhsp5Q/RUB241RE4Kp8nDq3BZj3jwE6yvISsA/8fnv79kiB
OwrYva3IE0V9HmkXC/Fc+MDFUUsTuj5G9Rcfw7G/aa5pBYRt3fPdEHPNYD36tLeR
aVDj8FYmAa6R1mJnRpNHsTa7w2W0+UPA0xIkSXxvRXe/pefIViE08URBQNl3gpHM
GKbeNzEdPrulOMzI/cWGeEv6sYJ1ZJ83TVkIFXSTlplyhlJqzT4wG+LpCc7tlwVg
+Q+YEzmhmPZ92CVry2i2QzNziJVRAkEFu1L8Hnuqw7TwBj12VQby0ahQgUr0F4uO
bpBJZB6krc5WPPvJJMT2HRHqKwQQLXs8Lc9e8rRKJZlHg1V01yug7zH5HTzXbcvV
ro6W12vqljCdqpDroJ75GE0PnsMiO0cyobcAkxphlPr2AbgbR5s5hf5pxDpidEi+
6P/96q6kBOKECbIiP5nbBRuzmia448HMNPDeVvrIfnpFBiDUKuM4/firG8gVJzc6
l9SDgJfDnqXjvzt5iy521fn0yS6kqcyd6j91vsW9YROsx7jA6UVdh0Z7WL12nEKG
O9TRetdiMkYr0Eb7eCAVtGORggSzfsQ0o6Kx6A0izU4AGHt7GUgQxaY0y/IxHPK4
S/EJUO6DGHlBx5BPGEtMp0pgcyAst29rELDtnaIgHkzvmSBSd/ykQ9lnbcxWlFOC
uzOWN4WVvCjkfKMY9m93oONqZT5WBLoh8mSAX6+pG14Bo8PcgZ0aKyCgcOD8/Mam
QpKVncmDWd6fmRkQb7SNKCSX6L4rsneac6tEeyLQgPl/K1xL8w23auXf4fvL3jGl
1kR2yB/Hk+rffC98vbOQIFi2j8hBNDPSV8F1k+foMQDzTERAV0BFVRQ7YWuzpxzV
B8dWml39M02jje+6g9+GP6+m8JmDx3gh4s4I3ZwuHsQWRkiU8COCy/It2Gouzk/V
HXMZkgamJjC7MvMZM7RJrM5F9jMHsQ8NvY7Ny2VAF2sDQWDZIm/MwGe7/KLw4SjR
gm9UTPwI8+xFtroh5juR/U1EiUBoSQPQbScYW2p9+05mZFLKHmQnUTfslRMN4L9e
NAcovvU0LSFVLAUSJFoD+Oo9teXSkJdZ78EQqacmUrd667+xZztY+k/VCldhZYdB
Xwg47rd3b0KMSQ4SUF6Gy8H3VUzCy+50dNcXRPLHrliQFQnhqHFr6eGBKQcRpdUf
Pbdbjx74ionhItCGZ3+yBeAorrBjJJul74x8LJNZfprW4ZSHzPI+MnVJWq7qB5Qw
EvrCG5PJmZz9fKS76kmkr+obGNFV0Y9yXiUZ3fr+qYm3MCif8KV8yws9zSJUd0+x
InGY/Kplny8OPDaLGkAIRpEJlwxre15CTvoeTEEHn7JcB9aqw+3FJkq/prSXisSp
w2TKoiYvI9d0Nbijrrwcgs8m1hj+N2JGQMSYyNoMO3OFvFP+DBx2BdhzrpBXl+7x
jSjtnbRQygQHA8viG1Tcepe03yqeuydZ268TcdXdQIt5PqhrhOLOPFKm+oqVC12q
+ZbFfMU2nPIG8UWkZN074ELdulOzGIDg+AAXtX8hWAQMXYijoQ34od899hWRYcg8
TkPqOXpSqcHSSDxGTGSc9eiuCmN5BLpzjx3BaWVr1wLVvhk+PCt4la2otFeJbV6g
Pi0bXZwxWNCK6X6+Jo+RlMQNQCmrlET/K15K7S9PMWU811boSuVPKzt7nNttB769
oYXBxPkl8R+DsHBiWjpGCQou+t2Drg3PJ7GFNtMU4xvkqJbPPAPy/7EruQZTN7RU
TTfdqSZdgvxywy7lwLbtt635ByCGUhJb8khi6FSvAyKhEZROGNWhmU2hKHqDYNKD
2AZ9sSk9aw3h2hBmt1RhJseV0V0NgdSbhJYy8YUyvRULPJ/Lu9g778bZ4YRb/s2K
1muS26kdRs+hl+2PLcWWQwJynaoFag8qgi+Te+BAUl+ugDFEXIQoXtTj2y2mZnCR
65aFnsDtxZwsiFr9D5AbI//rbs+Osq3piTEKB2PzAB/kvHs/Yreu0tiqmR3JqlKa
onJs0mmJu2Iknp+Ys6GrGH7nbM5PH+301RyA75ntiNs5eaBD4IXTtTy2JGIqmnfk
mK8rc4Z2elC5+eF3C790cqMqd8zgdkH+SpW3U55MPapWZcG24zXIZgfH6I1TnqP2
sVZ5cnAaHssBN01goUCdwc3SxqUVzps7e7yAEq2S4poBaWl5cZhCjyCp8m9ZmzbE
YYZdvC9b9jvP44NTxNFFtNwit9DZ5NU5D8zUm8OX4n+Gwhdq/xx1VtgC6MII0ief
fI8bugunxfzDvfuhCRVlHdSA62MBkMLfcFOOied/qiqfUHqPj01YzUcJnx6L6Wgw
pPbbvXEVW9hrXMonYhvJeX3bj8rLJhMmu51Q24wY3Q2UA991C2uDwJudROc28Vtt
VuUHQHcVYKgpyVmSrVi75/hA3INZjN1pKCJj7l9Ms8qBJadetjfFASKjtU9T6wU9
Ou2mhsJW3FSo+MlTcg76TseFXhoSIpiIiwKPXXjIzjrRi+XP1SouuUiov7MNp1X5
4sxqnSAX2po37ir39FO9CljcxdAeod8p3w3bhi8ykFQo5lKoghXDUsEcwsZuTjwI
Qm/01PBoNsSYBMBVl+Ar4vN2b2rPnP3Kxf31YC8lpMhF+/8mt+6HeI5QSSlg21lE
DrjA4DcfxEyc+S2eyF9bRUfZ7dm/f4icFpAEihkcz4USnMJgWpmpYj8BxTvTw/hu
1czu7p2gve+YtxklQS1dDH0msp3iLwTG7KrvtQU64kJlhXSEOGzb5XWPMvKoiwv5
gJvHjXT1AcY/S9xkmnfX96vcWtJHt0jBjXpd+o2YAxuJOY+FVP3DM49jCAuijiBS
yNYS4HdnIsyJQAidAfj13FUErQH4F33MVonGxpgDjNpOy0WKoi33+5ccxYz+el6i
vQz/9CV9KV1clw/ApO4XhYclG2icenPYrgj3z1zEdOee2juGln//wAd8qEEQ/EqG
CDn6RHLiPFegJSVln1kiqYTErRVZE8pwQcblcKgsCE45xFVOmkifnOCPSk5mEaer
Pbu3QwL8LdHaT49JE2SzGnJT9S7Qlvw2CaEj9lhWq2+TmqHfSMsnnVoxhkpkZLOw
ebTnGX87TtWyVg02X3CaO7yCaegNuFF5VhQk/rQ2FGLoK/rlRQTLTlvH0e4ZAzHF
74jJo409dCQJHYPbXZQCaTLk0rd2Nl/Ci+tB6l7r3/zW54SEW1wr1wZnEQ0kY1IC
VALsb7Ib39KqjK41BD1xq6SmXRIB5L4pQyGQiRVc0JrlA4dn7U9y4oqi/nvnMfkI
K2BvFs2HD5CtYONhZUPmmGRpZlPuFkfwoiD7Rp+HUlY6p3ld3AbomaXsw2xGg5JH
Wo8JelKlQ94tLPDWN5GNWyvMmWRNoCEeBhS4DaUgPwiQZabYGK8wjWNC7syr3L7u
LlYnH+1tZK5EqZxzofOKzeW6oleDGy+RqPVotodz7SzRVC2AHw6fOyzBX3IZoJQD
jxPtjKLjFcVb2PYbQsskuV6QdP9LQn76yrdEfDKC5Bjm+gFuax4DutjAnH38iY/f
I/iewgMZH3IOcUSxTOH0eM6perBbqLmT8khK09SUvSUl59A3xWwUcsRPuAjj5D2Y
CxUEsnK26LM8bHOLBdLGMDOLbVa3nV3q96C4EKvESM7ne5uLptpVHG3RWhOjQEyy
d8gj/1UUPcgTLr8H1pMeOhs+pKdTNVMs3gCJFYh5guIvrY8y+n5uWd56Y1bNwJHd
M6VDuXTUWQtYoJGwA0D2NB4eKo3yq7A7oXZ6wt9te2hYd0PNiGiwO9/NVDdeMAzw
NDGxAV5vDeccH30CnImkwtoHpWT+FyedV+DiZiIWgO+8SGPU58iqjED+aSkFbdZN
cDfllffUfpkGzBmQs+GSeYLr0TSxKwbbe81IbK4yUw75jUbKxgVFZyVY1ykq1us1
mbvuI6drGQS5Z+9SXhjdFqK2xG7UAVywXLn5OK1ci0BLfcQ4Ty5+MshTx+Ljdvym
YTscoK+zoETIwSBu/Hsrv4tOKrNdO5kM24Qhr6KzIvus/mqIGXvP/wTBXdjF5WVx
UjcPVPoFefNqmi6go+RBIEet9z1QANhOvOx4S089s5jPW9jNnly6Y4FefIopGy+2
OiVvYLdKCEm7WC93eSZkuvJaxpnV040hM5HqsBCkVcKwMEF6+e3ZGstiFKtD7Oms
vtzUFHK/L7nMq35uyFsiZzYF7UKpIYApfhmRuUd4EejVeIkFMekKiChIZOw9IvbC
V4jf9bMjoS+DKJso8DNr7s7s846F6N9tMgrhVwa4huAtmkd6m1PYsgOkkL5vizK4
NKRSrnUTmHRpAIqDVlEDm/VKgU4AV1CyZ4BYtYEGdqf0UGfVZHN/ZuD+l1P/hD25
20eK5Z1bmw8RIDfICP36h6Zwr0UnFbUo3eEBdywnJU7TngrPc4Q2G/8a0u8Lt+Fq
LO1UryZDxMEldD0eiSUnLwgq+HTmTa45djdPJMh1HXvfjnLwARRtsEBtgOGdlGEo
TSFydKi3UKavdgwbbrQNV4MZew0CegsGnADuHQfUIF/e/Lpfe6A+PVtC5RSX/cku
RBpJrh7TP2Ua96YpHG1IFXlQJorX+0E2CA/mf+04Ue4Ug65QLglAtBiEfDu9BeKE
kUJV9OgJf9y5o8W04Tp115g1Rhg52fdpe9K/gUMmk/HPu1MOBvJ11rxas+pucp8f
2kLfGT8itQnRnKxRyk7IqF4wWVLV/x0lp4oYhWgMXxuO5ivgyLVr/vHMsx3jJiGW
80qOWavpxHvfx0gRVBJ4RBP7it6JWtOHPMBT30ny/eX6sLsB61GDMG9RdxpoaMUf
UpUMlx7g0DVEANZTglh1YUAT1vTneHt8TqbygkMU8fy0NEoZPzYpnneGFWoNyc/a
WGq9Ax83tnQC+BtRBhtqkdaRqeXZSpc0BIEkNrw9qkXlWDPqfvmK/VWEysczlDdk
lof/HZpzqTTFgR+q+3rllMxE8z/3xqGFf/zPzubilzXk1yTe9GRy4KCgfAVzWPQQ
dudD3odTYh9nOax0tKn9TVaAFjDGKq74KblwHoGU+8vwVi7oLFvlO+xDjlWw1B1h
SOfqfbiALsIZBYjMUyuloA5FbrE5Xd5Ygu21ajQIPn1JiR9WR5zjcwhYzzA/84eO
8o39NpJ2qyxLEWGhz+nTyoM0seg6446uO0YjSUB+6v58oXGrtITDhAKM2+aYT7xi
9+cWfuTow0xAjdbpKjGO+E0DzMC5pkiUJHfRhtP/Ny1tQcRtulMXwAlNQZQzaNaU
GTHr50UsiliVAXuw21YuOrz8r7p14yJrNGb9XJ+WJL9G7Dc7arGGMUT08CjvwGRx
WK5qEMI6wzCMviFZZ2RdJEYiVVXFSXfLLV7sO9juKb1ZPE4vEFsjHiwd/a5J8Gjh
n7LAEdj4Z9TVOZh0qEJ0vl0jOzwDq4RMG8cpYhotGwqh1cS02yrFc5c/9jwA/4Qi
xr98nDK6WlYP8PJ+PZ3+0ZZPkbnnxoWMLugWZlyw3kuH4yy//KxmopVgRIkh2azU
lSqDard2uAqyYkB5QVhH4kftac6sUcdHF6gaTuMSw20zdkoDtiwsL4WyL5YdrwmP
AyGN42pLz+W2kPE8yuxPBmiDO0mxg04XQoA/IMH0zJ0vHJLkl6wV9OasJPcYy8YG
JX8rhZMcwxd9kF/odVoskxr8j0MBBA0r2vMsdj4MjFP2VQ+hzbigj/NXw69weCYw
0phm5J8heOu4g1gC5Odt0kSjXIcM3+RUUPKz0ZJVijUwtH4+zFtpy1w/n+diZyQ7
/M6uvm/lTj2XadMzBuyRA86bngtmRKr7dQFehUrtptM8V0+t4VoMlcAO2CYhCLAv
h4R8w33g3b/G1tKdKCFdt9Vski/rBMyMvza8MoGO00XncAgUMFBtjNuAtQhSBDpM
2G6B/mo6YtTRD5ZTSv2ZOy691qII1Dao+ud0m4ueIDddKbNDqOc2u7cmes8qUg5+
uEtw9Q7/ReT0HNAYkxutGf2V8JOhcSbbB/eildipee4Z8cb7vglI93+tYHwK8+eI
GGU0L2tW0hoQHZ3+UxuUsBGthssn0mBMOJp3BgAK0iIzBQakJW627RmWl8VyznKn
UjbCPWN+pGzKyuwcDAhkGqUDxcxtcJvLtH8ScjILRnaHHLtQFQO47Z4Dkr9WmgEK
FkDFgSQYLtXXuwJS8Ets0ZCcjZG/jpzDMsEarb+N4wEai82uwCCyfgGcryd1gGzU
19iBTYp0fbHVvSOES6um7AdEbtwy9JfE7O2Fh5yRjPZ5cnh1PmdHpE+CA6TU92wY
HYQuVOgJu1sOTpui1Qz60S9p3WvgK0YPR2Ps4L8cgFR3WnVkEk4Wrk5l4yRkWUfn
e95sRBCujqnZKDTOxdCXmVsfYITZnPZ1DJc22TOwJsiZ/Yz8sprUxop3+Sx3LV6c
V5tNrP13M3AVCdCbAQQ2ZqjMbIzF52zs1v9cyfN8c7+Xj3lF3iOPKbd6B7J4orqI
h5SeJw4qeT8sHl7ZHaO6Rq593jm3pF+jg/C7xpZ7BxnMTBQzNsxL6nmxDs9SV2ta
QED8Q6owuWbKr+izQRHJ7qCNdxWr+Qd+blV9HHc17WfpmJNqcLs4abqvSVNyX7mJ
ttTwCAjPO4eMr+0SznZP307ZFnL85LN4S+R6iME612GCr9TnP0p/DX+KSW9vJGO4
k4Ek4cJX5+8i52vFZcJaHP1oucaLasqHjSno5epxHPHWHr7X4dQ8o7lxuJOzCLfZ
5DgfFQkGy112lxpfJhD03p6Q+asu2JJ6pwpKDibdm+3gsLd1XZrhNlM9oT6OGkvF
ns0uTgTbMkYGc0oAtIrJQ3crs7c6xxX5xTY2H655Lmr+tDLrRntCsLjGZvD+UO0W
ntDF6G3CLho7+0uq1BKdnbn6P89R5JI0i2b5xRlDLA2kGogxY/NFRWM8Dh1jawTt
TLXzMKRkoZ2F7XVfv2Qpox7Z7oK8ozQyPhfVciRwxYvB7xje0Gnr2zLWAjUyYcts
Q7pkGxrEF2Dflm4kJiprE/Vr7qUp80JnMF6bFaiguT3tYr821YYhRlRez4FbvOyX
azuTnGiiHmR/nt+iBwpg4cxHaJFgATGxbgVX2MK1yIvyC5dJIXKUzXNls5i2wgKN
IrVMZo/QjAUYezzOcDbb3uQOx4hDyCf0NWpjIXZV7RRaIux+W0xSmeLxVKgAldPd
jtLA50saM6Xatl6Wg5AwjzR1+CwqUGaGSaoAJ80oF4ZqTXLpNV1kzY/aUKhCA2Wa
T0P9FdalYW68XXCYC1xzHIbrekrW2XzvCH4VmxwWCv32utbdbxnA0bnTQG60tAH7
ypJWAb8BU0cBCcZziwnrFWuM4I2RHkvWxgDyxFWICRlKAvK079W74dEWJKD69Rdv
P2i4Q+pRoPp7aeyCi164CNQNl/IOSXKn22Kd9ttLSZ9gooPmdNS0HAMdZwCddjtI
U9RJgtEA2kExldiQiyhvPMFaCh64cZ4+iYjl5zzCPiF4lcVKVDk1YDF+1KDYA9Nj
MTyrt+PzLQhQJ0EhOb9xgdy6KTeC5YqncWHZm5LMav+RebWodbOGFeaHH1b/fcmT
Fp0rBDPezOZ9O+zyxecoSL8aq3tHIcSQI+9TlUOdR7lwLInQgHvX97FPnT9zhzSy
s0eYZ4Iliph+F4KjHIcAk37kGIj8BAE7Etyohcj1tS1/+31htNakJyotYpQ3dXDH
qADiTnXohUuAMmjHqQDVs7J9h0DfrJTWJ1urkYe4QMPmMDuFwrzO6IiHfNcnaLOL
ZwfIeA7RgjSxBOp/ia8m81G/T0VEYx/rvdqezmoQKzw+AgRrt67Aprv+hTO+zuFq
zvO7pxUE0Np4xLZEVULJU6r9ZAPIye7nLE4L86IcY6uz5C8ltL7pvVKQpqLzWUXD
J2bpSW4Y1mXmN8cscF2RWGHw++HXg65MOmQWxPfZn37Qkz+bWDfyzZr1N22kWDRL
K60eLAxVdxfMsusm47KdXDQl0r+IME+nAKeQBv5JBCecobNUEYPEUqdT7QafaTHU
uuS1BmNViyNMlqIQJnNDQnTb596Bjramd5DyUJFEoREXGrIOxsS/wqKBd+136PW/
ZBXYigHbWf3u+bjb9aPIreJU/au93B9U0rEaU6Hf/pHuM5IBFbd7g3iJS4/IpFNF
7auaTZW98XbVMihuGjFmlylZ7X19aVc8+/ZsTMKnvv9uQSOqgvL7RwcIqs6RO5mu
vtE3maaluxOq2zZxZJdzkIdf7DPRCZ+J1WSQ1INMgQUXYFoygoOvHEO5ljTbfr9E
vKAUlvQBsKNZllxrZKvYZe9AOsEudRjfCPiNjHF0p1mla5oJsKB3+n+g+4C7sXLw
mQ6DW8k0kUH3UStIJu4MiZSBoUX6gD9Ju6ui03s74vC0/89OpM9awuWXcR6tJisV
GPiZ1YV0WJ2K0562Jog/pO+WGJfNWgSeNDyfN05YIKFrIDf3KQHxEjbK0vWcekCd
mFRdseT7kPVLBiPX24ZCB59v95E1XxN+315uPqSFEkyKok1EEZYv8+iAgm6flN7w
cBPzxfxkTPymt2Bhccd96Ih9M+nPU3VWeWtDjCPZjFKX/uR8lbB8W2TOnEMdaLw3
cBEJG/qDsnIIgJUTokvQQS30bkHB7onu29ljx9itfbpxwsyaztSB63k+HJhqlLT0
pm14R0MwtOM93k5Do5iAfHH5GJOqDbBxlJNeu9DNxbuRCA/2P78kOwdV7mdNk7wP
DVcd5g3JLz/CQ2jQcWLs/xPiY/1qitS1L+h9t3/b6oJdzA23LCad4bvb5c2WXHjE
XCC5XM5wsQT6oOXuFJTxPIKCRlx7Hjp2gsp0bX692NWkiRzewfEbWymzLMU1Z4EV
sq/1/b9pfm+zWBQvX6EjaQrDUwN7H7PT1Yvkqg8mxkffMHoTGXPDYW1vew+mlla8
C7UboIXYwOMj2ITPZ5tfl7qRPLS5jtyB+n+ir4LkLBfaV6f/cngcl4UuXwcitDaY
BXJDwLTKKx8Tn3AylQeUm507HUI0AcSqQagAcyEN1neRdAyh3NNrMm6bPVgX6Sta
zwe+F2hlogqFZ5bTDDs0UHlOvg3i9SEUh4XhUExcXQlm+vXiXaSRV8ougMgG2FqA
cx/rCjsX4r1+FXSryQhJlmgyMZGZDKZNXFALGsZNAkF85pKYsLkJuqrLzIiabH6t
5xanesJuN7t24a9OXm+XXoKIeoCJJb4du6tlZjXK6dP6wSXYq3eTQ3t3TfFk2fcy
GuG4R9jJUyfHVVW5pjTJCwXReZ1DpIukjwCQxVXfawA/7oiD0NEU4ez29SYRGWg1
9b1/AaqJ6mJtG6XqMUK2zf6hpF2UZiWbN+zM2BTmjFrHg+2Bq2bfZZBYV+fo+JqY
6GBqx2doGripjuxaNbF5bwbY2ijGvhkS5cYgH+oGTGAZawcIBDiK45APiXkPx3po
DLA7tVp0XMoquGcsnkaEJ9FVCbz23ER8985dLaHxrr7+v+CP7stPPOi7yc6KlV0u
4fkoayT8MOjiydWHltVlIU5nWLxztrwMnhdVZR2qrbu6Jb9UL81j+UVfF5B2tROM
ATn0ssyUx+UQmiPJWmep7czZZ7dTWvLHiCK9VRiomjkXgcYxqzYgsEFMozErZseJ
XC/1URuw8qsXQoGdxRts1uGYp7LbZOpSE4+Y1XvR5dOZUciavGYl5lkBROXKs5B1
PRMOl3BP9ZpUwGlsh0cLWA+zf8K753NP0Rx5WGafmYJZPsqAzLawZVNXrH9xLZsu
essqYujHq9FT6GByXVigJIrja41UPIgKgDXIGumjFw68MMeVXeLjfG5mJvqeSQri
7IFq6kAC9+8RmvFdgkGa5yX76zd36xuPtb9eA+SVPvdGl321acw0rH4yWnC0sBQG
9xjocaYr2GRXmMIKf0rZUK9PdM+UBUAy9L42OoGuXy3jNBTf18x7TRHH8dVoyjZz
6C5fwDQ25adZellz52u2mjWk4CwIbvr3WlmQ8ekswyCO8qGTPli6HamyahYoce56
95Af4xuVa6WrBgzWf/3a1IY+XmURqlF9byMSBVv75zH2AM5KNoym3ay/lqbFSrIh
9bsSLMtiUmBzvQd5qoOr17x4kKmJVGNsZwHB/QdTKutc2o4ehi4EMwUUDqc2n8Au
BUmymKoD2YhH5YbVR2oRNtiDNo07L1M9gM+Jo2yyPOtke0qU6Yty4BHFJS/aYGfp
3pfgHcEg5qTRITHyauZYXdGU3oUlGphjfZVDz7t9qu/FzvP/ssMmPXPjl5OsSpYL
KXj6BzNpe0KOp8TQ4uU5ajVULBGlkEi5WHg0XhxEU9jUClDHK0finoS9uQgvUZGm
L1jymtNaUAkQURE3Iix/t9UgwYLCVIKihLD5OdbfeS1C+HJxpBJihQI+w5EiXaVg
ROUYqFzDhvzB+QfBfxzsbupwdu/GHx8NAOk6NTSHvIXJlM0E7ZrQKqm7jdl0yNDh
FPKaaz6435ebgycs8Kg92CJ6kNQ2P4itvWQ+BzheIT4Dt9p8BJqV99zLTrrKLg0I
SeTYcZhEp4pqpHQu3OWXHvudmzqb+QxPKbT5UY7g6FMCKRaNwkKmSK69bHXvfAx2
pYll6heBRXNLEBzG7Vm81Ipj4sIjEbPSAbzpevU5JdiP68CioQXLl6pFmBVpeuS/
jtjAP2cF80c7Se/rUbavFRE4o/+6O5gyZbqq3w2UCAG3EoOigsBJLA003I2zzzHG
Slx2ftvrGGrpaxdKS2cd3A4loT7wnLbAWG0MqSb0C9caLeA/2hecGLQpY+LObZIN
tOCBfC8PBSG0AaXBbtObuiQv87/Ex3xLo6yihJbnFhpcHJ6AaclTlqvT8nJ1R39V
YHu478YoTFhcxahSdqicrVRoXGNtKyufabIuSjyyPiN/k852mD0jnUXPPOXDduey
1b+iXKRfkfrVeIBs5zN6L4aJ61xLoDYfxHuZnjvfgmKV535IQJXPKyMIKbJ1P0Lv
4fbbxC9DF8quFwM9dLdjXcmw61CXPC9/wKoq7f5yyElRdJCdC7I6ZUSATrPFd9HZ
E/ghE6veKSf2s5fUG2/8cX+VfGAoEtVGl3RQ0lOcZ9nn7kHpG93xZYoiG62dPTaa
0lc1S1MiYXdsshWt4axciiQezkI5yks0JffMWWNkv49hz3Dfbx+kZfYDtlZWusgg
+J5iawOWHxkYq3XYUx5bdBG+PuLLePrIoRsSRN6HWgl9qIx1iNmiQ6e5yjwTu8WR
y7+smc7ErYGT66/MxD+/qnLTE8AUqqMfr8sVESBURMUaZb24r5iKUdSbq9Bw8C+/
pR4yKb4q3mKoeaBgK3yayIWjVoAhUdQPeOY8YFiP74ehbZWYGe8uIVyn85B+c0sT
lSYroLF2aOC4TCQ11sJwh6ggOb9fdAXlWkUPWsK0tUxK7Pz2jQKa8nvpDDRdmGUO
nu8EF7CK0vrN091wYJeez10IQXukMfrt8hhX65tMuWemYfi8ZqhgXvhjJ9eb9JhR
Z4pvjLNQaKtvxCOudW2D45BKNtMx9qLJZDb8F1uNOTcSMVLb4SCuelN+yK94dj1h
h5ts54Y65QIU17p2ZnNnklBtt9Vv4DIVvKNLIkVwz9vc5yMIRmlNKk+hDGW6xXgk
eHulbGy1SE6g0/OqRADkxmc8lbm9APbs/xCXNJ/wtKfOGtwDmcrX/TbF5xxmOEy4
mbsZB+Nf20zTMC9J0ikVAlfXoKd3RaXSyX0i6+LAaxVYXi1AcBG0egMU2XOTeMFD
Xlw4WRbcwLv18ZTRw7VHYyTKVWMxiD6ZpFHGobdTfCMxIVhgWBrYWJQAdPeFPtU/
0E12gc+57iKNjbxuRRlH7snSncNkly89Etx7xaQBc0lWFa8lxklfrySxZl76Ztao
QKFy7187OHSE1ZQpUHitOKOIAqOD0BGL8M4WhnPXkNxgHzlarerQ67imvNc3kvUx
LxFzThweQQ+lbLooOWtcwzdU3HdA45EKshBhArdTmFLb08q3XrCdU2EKMgbZBVoI
H6xIeQ4oDst9CTOWXCbtLVPDGaO5XH1D8qfe+rumQ9Ck7VGGrorpYOeXmbwmlhai
wgMkKbx1VgQHGK7gK/aJ76GYJo5CcTHftWRfssjbL97shzRqgsefM/3+5vyyPFUN
sTMmz0SfF3/VDq7V7ueayRFG1KXNJ9gUKG5Do2Bp3Oc/nyI+jJFjdRGMahuaLxQx
5xCkiwyGFR20uK1M/smZsO0Ho5WDGfiHCaLWseRk1J+NyH1IIiUrUulQEyzO6ztX
YQe+4cOkjcgyNoIEsXG/gohjL2trngcdjPnwq0b+YORMSA3hfDJXIWIVhmJOjRzs
mXBtQKQUtlG/ICdIJNxIcQ++yfTr4tt+znwJ4qBLOvKfw8Zw5Bb5H4LlRs3CRazl
v2NpZjJNSyM4VxOYJofwSMnLScIPyySyptS393VkaLcjkwMRSHegqpnuUTr4qqgH
dtTYxfGbalQB8VHxz6th32rd3u/2Bkg0GY8kZriJm8TkeEUsnlhD1zBqY2LI1l6g
0tBx0dJhIasY8EUx8maIB4kyb+m+y9NT0RsCrvKHO7tW3vs80Y9gOE/l/WdJy/Tj
5mDe2fdx+ErYVOAylEnh6VidNA15dVE8eFGTmSBCjRm8Kuz+KBxqqJ470FBSLywK
pY0asRiwX/6PKmVSvVXQAs9L9SX+kS+BLR1fhVdZmpTkpgQlHYjxL0v9LWJpT0fO
1ffolAOEpKG5/6WMEWm1S00UfszQDaLW1WkjXl0ZXuyhF0sxg/Z7B9UUrp7lXGIO
eAbVm+c4iWJFOTbKiRGdTJx3j7tye1QCP6MZHA1PuKFWM4q575+EciC2skkyrd9f
L8OyZpsq6cUuPgqvgH0wutUvIs4r3s08N1jCWC2bX64qPpfTtffhOlNhocV7NllE
ivX12HuWVdpaZyEiPtFjUshLDdxBD+uLjxJiWtxfUFIB19wTKPWxXubE+CqJYRER
3x3tcRkx6BbLqTokA9eY+Gb63WoUfJ/5ge9VcrJhtMvS1eOU5BFrb6eCSzJ2qkdW
llD1X8z/0oDK1R2WzQj/K19pum1GM1gKfJHJ8sTHGg9WI6vyFFFo+3Sb9f++WCBf
ejHrYGMpZ5AkJJMIeH5TWng95tG9bWDDc0uMTXr1I3z2NLAAsHoqxmwLUOfT8W0X
Iz/8q8/wTGlD43OoEhq90i3DOo2feaTSFGUMSUM5SV+AqlFqARmf4Y9aLxMan2Ie
7phTiG8phXfTEsHh46o0wcNfABiQqALmBk3XIfdfdEI3+yYr3SmNQ+LpbY9U6mT7
8SAke28h56jpew1IXPPEd6LY0hgAln0msmXf5kKtBteUNtn+/vnXwdlj0/f4syPg
vIv4uGFjuedmcjgqT4rZqnMcHQLTPKhoEzXO4llZ4JtizjEpRNDEpOTXpsWPKffU
UeT009b0tXxmJGKMMe3RUpnNmItaIl3ZsABaVKC9m6mo0SGob1JFX95uRC97Cib8
5eF26kTuPlKZ3hjSfoCVLboidmd7rqo5t8sX2kpqRTpq8Wi88j/oIQlVKkgwbz/O
3QQkM/5jNx/aVcD8/n9gB1xw/hV7yHd6ocQms7AuqMl0C+P+GouJFQxT3D1Def5D
Q0O36B6G/6iMWj8vqXKAo3Aw99YryLp9c7h39piJYvgNmmN91wbEGRjZd3Db4yfb
MvFRnUIgGkrEh2zgesbUSCR6wD9eEsq/05X7uLgyz8Nmt1TNG+ZOsWL+F9oQ/cjW
2QMgNN9/YQW+z1ibQ1Rrcc8QblnbBv5Yl5WlW33h/o3CuFdvfq5QC9BZy6O2/po4
s59kO9vJPG214JJ927pqdRPbOcJFRAmuQKjkTPBj1aqhb7i9e6Djvx9TqdrqOZ4x
7Zpd+zCle4/uFE6y5QRLAXoYJ5hDhFUL3lF4/aaNbWSCxxlYdxa/hACmDB1EkBAg
b8b5yv+JyBLRfzKStbMa/YO/IvMtEbw/prvBNgCX4kbD2MQTPYWMQFMustzG15it
8iQFOFdzNTV0rMoz0CPIYezKVfUpgEXH6eile0/XSeG6kzpIBsZ6cvsEGGDnBOCi
R63QbHJWzzY2BSYZyemlbf/AzVLv1ijLzi4hsKaMFZ7XBiRRhOLY9dM+96MWJN2m
0HZtMsndYhQQcGFOgxUu+0OM8fTgiRLjQzegrLZ62dKwe9p6RuFnPIgBsP674Dmc
PCS8oshEIAKt8N6ZR5yJXZru96Q2AgYybGcBl84KKcVMJXDMs0qcGUuGhqR4DddA
yjmRrYNxGqEo//ZGTXPV3msRmWMY33yQsubIaCw7fIryBCty0VNSoPPfG4cKkI/U
meYgHvUwQjOEUqINWakqKoqMpOfU1KAaIEn8dPojB0UjIibxfDL2Iab9DBfPSzOj
gaZFIAwyrdGK4USlguRfxe25Y3EhsP+bhXLF3hiQq28+9Kl1triNZx0UN1lmbeIe
n4dr5OLE06XmfbWgSv7uG+d1m1OFRvGS1Bj/yiOsqtxDhSCXf4eUkRcmVzv+q+iE
C5Axcfyb9KmFwuXD94bN/Oj217kekjJHJXkuEOSeEpZKVz9cFm7xqnjJIitXK6I/
JHm1F71MaexFt0EaH9pMD0fr2m2sM2jTpaNi0gsWF4kwYuBLM6iLHiEr2gZyXZ3B
bxs5dzFYqUyH1Kn3YkxH0ZqIg2Xza+UD9GANbe2BZ3ICm1U+mAdSZ/v5f4qM/Fa3
5m0kqqVqZbaXg8w3TqB2Dx7D+1XkP1mdAyzH2d15W+svBREKOAU7skdIEZC4wUyD
1NpWHdoHYZDm7t6rIrEyK+LR+4hg9Ys9zdHYf4B9axPpXMPkGFRavdyJKw9aCHbD
s8zEZP4/2GQUfFLxnRnjQ5YKAIYDTPgOVv19etc1XMpKbtf0B1c8nO3QVsfkXnBW
OKeqgIiOfiu4UZ+tvrglvzrb+H+vA1fc3DhZX4inwaIf3eemySi7M40gqezTCPUS
ucamwIrtM1vne7WXhoYaw/FV7aaItDImVSNh2Wj3g6H+jg6u3SmhyvIxSJOHNYtb
vqew5GKibeuNFLKBfPRrmK9mqbAl75FVfcWDANIKSguG+z/ut9wjFf+w3sHHb8vo
JS2vXsdHq6jxJRbY9fxDiy5c6gg6O9wa41KT+HKBK5kwyNYH4Uza44i6Jujib/Ku
WA7Zc4GEDiKTX526IUgvHmIGnkDHgloUB4k7ZoccRWutG9cDyAx6GGzHfUdEEonO
pa3z54+9T9ormFotB167x6VFQQx+Ri4Q13dRWPLzYJsrmgBRzuZ/lOrTlgJ5Ktyg
mwEvF0fndMnIFT+373pUafFI2HYybCRLRKpp1TziJ1xjLnerVfwRKobV3mjGjmcI
Uf+OK9nATx67THQU6wB1XPSC18CXbzPXVuFJ/r9NOOFtSv3el3nKnCpPgL9L9ua+
1H3/HGLifIuK37fDinbgJs3M9nl7xoaXde18P0GDwF74OsRO0ZufSh+GA9G8eU7L
7NpBKi2F41HnHToLhDO9dmUi3zfxqp0Xic5lfbqpUI8UNNmgAX0UBQwudV9srH9e
3wcH/CQIWIXxVFRYicyPbX+uXO+jfSGN5in74KK+KbxuUU5sf+0eF938Sw3Ifz3P
WJfkdWGGsWdqjoKlN5+Q55pLbEqv7bC1xAZ6NZUTbO7noN31+m447Uzzq5nzmbcc
adSLMbCABF7/SJZ8vLmRpB1Nawa7bQ11EKUiHN3Mq/Bj/1ofpJnXXgYiA2QkBfUw
lBDTX54Z7zQzSnYzxhc7leoHeArfDSENislIp38zaDLiguj+/xRTA9ctUUWbvfT9
jPEjplMN2sYfCMj13TpZLB/ZeTFU3kU5yHjBJ7NsJnQ9H5WU972xBp4xh8mN4s8V
e2ZbM4b/owqbKmBV5Yl+x3imEpNaO4uxr9yvnK7Uxa9foHYuylKlaK1/5ftNf6fG
kqPVykX9JlLjVfpcICGH0XYO93VlTREJWj+lfc4gldJPfPGupc25m0kJ+sA98NLj
SDgpi4LxBf/yyaqhHcK/gAuyug9LQUIAQ7C9aVZ5feUyx7Fqbxelk16/MslrsZAB
yY+InvKZD8hX3BwY3id1YWX+RVbvb8fBguCMPChcxFOxEPPCKONJtCK7lUpLxmIT
ZtLXAT9SunJc1kYz/pnDtNzf807AH5aZQAPGk7HWucT9+I6Ft5lKLAr9KqgM1uzZ
9QX2UdmbPJR0gu1acw5h7lde/Rgc/kOyluS8QT+fv/k0qcXNCJ7ubpG/4rfj/gEg
dre1+LU/JgIHz0GtZ+OieFi0U7WcMzUSO7o2ELT/9mgnDZC3yT1l6b6q/cwoxyUJ
PM5EbQH+HZs2Hx56FoUH6At4uiokzOoKDa+vzBRuZSpBoxQdvkJXFzGri5eySrDt
AOQfd8ksfk92TFSFitf8+1OVg5cCnjrIhMQYqZNofJSafG1tiZGIh7c+4WANyp1e
Bag2VvT/nUVOHDw8aRl+aKicUkVLfn9rbQE8a3ueS966+3IiCInj5HVL0tOMxxLA
xZ5+MTJ6kjJU453zPgF2FtEZueLi73Ndp1EsYzUaFGBvJULbqR/suzf/hLEYwblV
egA/nriiDZj95DHuVBmQH4CZOxn60gakn4LFBm1ny9hBKaYDBCtjze5YmOuph9eY
NYILDUkVCrWS630kCChhIadG6vFTkcvDhcy5vgiUMW7e64QchCzxOTcGLXH6D0IA
mxGhNqj8qijhvc7dVQqSol+Bx+r5Tduk5X1eR0/tjFJpamdbAfZvsvYaLYwhFCV4
9MIU9LF5WNmfpOkD+heCZwCfNFsgHS+mFg8vNKRBD1eeHXkhJBzYeXAf/3A0EvDx
ILXzvM7qnooDEPKsyIwWF1GaRtNaCkX+rP2AX1BYFO1hVHahhAt8TQZVyMP2fIiu
LJzL3Qd+WE51J8rqhLmXVVHjHtm5Bv41m7f+gw+a9bBr/k2hRD9JkWCtSr678Y4H
eudw1dg1bWt0g2LWotEveFJhw9a4LgzL1OQBMQZtfBaTPBL0FFxMLUvQ6+BpSwdi
kmyaSTjpbv3XxMqrnePCNACSJjEXA5MZ7AJEaF/O2plRECvlFxPNfaNtcKD8/xvp
FJY56Md8yUtk8qaPVJaxL3V+HzR85015N0rUS+fWfbIqRaWbxYIcT2pSftaS8O+d
rkhYu35tK0vWPOn43cwOa0z01c7BGLRkk5TNFrCGbSpttDFFlt1bUnPOEMdCxXDJ
eFAkUupGj4bbQX8imE4IWFQpjvU7/Z9ddTw3NDmEY2NYBtGWYq8PWU98XbmIDA/0
L9EMWZml7LekULADy36bB/8e7FhfL7SwLo49bMK8oXdPlb4XBb2DzUV9XY4Bi+lL
MlHai9o+jW59zUsB0Q+QNQtKYw+6s6OBGhlDpsmjd2bdH89DcRnoT4GxHDLzv1wK
Lr9p9SallK7+pAFLKzaWLC310M7cpB1M+F/8cjacfaCWdlapV+AD+mapSTAXVPrc
0uFZuDVFCdUKx1dY1XNVm8Y7JfYlOB/gS6hUxCkPNc3mMNAJOtP40N0cWPPVZI7o
gAn41duJ9xN8MPebxMWrsDdwWD9DoCubxsqoVL1Tq4ho0e2NjBEmcHLXJLOc7HGM
FXSE7skIF4XjExOjzUsLdNEblg219IMzBHc6zwwr716kz6hH4q65Lz5K1UUDsjPd
NGdk1vuYPspXGuVXDA3P9HuNIGCkb+15x+O1nh2Slf/6e+HQ1DvAVlwwiJ25lMPi
sNSvRVWbhaod/vygY8xAhEeWBKDmV0IRzRwvrvCKBILVitCRMOx20gDynyt4/fQr
q5zdcUCN2CYToDQTnPJ3OGMWb0Hteavfo6sTFTdMo7PbpxEVXsUVVk1LIax2dnP1
NASrMFUjhXBUapXxlHbmap3K53b0TlczTv+kxXwVBWuO1ZwVv2c6JLSrLlwoiPIZ
uw9nqL14xxhiZaIhccRj24aVQwioO4WxNIY3oNqOPGny8NyvRr8hqvV643ZAQOZE
BxGpJQxQiFlGshMnonJkjhjv9PLKAvuMBeFkj3D0jYHx9/wI1C9jrIJN/JCCCeyh
cDP6lV4rZXYporJ+amMHexa2RheAjyGmGptKwJU+mkd8ZsQYFeOX6dw52LI3jYoP
ly30BMPEcayKteUyATvCTSs2Xs/albh5zwt908C0IZMzRt/fTrwAtotv4cJLdQib
Jf+xQ/hhpSOBBlgU1WXGXnClnuERwxf51xBpvgrq6NWXF77ANIoJSIoGhsk0MBUi
0S8zWIc1wj7q/12y9U1qBpNdS9m91+pZQOedsOEI1+GtpAMGVq+s3ESoCWyJii/X
yPB7HOkdLa3EKYjYf2VQelo3cCVRlaCrWXBHWjNd/+db4Gf7Kqg/zuGmIYzIUyU5
IIDgtGIZfvXE6ylyv/C5O8iqqdJTQyOoeUJleUsP+a8YUfLFX20wJs9xTh4p2B/k
aHxwcmaL/jSterjy13cw93T6U/o9Myf25M0/2BNsxEGDH/5QttDnyPpUvF5y0nMj
7wASzDlUXYAsndMFsGcN8IzGtQ1c3tYxycCsrPlPHr8YmVampdy5YiYDuB/ptJ3Z
zrRT2INcLDPWgZvi3MXOIrCNHZE9WDRtbCvTrYKT3oRLo/DgCskjy02LYucCrCgx
zeyV6I9QElcMYFFj0LbmsZrdemlQDvnHRm5i/FFQdxXxTMHFRFHaZV8W8f0UwxAD
AWiApygkuNIr4hfBPdft1GnDVeUKqYVm1kEjetAruH+DwYWjU3VPwfZkATftMHLb
RiqqyiEYglE8yDpqfArNDfQhAIl8pZ+zblf2a21idPGUk5mqPO9R2xAu80P/H2E9
gdwuYDDBsPAaRHq/JW1fFQDm+iyvTsiYKeEv6TPg5hLv61If33c3h79ds1479GeI
fnM8T8R7nGMOCYxgI/f5us2UpzD46Itr3oRK12B1ZvpKr09knDSEnwpBQh03p8pF
e20QrULLa0oMpRJ0KMXkoAae00AeJdzWTHh6RRUuJh9i9dh1Bj5MkJypOYP8oPyK
wJkFtC3RczQWX5O5oJiAvrBbkBZK7BO69zcrLkUUaM2Wc2PTcGFGQ9ooj/DOuiqS
tMYOgtYl8nq1Ww8vmHCsYoHxo6HgMhmGwJoexbb3P2kDMpNpGUYwFwS7HUKDcMoz
z1/SZiWP0pWf/u2vr9P3n0A2m64wC4TNczeLN5o2v7/UWHek0N1YsJFraJF4kEmB
nvl0f/BoAQNQVVvGX38AIq1qMBgqW62s59msKF4qqHFk+6WXvO5eXQD870p3kq7j
KACxYvHDzI3H8eZbwv9bAVx9RFxEeiwpjQ9DTYOORKLU+wZHqQ8UqHaUR2By33cd
7HyOeLBUQpgZx4BNw02ZK/NcSEC2Z0iciTZklFXKLUjgNB/pOmThc74Thvl55UZM
4wI2vcxZPXhxAlQNwgN+cpxF0qhMnzyYZWYgWw41RRgcMCznESLDtBCIFBgXEXCG
B20M2pBycUhS9jWu+VVMpBDOckPWO6VFFQfcR3XZRxYngz/bNDvot/XNxm+clXGc
mJIW5RY95jyn0d87se/vHJ1cr8aIe9F7Jy6TfZKUO6jVstyt07xxNpxczoZ9CcpG
5bbvx04iS9cGezR9LssMt8vD44R0oY+6pG8s8R1A13hWYUAZoNatUgVc3ixwmO0x
PQy5m4Y+7KYJd9dTGI0J4OVwRG2u0FdqPfaUR1O4nDM0rWtX2WyUmmOxI9bFansy
aQ0mREBz+eIPgtQn1rzeWVz2y3Ub3C6nFfrAGHzdB01OFKYQcQ7dJYpS0H/+RXpw
YtzDSRS2tveXqYyLLFTHW95kTBmSAmOu1578dr4mtQXlxcoyw3xUpbCpwCbxIt3E
u63KIMsNzb6fLgypLfrL9RnM8Gv5LblLZcxDirn6r9V7Yl1r1O9aEOuJqFSY1ckw
5aCty5Yx3rqXTjyzMT4YPAp2x0sOS22chGgOKx417Clc/k1nL16uxkRac7CXVGJZ
WdLvPaklTmijUP3juSY0Sal8ATReAZ0l9P7xbCi0Ps96TyRESwxCHn5Lz5S09GJX
qSWspUzGjZ/+b3QzOfQOS9HqKol/xyj5RgJLyK79Gf4x6fkdvu/ZibIFHEc5u74A
vTS+7jFrssx07hZ9k86NaFtTaQJAraeMKBBbDSWMvmpyJRa0gdRPO/a6Uj8hD50b
Krb4STaZZqAj/rVzDMKPcf7XEdxUoqftSB4xxzBond3Y7mbBBP8YD+EfDcxfHhfa
Hm6U/GIv9fIrrSMtkV0IQA==
`pragma protect end_protected
