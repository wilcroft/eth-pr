// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:14 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
s+BJx6rShCKR7n/qzsTrYuuD2KhZAOMtoBkfrVw8FoJAZzB85qozagqhzS2snJ1K
ZqsMAUvyQgJhEViuql2MO/EDor1uHJhITU0n9+7qCo40roEFsZ7sJE55todiWtIv
BLul7mRlpbUmSG0r3r/wQTeIwXFIAtA/RvzHfI+IirQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 50800)
BuaVd8pfUco0puyOBSR+G0EYF3YKfmqu6M/eKFpk246JBScVadii1/FFU33/4Rkq
fpN83c6NYcnUBb1curskajivjBlcguppWHazWtbPGJf5gtoIc4O8h/haaHVXgRYg
1Tf9T5fg0JZasxs19H8QAxz6btktDKC+2cATAWcLBOYmaj0A8O7VikNbswL95Oqm
qWGL7KjWKGA6NKUPdQQLwv/eJr4lXS/X7IgC+/590zcIKM0oQSqPl/1OAWAMefGM
Gy4Wb7cl0DWrg1xcduCl3nOUstcv6/Za0zBVXTrP8IvZlWbdOWKwaE/a3cY52xM+
Jw/w+eUP1sTX+APErKl1dxTRp4fvp2GNqwCVAEQ1rMqyIvGOK5jt63zflR0cVHwx
Hc86b3MQXDSWgO+OOolyaJZFGkbkEfOrR7IBvJFnMql0b92LNpVS6+UyUHjNq9Fd
iOctsoeuNVRowETdDBG81+QhXPY8HrGWgIIqeHskel+3d44voltIeo5wj8w9/jKU
3OphuhvPr7KyygDS6ikSPazqW2xEpfOD6nthLQSSQIulTUbs/B7dRgs6GVuBsFcY
gkDqB1Zu0VJHSnr3stid/pz2GQWRdiIwZLmAY6aPbXoSYhdK2jBGV5ffaI/GAE+G
XNXLUXtXfgQF4wQHKHqldyEjcej7JoB4n1Xu3CP9vMELxaL64VCyuH8iZ9isP9Fn
663VpMiMV6Sp/Z5368NYl2jaHGxe1GYowD8s6n51ctsJHN+Gjn6tgwakNk09nq3e
2wjir9DC7njs+qYuvvuRVo8Nn7TyZE2wVG5/TD7ru8+hGx2B/ib8sXcr6O2OdS4e
sueKFyIPXXqFM0ABNL6C6qH8kdduWSaxiwpbdAB4uK81K8tilMelAiS3aS3Up8rg
4nl7ObCl6vjIuRzMtrWIqG83DqNLREykNvChxeRGyg70e2zP4hHR7WRNEvoSrbIv
b/Iwg+P26N6DNCG4pIsyCPQ6p2vlhxJ8ubc7aUUGUsTgw1h9YaQH8RxLIMFv6hHh
mIbZ5FSuvIOCFIq0LxT1ZHDBkmFuWsld198WauDo/yZjauGrHPb8jGZQkfCvw7GW
aFVgdbOkwGHIwYZRiPbpf+Ta3i/WDo5JkybhiZQPsRTblNoY15o11N3dHU1tG2K1
R3M7RTx4kASxBFPcopgCM0VpOlPma7coL5cAmbg3EOGWvMh+nogLBuv+9lPmQRkf
UrAl70X6yNw/16axFQHoYvzHC7o6bf9ye+akW49MXkDNie4DaHU38J7tMy/do0l1
pkYP6gf5f9XxWMXArl7djnVSFfIbEw3T0KJU1DAUMKM7FpG8fJX0NZ3yaahQIKwa
NnhTA2Km3DGTQeCeSXpfGEc2O7aK3SKo8HEWz0/j2PSRIDix7wanxe077xKJDVHD
NMPmQgJI52m9+vsKq6aE8U6Rz3DhsvKdt6zoa31UiDZ6xuR+xYlJxI3o3f3ZZEGE
gvIXF+JseDVRaTgpk+3TLpD+tT/jxTcJfTdLfu4GgihETid2yqEeT3hOQNece1oI
UxwXINpL2LZN6buWjzBhSj72lP0YOeoT6VVG0QStUMGrDohmfysVkGoDL3iNpbg4
quc/g11uUqJAVcHW+7x1Zkvrkj/pt0XsH8y5ZvPrF4D8uqxBPNH2Z0sTTTtXM80h
chX0L1Bl3kb3RiSkdog/v4RyzyfLV1t78bFSgjcNSeemj/VLpBYShNSNq/yyVi2L
Sk1orOzUcqURRrVnE5TRYtIrcxS8q2HGmUB1z3J/1ghrprUB6XDIPcgy5M/5CIBu
dDyIGbVzLBHKMqX4PijyWvxdFkFxgl30dUIi6y4G4t5p62Jyj2ZZK/L57I8h9ngW
Fk0Ck7Zz5NY91aUPKEesVdtW5lplj1bYl//rNZiw9mVGxtuBuhm6Ivy0Av2xrAF4
D2j7R1OX2ooFsymYouihN3YSxFA7j32AF9NcnAtYxmYmVDW1MpP+hgBQ/vUmvHE7
bwRLOABuyhYeVuuumZmAilU4DL3xhvzzHq1KTUB9yicB6Cmrheuoxefn0TsbiYar
xOabz2dd2EXIrP5KOwqV3JuY9UASz4jrYd5tjF2n1DGgwFqUWevZ2/pexOKU2rHd
XE6cXveWWw56svw4msTCgvT1Kqd3C+5h7DTYGvoH5NMYQmigNHdYkDzJWRqWG4mJ
TL+akZGt/VXhyfJDXpQ2g953CUKTFjofDkywIsvM4WP/4nftDzP6CmS58SxVKQqT
T4fEcopuVw1Qn5PgIOF32OwfY7EupWBFVSGG1lDpbKiTWyyBnGk7wUa6VYBLv2yx
7t2jv3NiKLjxnyUynxZykIODD6GoWjEUNS+gT+KkerWkeD/L7coyPSYF3hcOPRPg
ICmnQL3qev2I+OjOS5Rsk24XZTnwusPSU6SMfVoGU4jI85IFL5W0eouwH7BY9zpi
Gzxk5HPMt3KjGF88GMR/2eMW9ot7Zw+9g7rtVWc+Bv7ehCX4HIJ/6amSYyRkmUNW
J1K0kozp4VKq1UpNZHO3cqnvFBf+vcilmyKeTj64CEWtBMe6sJqYHqGX+HLkIJa2
0RYhqZwJL1STMt8o/KkID6YgrHSncjMvulwh/erhu0WLgOLB0ZHR2syQu5TAj8kW
T+tpfc4Vo4NEppLkpynOitCcubShriVrXQtNKg8uQQ66n/1gOWjjSJrUaOHfaYoJ
4a8k8R9NBeACGs4ajZr15QmLkDcOWVq3qQXKqqJBSWOOU6lcFSivD5Xw8TN+gFSv
09LwvEzJuolSNTW90BFkW+cFvuylexP3qc7q7ti3HrRJGSSS/sUePyVINKgPt7un
cck7locdycDsFlKTwBvhYvQUt+uHUOcTGVqpXfqfpJzVgecbB7yW5/rwBTU8HKQy
sNElz1wgRILkxtonhP29vGG9RRsKLr/5G7WqsBTt6jEUd0Mw8GN2GW1aNnOCwi8Y
IVibD9wx0YYWygcGAgV+X+UoMj4ocXApfKYY0Ru410/+cyP5JuT3V0fDA0qeORip
ZHiv+v0uwpRz+vATKf+RjIAPbbwQ6/E6tUKEbqtOcvd4OuHJYDv9/2dyQyh/+60E
0iN8PcU/pw/5Mi9s5hM9sySOCFPbAWjxaPJKfrGDUCPEpwB+VDHAVwPgV0IE5D32
wpKRgYagqIeEZZa+UhbjexeeizyUCECOaxpDyIDpY6lz4n+ngpmKSTwC4+xXgU1I
Dgemj6PYTZrfwqj3TW7N5dKrITyou8lfQfMlXvbqS9r7UhGxOKlIKZ+U0hbRi02E
j1WWsW6gbrT9Q/6j1dojj+fY+sWBj+h2W1Of09jCXlpDUK/DLcDdq70Y2O1oAro5
JYyEdJsA2FTXweeuTJylJSu7FxppyoM19esIAG5ZAMonEwJNf1n21xxHkNifvmaC
wf4eAUN1UKeWdW4S0jeofiCC7WgEY3q7mfZMztJlOeBCIDqH+5cR0yRqJoymO8H7
AsPB2y2z1RE5AkMVjyyjrAqIUtnQv9qCoVpz7B+TbtmPcYQe7tT4w2hBehqa17Db
H85xXWTdbDkmYl9sHs9cTD1v1XAh5j5kYKHjEndQG9XaeNO1HL0sYruMepUsQFpN
VmdAUXqqsYXl/CnHpk8nhMdxTVvLOUtGnnUFZSuuBW9hdeG5oIcJ/MwKFg2UQK1K
Liy33AOkjoChlMzUAOyr2rm3suLxkpd73QwTYlnburHl9+GTb7HhRWcXJgIsq6v0
4uEsVazNZrEkOSqjqwYLZdL2NMzB5D3DdS4lg53+3s59QbGfsZxa5Oa+Ep6yFauk
VASKbUu8i8w2zsT3BOC8DhratmzX9HbQr4Z80sWfgUU9g6G/F5q9EE6eb4XqBH3F
/YTYaZmSWZmpmCSKWrf0PxDqBAcRaGTu6M/lmlfPLjyHQ+TyLBMUG/Ten9XQWQxq
jQx0+/UxOW7WVM2aKsFOszx3MrYMRnnBaf/TSmv8VQED0dDrZyxYrrCgAHnz4A3n
f1dIU6/L/bdmdOw4/I5CaCaE3ge6GozXZyDG6KAo3ZEEBUI/dUTk1SM3nApYkiHF
0mEj6a177jwhAAIk6RqubOqpG5OetSbDL4zeHRXflkuU6oJJXxmRUO66y+xQ6gEW
b45EIPDQncwsicWrU9SxlgxYaLymfvirV/y4Fcgztfs92PY5kLwZtu49Bsvb5CZC
Tp+4N9B0biShsD5YLEU2NtRKvVT1XRHk3KOQBNL6WgBhnsPo4d835w1yPorYuwr1
LxpNFXuUIryzWKnxyJ0SuQhE3TL0x3E/xAP6/KHvuzft4p82bfSq5YTZSWSvOvYf
P27zBj7/k2H19gHhz9oVVH0ujDAd7IG9h8Oi6Y97wVgK7mcCjW/8Wc7xH+qwrY5G
WvV2eAUYY71gpqSRmeEccac9C4LKEuxfSGcIDoG5ifaoxZNewhfPHOxoa1EkwQyS
ru7KQNHVWH6dFYPoIxmYnequVwnbLsWSNfHFLpODeiV7BCnZnhNVQvxJ5rA/wCXy
tyyl6FG5hCsUuoiLURCppzmn5fYAyxLgkPHPfzg5P93FrhHDgobFudkrDliIlyl/
erwbt2Nf0FkEH9pCxVseqTOJ8LdV3UMfr51XLa0+e1Zqc5s8auelDM6mKY92tQzD
g9GA/966tfhemPJz93w2mbGdFI4Tku4eIuSFf8LnA3vyMTcFGOjpmJYhQCQWMGd3
gQuyBLadZdxNknZGnCZwJLAfU6YW6PKaOsAHz1aO0/JFbYjiuI277hD/1GkVi212
t34xZZkN1NStGQ2uhafe2Q72xjcgYSZJuJ6Dq6Pbs+lKAjjVJ5rTp+o0h5NqQ3bM
Tlzr4tSiAVeZ1i89XwpAINnJiecl2o9rcnKlj4MGh3Xg96Ha8Z2Gdv+TopitZ3J4
rI0Mp2jAmt88pucrO19LFEVl4A/8XEcAfpha9m4p6AJh8MRTUgshib4YW/YNlrHa
AO7XQXMc3Wf57MEUWDtQjaOjOFa50Xmb7qSOSawweF0eGEZSq+koHWOS3fRxoi0h
nOSb2rhlBvGt91nvahaRSmenE60BpFSj0AH0552jrsnWOqRi7iVAeeCQYWNLbarQ
BkPP77kt76ickuEfppbpQYjUkLKTltsp8Mx/x0v8hNOPzfTm4oY6NjiQy5y1sWIa
WyrwEYVy8YdOiB42MZyfMoFVdob3bJpRWDesrdHeE73cETN35q6hNdwyKxz/sG6p
Wme9+RJ4thNtBkJAzPEXxhT8CXtce7D4lz5+vIQLYSPVl36WghvAKyt2OiuQL7vF
8xkwgfy+LN1J8rtoqpJTgal4Hs9MKYMdwSiTMSjz4GVf34RIlKdCo3mi1E3nPxF9
bvy1KAy2Crhj680WM7R+GTUTULGN1pLqEVtiBlEgOhJaEYPXimJClF37X4yKyTKq
qLlS/3PZ5SWuT4vNUnKMg3zsyc2sosB9FpaI+LvFusDZeFsztqF4z5+EqKq8pipG
BPfNaFKeX7VAEefiTzneRXEMLvcx2Bjf1WNINk+P3D1GkaWMVPsRutG6Fz7yBzK8
ctcFpJVOICq+suZAAAaES+8iXEMirlc5LGgQGgrK2mfO27ByhcsjEtb/9uyVHJX+
EiAlY2EfcsOBxwzuYN/XgPQN4lGPEG9hsvsJFC4Js+LwHgkvHFrtDo2vcOSKoXdl
AzAoNMTm0Acrx9l0JZub9dNHvaU4DhlCTIIKgUFL+VqhG2qShOVjhn5dzfQLCfZP
sntUbhHtmDChcxXEL0363yvcsEd5diyijEHib5QVucqr1LqjrqLfzoRPAad9YNy5
XK07DfOQ1czvEyiSA321UpCpiV+lBKrx/uN1/frvbT4t8OtAEPAV9kH3y7ztbj93
ZyWxF/PSVOzbGoFbduVQbmCDex7+J3APBoUUU2b7L69h6u00R0Z1YYa8Bn0oWsXm
ItWRr+2TwKgse2MF8H7AZxTUxo1Fh/f7WaQ2FayXqXcG7guY/OLMaLXxmpJGBn5R
bu0MYfab5mkKEclmK6/wuV+X9R0o6ph+39IW5wcGSh6lClIFwpkNG9l/b/vLeAsq
LgtB2LkuROz5bGsC7wqC8pQa/uedXqnSUUr4EG+ReZlwYU/1/P3HMFzi4W+IZlpz
dUn5DV2QTEjL1IbWNREIF4XZqV0w6tIIw31S14McuSbrCZq0E09S/ogZ7ctthkh+
nxS2k89Z7WE41xNeKrK6L/LFJR+6KW5RYmocIzJ2jz9tblaC+LSji48tCtHacrXY
+uhFIwePoqvgIi4zdg6we6FEghRyxpwUhAcXa9nxtNDUoKB1RaXkK1OEQs/jdqbT
OOi5+oMRWjdF041QTHMID37oq/PqcaMJxw73LT0CDelI7doywBkTiRsP2Z8vkZXE
Qfgcqu+hZ2ie2ZBrXq/0ge3eBQKjY8Yg16ubZqhvsZs0aJAo22M00xJnpqK0IK+F
L6s7BcdmWt4Tb51TnYjjTRfjGA1rOKLzM8OamkX3TfUUKEeyiEdN04/gM2HtRvLm
cWcNo2p668RvOtciXb0V645PPgSf5TKkIqifFyKDmXWCWQhXGNEloQE+7Of52fFd
wuftQageIbtDNwUhYk68NEAhRJk36xc9oIvoOTBOkHDfnWfr6A/Fp5QekgWqZFfp
ibjJPRfdeo68F5709Y4JVOVUpRp7ILCCm5ZCI8KcVrC7exYnAnJ8+t19+ORdzNDF
vZxNSjWnE03amahsOgkY5Ws+OWy/PUfuI7lV/690qLtyZWeMZZZ4zgOh0fIifC0K
pWZXbfGNjedyRe1cOoBloUpmH6huHeDjEjMCcAh+sQnuj0w4qVztHXpHejW02U2V
HoxSZyh6vlMLhCL2tk62dUXf8jslGN1VfjAl55iHwoq1r5B+lld5It0wGc+1NtfC
GImUuaAwuQ59GS3PTpiNzZMnMFUPgnwMGHBOY31WPeFgCYJaP33BAw9Q8/tIHVgN
kG4H2pqwkAiUOlUzSXYE/d16wwsKpiEJyguKmI7Cxw1aLU0OmD8pLB/BD/z+f+z5
PSJb8arDM2zNci3enSgWPi1OTJx8bB6Do7xSuOdI17X9GhfpwAZWUujDZrcjkaei
6tr20c6FzSyijk4a3jXQCYjRIpXAqn0Ew66NUPnTUn+RG1ueadUHsnZVBgGmIWYd
gQbhdbiygC//jfwColfW5i2ATmV456zFmOEPyTLfxqGjqrlvwBSl9lOq2/a6yXxe
PYZi03Uupkj4TyWUWgNz69SdN0EoPctZtWAuh7IcoDl9OOAH3vbarNqzD6IcX4rr
u9jZFxVgX3/nBlyJn7DKRZHVvZBLioSrgH1bdQUTg/0Xdt5m56QmYl15hTK6M0hH
pRCSW88aScfTPqI6d8uVw8iuNeFKkLjPtxZppDwSeNJ3DNXExjMgNa17iwD58Nv9
NHliVBG0bHwqOwwQbQBVFu8qGwr+Iy2XlxRig5csQln5FaEVks38OXC/Z+A4kwyq
KPykc7NJaD/QA4M9fM6haz4THTE85Sw4w8a7vvEhwyYDZ5DCbuDWuhyY/r82TAQu
z6BANUCcd7yKaZ8pedAr0O9ITCZ30/PG8rf5fYtyUZ3JcsbNnIkQU8E6+EQMzE53
i0jDJScEXZWxh6Y4ludgIaYqhjIIrwwYVFmgjCOkfmHz/LFrdoLDSr7R9EWMhptI
Vk9BoVLL4fbC/RgruRymz/7Ws9JYOHHAyjyceLcHmngQ+JwgoT4NXSTqj4SClsot
UmBVJYfkYtNGLV8FbdX1qsMT1CBdKswoH1Yk9M2HEwUriLyVqGC71IHUYRWwBq3E
R2l6G05V6enVrfBKa5sxwtpJe+0/VoE7JFR7HbV3xd/GHjHEmFBYja7KWb8O0l41
9bsppxVw7Z9AyMlVPrUUvkG/gU93JUEC79XOe+0FO1p9YlEurUw76VLTl4RuNsbm
NnjecjwPyuIoP4tMjTFbEMmesU8GLnBD2fLkW3f0Tmh5fNE7UpDrgx8+GsvEj6VI
3YUbar5YrLlOgLm0wvVw00lTuhdj35hY3uNFBiKJlru3PeJj+JUDxftL49UCd8tn
O695waGbIyUDx6X5mqAkS+6RcUtf+aHn8vdOLuymje48pw8r6d1uhWreG6Fdd9u3
+QXxcKkfmpCKCkryzMDeRNh1PqCTTSa/T/YeXUud0+o1ync3FFAuPZdmlNfUM7JG
hTbvN7U6g5U80f0V1ypmdsJxlzLBhLUZYPREnYvPPFn+BTVhoXNEQsyU0X+fYVbZ
wvTVRd72bnQDf7bzEwErLhVH48SEHstEAXFyUdmA4kJZLvHMbREEfZ7lPF+/+6bq
HNe/yWlmaIsc13l10ZuIN90Ca0BFFLckQA2XadNkPzlKt9QHAkwmPdaJvoRAwJrF
2OuOHR5fnKeLda9oaP5AkzwuHA+lt5k+N3SRWHhNQRservYjCNcH1HdiZfzR1pP9
jdLN+srYrp/UzG2hl+lFgmMePJm9xDIOwt26Dz70P2xXLfNHG0tMo4hO0hK29ej7
CSjpMeWi0dXleectfkwQF+/6uPKW2oIBLYbpA87bp4bwFxI7W6J/WjCJaOH+ZdPK
40TC1/WRu0IMjmpFrw/fjNiGdi0DxABico+cClCWOvDg+z55gMYo6iFnHS1thUAV
lXMfFB12pFQ5D4XDV5lxWAE17XvBFlsoUGsFxaRsb2w6IU/QfhK64KeTwqLlhvoG
eZ8vPMkIY67PLGunEyJ6Sw9V/0o9TdyH/atBzfCIvAZepSqlt1koQvd647ei331T
FU6u1yn1ihmXDW0efRK7SetMI4iuGWkeoiB0tz8jhKy0qFkEx3QARAq43q0UeDwR
1k4l75p33PdonZowcWV6ybB6SYsxITBksxmHScIuJsSXRiQNXQKhTdEatZgaabbj
3eJ4/7YoSjI2F4EkWwu/3TfALztf2wMKdLSmcfJA1m4Tj4Y0Su/Wb0AAH1rO+ZEp
LMba8oRPsIMoEAV/vHobf7lGEdKy3TmQvaaRFtt+1zKgotCWdjG3MMaU7gs3qABq
zyx30sqLfghBUGwo13GBwGxXDxTSf3+Lt9wExE/ZKOHBYepDCSxyhbDySTY8GS4Z
//nH1nU22gCzsKkXDywAL0RIli/4CA9y9GOVgKpWPK6G5qlU8xnNsGZjB66/PPuo
+uIO38nTmwT1pOSKoCISHwVBg2UG275CMFrzdM1oEIMTHgXUuW6NON2opfxuwlk/
k03Y1lQQfcm5pLSqLWrc4STmtKvpy5VQ7b+BRgmCkCaH7A4BPCsr08dzKavWXLix
1vIBMXWfGdjPzRlNLid1O9FDgN8VmdMvVlXcBzQg5ng/byA+Y+zBtNwfUI2bjxxx
EB9ltj37/qXxwc2QHcdkGWdij1PGj/lae5CPwXddBC5reqRZLnPdchIBNu7jeg4f
HoBjwyTZeUhbvjRhLy+Coe0wylEe/Gev9G6IR/+nemk1dErhph2ls2qe6LjOwVz6
DtkIZDkju+KCPZq3q/4ZcDPNJVR2P8p8n1EwXed0Oa3Ea89r8wjtDTd9Ggjpk9E/
xPy/2NXc4TpORemTUiH8gEgO5GJBPDEUTdhqW8COF/X9h+rQSnaMj1ZldxzPNyM6
Jxx9jzkwGcjQ++NdHgorFcHP/j5mP63CvV8nH4z1T8dzo70eMriQFuHJar6dg+of
ESHEecr0gL7q4TYuID0MESUklGf62LqBgr6VScbZfI7xoggU7Fx7GgzgRwbkRZvo
vGc0IqJ4xzbaBSCm32XxhyEE3jIf/vqgdaNz6VTl14Rf8wy4SNxaMo6yQqaJBpnr
5bevVOiHEissbC09QONTjn0AjPYjF2W4+F12wGfr0m7NkNilRuVMwyPOZBtVohCc
AnmjDrfascFg275rIPr7iDVuXg0lXpqvT40xBojS2PbVyTPaKXJaPFMSM8bXg+I9
R1Zj3eGW+rZDf6fMY4EOBlE9vHL32d0xHJJtb07LxaqoB0c8vSXT3jQYqaZm1ZTn
59gNEf5dFJUzpSkjx74h95eUKCXzunOCGc5wByME6QlB2lVeXzHjIa+JkiWDJBuJ
qgS+WB4L08ZYR/g8fl39cgBv/S06RqHnBCPRZbpIx0zCrugGyNJk8LyG/8XwyYv9
oiSVpaa5ljQk0u4VdudGch+Ev9iIBer5PSZKQt4NuxeP8O89kBlD9xblPFHO4HL8
bpVO3Rf10UjUUAAtC6SbEPcl01AGfB/vY2jy2ONQ9yT4+HgWk3RRDXBYE0fVUMEk
ZZa5mbk1NOK/gCHeSTLkQH2xGmqVFXfLtlpS9cbeJjA+BPkHcfC8tO3AKOiTE2h1
na9jSOAZz1SyR1LdC3+YZQLOyUjQvR1L/R8ajiCEAK17mWbpz8H2lLdhv7XHTO+R
Z5wtmr2GYU403ytc9cxPJ+4VYzSVuwbTtvrXxdF+kBAbwnp4xpj+jHyFCB63tqby
ULQ4CcvY0oEyoQlbLW1FSeTBTXQxZ58djhh7gbxyLu3TwLSrStSEzDb6TWLM6Ipc
0iO8uxrpVuLDkejY2nAsQNcYqtNDl5pJW3hbqEhYaWPQpDh4RBKdGmG50TOAcbPl
WYHs5Xv8Ly9VA5y6W2n+Kh2e+nqPPzGPhN7eUZT5RGWV14mgD7A0tkiXCyd+++iv
Ym8N+jQ57BF8+i9LFlOI8M/HBlN6MY6s7ilYi4eq9wm5bM93SUnhlNApsWM1OqtG
m3fPzNEu8ZzPn119MTa6ToD1+seKWb15QupleAN5+ea807CfFGgM2nwSnxvUlv/k
JmEHRu0C1MolsMT1O/QpvIZBi/zUP6cZUFWLjYpnqHa8zSr8thtZ1p2whirdtxc1
dHmHUhl29zzhztvsC8Rl6vwa8dF+cpsP0REhAPzOmlZEu4e7i7Gj3Bj2k5McdFsl
71yGWXARauu16zFJnJT74fAQFAdVc/p2deONVkBNxaW0UgjVXKAUbBCej/7e+tBz
JHnn1/33eJxEvEWsXZ3pMKoyVivBLdEeFXfr3WYIY1SQdXVUnBFVsnRFnCPX14D9
VLjtVITwMHRrI7UvHCGY0IqhaPUiny3ETOVoyrNCQEAVTxUcuX09SB2C2OSoCi0J
A1wrjldvlKtk5khgtI3DzrkAHM5g2RTxthQjPtZaMDPrldM1yWo3zPoOjffPuT4D
CmMxr1HEiOthIcmvZTPXiD8mP+TUu+7bVYD93Km9TNRpwVubifsIQOBZaIWC5sn+
4ZZZ8WooIEcSBrcVffPVgRUDYHElKWIS/r57PIsToxOcS89tde49dgn23qAsXfV8
rLf9+rcEmOCkfHAcIUxJQ0FRubcJYHUur3v0gw8FPVZc7QTSmtaqtyNw2mUV2gwN
kwvOGMmYdPI1EsPPjTMBO8euC6dUa9Af4vh3tooQ9OUnTpJmQMaZ2QOHt46mV3Hl
NGow/00uMdnLI451d47PGCDtfC5GKh7s3n/MiUM6TnSO/Ob7/rSmRCUUf1BswI6b
SHtj3HB607GKhUy3daPkopKXi8fehWCafrVwPvrojcsTCwH2flR0PwCWlewHcpC+
S1JB6lyZUMzV+nZLRJ5EUPbh4KMWzDYWxQT0OurUxvzXArXoRCUNs7R0gKhnusLP
XndWf3cbkb4f7jZOr78/LjrHqQlIa8VHhp5aoE5iVRNEEyzC/to9Dkz63NrX9ZJM
+XYRvJy9DNTtEJAvH87CkLvloHY6SyfIgVxveyVfOkdnIELJbulCfckxIlrfEgdT
aaPH1UeSXl5oACCB92lO/j+LsEhfYwEUXT3drTmpSFvG1eQkibGrLW26dZa+201C
QY8MEOzWfdxhrlqTTpMl6t9w35A/X3Yz8gNq+JBmhzSlHui50HFczsdviSM4Ik2/
iwnyo+Zwx6px3aZKTagxUry4TbQtd0+zfGCTBNC3pjhIvP8zLsZHJOgQi/qbdpAj
QlfBPAOMnxxfXRR9oEZ1LvnOH4rRjbHbYwNxe72QqfVibioeltptIcZE2WtbgQYA
M+WcVhz0oj67L9TE35tnNG8IkxK/gwt05aJ4KIv83xcWu9rg9Rdpn5emBdSW7SM1
pphvoq12TYBfRMh1hddYtMPj6tgqOqE8y68yLLJ7a5Ipe1oVdbGmaJRzWa8bEgR7
nqvj83pEcGmUWOmg8Ku5OJt/zDggEakLc18DdP0F7Gp8suNpHfHqjfcLvI5c21jO
O3E/YPtV1AzgrWrzXO9FD8WpLEqzD+7kYFmGRhTj8mqOJzAdpoSrrsIe5ms69zkB
SCEGl3i0OCE9+jtNPI3tMdMlUU47q5vpGbFMqL42r8urBJzj0MXTAD4o1aM+9OcO
NRn8FbJC99KuukrErfbDKJEKBCTCs/BnMTY66UgxA2wXRhwbelKLmq1e4387yP2c
FDkw4Wry7ymG13eMLSsskLxnKVkbUrYHlqZkOPi8fLkl5IRjbF9oPPFAhCbthoXC
A0sMvW6mlLDKqbaYDsUxLFCLipLssFVa+iR1DYfAxvJud6Ufb1XZtX/kyuj4tiPU
IF+FgMVQasG6u5HWzk++BJx4SGQa1atKr7z6UdaKxtP5RnNN/tKNNF+5pB356pJE
8HCzMnR8lLIpl6RR8Q8yzU/4+8A1zOtGajTRDebgBd+sDe+ITJz1yzJm2zzE+yrD
7tP50GS98f8+rC8TZx4wzk1T+ldobZaBd5Z89bReUvKx5t7oVpqM8n+vE/Z8V3zB
RSbpnMkPjLd5Qojd+8wVzflteOSK8qsEa3Z5quBTKPQupVkYhks6S5CqGbga4Ny+
ZxhN9K5IcZ7eF80Nz4vSzbLDUiPuO1lNUKcStwD5vPaxTlZejyGMIY1nRJWrHzNG
MhttD/OLjh/zcua4hRxqfInzyoluqEVQGYNzzzArNvOi0f4GDcQgd77SowSBPnaQ
TOJIH92V0WdKADHu8s09Fe6uk1CHYiYTX0p1dRSRLqIaTsLzGUweLTUIkfKEaaT7
C3k/Lb1gFIcdOCwT2TVSn3FGgNY1J3X/JFIYfFbjVz3+drNXA/iDfpfjW+IWFOIF
XG3bUGMvTKJ5ghf078uUx/0o0LHXSyNPVx+jyecbeak/oKpOjlZNbZS3SKmjxcy2
MicSmXetiN4J6hFH9qcfAmaprQUFP6MsG86Vb/2aK5EkxjQVcC5X+MkYqY3kSRjH
9sroVl+5IC5Cp5J6ONTxuO+FBx9cb0acPvYbPWGGe7CSH8XX6rFg8X9R4IrrCZyg
PDmi3c6t/zkXotS533/Qw8cMB8aYxVttuPLQdwbuhi++78U7Njunp0gj9TkjLgFo
NSuP1nb7J9paug/iqYzT4+iMDODDI6FSv+spPn6vMNqDCViW3D7YsmANqGeEoxkx
RPQU+QiAt/ZIk22m+z/Ga+piEO3Q4VzCKtqQhpP1NSRkJcoD801/fuc/q/ERDdET
ugo5qo9S5JZNMhfxTsXa6FmWnunVltIqL6dscwDupMdyyOfb5vfQngOvR6sl9Y2Z
mVrhRB3h4tuWnweWJCVjbRQbzXNgyZvt+tLdhxXBcnNNKD1dAPxOR8tdB3/XLfcq
oaqQEdNouJPuu749W8KN570nRX4mozkxnyotMWCYyxDAexSNHdtzhpbRutLwSX6v
gJyjWcS7LpJdVu5qs2u2NlTObiDtVt2nUFAsCZ62l0iU4RAKRRhUwiL1G30VjlPp
UEh5jVdWA9cp3GUzyBM9zrj2mzmR36ihJXygTEygKE3D8XiGSL0ll1UROsPj9+4l
hfNQdfs6Lxj2PCgCzjgSnh7yAV1N1PnvXyy65gBqwaIz3mRsRxRoxfHhdiuSkVs1
vLp700mlXW40F8OCO4WHwoI9XfYk0jgM4uODuU2Ds6L1nU5UyOz87zkziWAwW0hw
wQJSORTosG7buZgXKSGzs9cBr4y6miH9a2rvpT6hZKWZHLAKZ8/9Oq2Bs4T7+nk2
q9WkNdj2mhnz9WJfce12V9tP+GoeAyFrSzT9u/uWmFyGGSgJ1PeLz//c2vr53wId
cGg/vidovaWaS5uGqme3wRhbg45WAnfsWHVc4zmrj+3gC4OSqw5WsBSVYNus/jpe
h89nikJe2IQjEf2DZkeJ/qB5koesjIfK5Tycrgs8XWqO7an+hV+quAmFhnOFOBO5
wbwOJke8da88qm1QA6UWeRn6FBNH2be2lhpnY/ONQjGJ+9zro6ToP9ZISjrHp7j5
DkJ4pe8EdP/vKVm+9ELYFFkFvLRc4nJ7z7wxNQa8mHVufsgGlB8chfqpW7aJ9BV+
lA4UNOtPPfXLugBMsoPV+k0NbHjA3ZqFcrOKgjQVGOQBf+D+P8yp57qelRJu+m6o
Jlqj/kNKOfzBtbVkH7G+cfLvpha8PwnGlG+b9vyIAgJKH2PhTSR8lrJO5sc+4KC0
6MUaMN2n2RC5S5tE1PRoPt91ozhPqi1TZHAVUdbwmORtJZaom0wDOnOc5I9amo0B
oPEv94T0CkYuYVh79goHcrQgviMrTCLHS88PFe8stfdrsPGF3lM9HwYQqB11lROm
9yitDepbhODquh78bEYlTJ8aC9GDzJJgzcFOrzdbhEczMcAiLF5Iqycdqlms4PiM
yEECyycZI8sLUeaVX36tbyQXtTavVLOfoTAgiTjvFMSpcZW6s80QYj95A/zOYFjC
Yg2ox/w/9sPNQfNpdOiPIVIGmTwGj50hX9OvXfEUNvKFCNNbfhDTcYpeJPkkPzvQ
48fkznJj44pl6AaXlTxD5kHXZ4IQsTHQTQN/KyGTOZaN27UvczmzJqrIBLIAIXGz
EijcMCQUYiGLVi7VCJEjXogSiUzuidcOWwHamijM8XxQcScwGVxMSyIbJiRFQVPD
CQ6nbk2xtd+0o4bPREkRePvDceGUbGSanyxPG+3jhkrTs4ZVbbl3skYCvUU5cAMH
xc/HYaq634Wy5tVToAzaGVUn0f/ljgM1CjyBeMlzHCBvKjSQDuQN4j872PVpZGIC
Ku1VZ6izMvDviW2qroOhS//SqNcsSVIsMJRf0Sa9y+UwQfjyZs4O+KMX+LTMWrE/
NO09aU6scpgisb1HgzhHR2G8plE8lqZGbBaIeLQiGEcBqPKOIyxDu1650bCK2YGf
+S77rZ7wVNP3lny6mosdLj5Nuv84X2g1o4ZUAw2yjwsNyIwDRm7HVuHKz/AOgeuW
B/Ej8btM3K+UJalTwimihELSw5OfTxr1iAhkw4MYYVjXKJK//76BZBgQDelSwsrT
VzxYD7Q6aE9G5St/sFWq8LkEfE/T5gnAXmjr1SPRBPEfpJ3tsKI1xHBrOOgh5tI9
SqyGMj9odqnxeQD/s+39eCCNEW76Gl9aat1fMTMj7KWnbjttf6XeiXOIqwjMlqxZ
vwtbDyqBpxMboZTbq3FTkiMlH0IU4DYaDiLvSv/yKk/TLmghtK0UvAAqC1JrkcFh
7ZRUiSha2law2beLtkCtuWrRGtugwWQMN7Io6Ybweqy2zvW4jH5WNmwy9CjB2osf
74uV5GOlditt0c4+MctnC/GmXQ8/OYCTZrqzjsghanDJBRBNwmFt1bvOgPspsXPY
ScISegIQdm/Y/UAOr1OpqKu/4mJ36cIx3ZTV9lzl55sQb4KSrHEHo09CGMT7VNfd
yqL8QCv0ejTE1BVIKB9yZPGDvze2mg8GuqIb4MbKP1e5UUJZFoKxpmu32KL1P7of
2qge+MgncUJBTJELg1Vtnn6PU1Yxni5qncB8WEhqE85WkKYp+mm5ajJMQmRfgjQ4
BQtornDFIWoaxcdCMYqT8m3XLZ6X/1t1tCpOaE3aoQS1do34Q9A2BhAbbHlGnHxl
ES5XjqC5s+DJUazj+a+BLyvr1ke0vhUSkwUwWvuvJFEotgDnvZrUl8wsk6lkk/XX
gOw94bomj7A448I40LeiTUCoG0zH8nRZ4JzXgYAboGP5orR4rYT8mCjbJ+EJUj0M
HA7vpxNZl8vaOordB1SvGx553p/bG3gx6NBjWQgio6MDAW4dl/Y9ojEGCa6HPQeA
C1JyAG4OL2d027UYsQef6gxJtbPtEx5BIDvy67ZjP3b83ahVCsNypMSvoOKziNWv
Ew/1gq5I6BOut/8Aka6xxa+LjWaFi3ucDnNFx+VSNtGPccsDhBJ9o7YfQemElu88
bqQOWlFMhYSdEu5has/VLZ8tQuaDPqF1s7JFYliPBArFuoUtK0Szd8u/UuL6Tpv1
b7y1xv9L7HKIp3XhhEwoK65eOEq/xFwROfXMkDGO81jVe1I2NcBUN8n47pZS5mAE
k/JXr9/ZJFFBfPBRB5cpWmdwDdkQyAyYFcTTy4MQJDkflk6xbNubCo2uD4xaT5AG
xpSiCFooKznJla8FItLspL+qGxtpY/Zd9GSAyyEUCw5suV4tynnq2+WZYAfCk6K4
CSRRnUAQdznwvfyZim2vA+AxMyYHFODs0GwBS7/aKPchr8WTRNeQzC/2RhA5B7cM
+iuwOhuKeSg7MhNWz+ldK6OtbKMNuDAtlBITjiJQbNnH+a83phua9uusj3Ip8nKo
Dsmt3Sv8zu1kRPXv5gvc/xClMybh//41P3vwhDUytG1jVy2kYVY1GI1f/2SU6fBI
W+RcQa/uCAWYMSrT+4X0K+mPmpVXuwgElqE7a3MWGTXwb55fXGvM5ud/Mfl/moH4
v9FgvCmDrhiXufeH1B2N944nDJZk7etS8q8Q7e2uZhYu5BlsVhV+uE44xDL/DM2s
v5yqduuriNv5kFpaB/OU+lCSNFQXMkX7Qc0TpY/0wSVJxh1lQbem7qEM99SmZl5t
5Og8gTE6izClhNPn+DCp6X+EPFVj+MAYpRIVQXLNOAHyDqHJbcoZfcnntyfr+UOi
Sn6+uDv8mCsgBbbyxCoYLDAIYX/T05H3l2TmmW9kFPuzLrGeJLhrLI2OLtERWMDV
hV/wdDTO3DBtVad4RbW+JyISS8CX0p9Q9X1i5K466anFHbG1OW8U/u7lA6XcCm8/
lujD4JnVHtos15PNsmmXCDGsDZQfQUR+uRzSO1p3FyHt+9eIlwKhPJN2RDA0NxGK
ROdfuwPiUWdOcRFt1q1+bciNz6W6F4lkc91AdF3t+v2ozJe5jgAAXGPwWofU1abF
uu9ZJE4tysFg5lFQziTUSC5vdORDPy9k3A0FLqT+COPo4NDLCNJf/wh1Nptitn2R
wSuSsSwFmfwsMr1Dam+RQj9VmjH9lhQxW4fBpvIeLMyM481msDLd8PlXZLofcOIs
hDMQX5qofMSGQN9FDbPgB1IobQdEKG8fb5gIfOscubb/YXVFGREk3Cjp8tEecMsh
D9X6RkFqhoNt6OL3nX+jG437BpUV7IotDs2kLPiwP1Yo/Na6UQZLTAsx9yu5ABM3
WVT9vatR1RGsCH7oVtuRoRS9G4d9Ov9+Vwjn1QaopFL/O+/DkLSC+PEPZai/TNJB
vC8c9htVIy1/3WK92Nk6YRUQKRXAx8Gi9qZE/ruPBSThO+FmaJ3MqY8jLwSy74qB
AHOSkHibv58AeIuQgqWsPQyHW/kX9aim4Xc3k8t54SkPux0oDiw+AloBPMR2nQXT
MwrSLIzyj5zvTeLG20eL2ClweqUIvbeW/nhMr4rBtpxrWX+P8vyyXBz0s43xG3AQ
UDm6N/VNubYcUf7Z9J891cGfZfXUwAJezMMTEYkt7VeqN8xRqL7/n7FDCpMzPDHP
UKs9iAURfDhrnDC4SURKznnYkJ9oeuSxgYVsxqOm09brLi+2UnYVz+igHzd12yqb
qKJDn8StmUyFqGyMWprmrU8t/uFzSgm7X/fYVTL7lwaxWCxDun+adi1u/qmtFx/y
oi2KK0pCZrTtpNAg0o/D2ktr+OU+OpT8U0ciebowRWCnmzoyTbsE9OcmH7ToNBd5
H6uiIPBkl5187poA36II/7Iuru6y8XQiaxATHmJ++8ixMqxicFmsWYg9A8JefZ5P
Ff5e76Go0kvA7R0529qaAsImLh6ZOgU+znh4SZZ8ejrwiRJ7Tc8TMeLKngw/UrTD
dKopIJjKPpnYhdDqkJpTxDZA5hRJDgWnG19Hv/QAxJUctpx5vePeTFtr8xe7LrjU
8/45nkCNko5DFlZZ/wFyn5GsbW1j3alPXjjaOUKmJGCZScnX77d90BsUIse3cfsD
z204KtUDaXWyCNMXvPA0R0BGpqEsFvSI53+uB7hIHZr6k5rcGFTrwJ7mGmb/1XMp
LrQRNFc0EcubVaP3uz6bl/6JqlFF6lEZcCBDmQ8TIamzpExAq5ci3y2Zl4vx6gBA
egNQGtP2/6U7b58VuS9MIG46Qq3Qez7TsDV5GM6RlXGtOXXJnIqRUX1O3A1gcItE
TLUKl6PoFK2rxgDE4LydnNU6lykzthmPpJ0w/SzLOjCrcdiWPA7odudcHjZaaSmx
LJaW4Brq/JdMuw+QTIpppEL03XTgZdY+FCKaW3dphiNCn2NtahjNIVJOfxgzva+w
+7NyPvh4pWu+XfsfIvIKII7RDbILs4yKU0iz1oSaHjJz5O69wenaSxokERvJKgT0
ijSq4DOqFrxAuQLVl1FRPdixBmJH+pnJLoT5MaS0ciZzTL7VvUmrAohLPbRzzSJn
vzbV0DXYK479gSkxkVJQJL417bsVtkKw2fvrWpuWqgi972bzS/q5bVcCb32pLEF9
zX8UdZaWJj1GlaGYNFfW1rtAot1sb6/cupoPUkpNrlujGmSNZqB+QJLPWTN3xXhz
xQH+rBH2L9mhMPMXW8aMNsKchOH4fgoyQJW/xPjM0P3zOWc9CJDrjHR29COgc+pj
PHhQ8PcIIpb/sF+Qwxyc8Jsj9uc6zjiPKgioV1DOuoupkpbxaUjrnIAxEj8jeSXL
fa6KDY1lGBBtSS3CI3A5gxbVbFca8ZVIVF3ilP68xY2898JK6vGB7IsVhwNttFs3
VR6NeuA0G2NbvDja7RBs7GRW7dDR0kwS8iwcvsRH5ANhmCri17YQhN95Vsj41B+F
4BMZ7peP98Mhn7YJPZz7u8nbywQf+mxz9PFoAe008pcHjdL9Qc4v4nj6awJqYr6f
Y1vcAlhSvKYnp8kYiP5V13uzJ7x4hriWj1flZcwJ4NsLShLq0ffoC+JPrWe8E1Fs
xTHGSOuopFgCvTH6m9cFACWdYX6YNog9k5bMMf07Sb495IUivz81Agg2nMLt9GSQ
c8ttANy9ntntAJxs+9Zn2jv/l0Cxmd2TVM63Q+XIc87OACbDv+uEz7vXPqhT1ce8
K81u/WaaXiwD0RuifQh8u1f57Q/Oeu+J8Z1cLm1E5/e0JJiC6sRydFuHZ0rOx/h9
Qt/mk88euBLgYF+IO2NAq+1SdS1t+OmeeyMjqs4biLeYS7oOXQYeTEosfZ63ziku
U1tmMh7KU/Mmd2wT9YXB4Y8KsvyfpFFJMQZwQHPLHZQieDgdBdByVIuB+Gt3oocw
JOLLLnkl4qhttDKTVXuwxm72RvXJVhqrLrmH9vRKwLrKRJdsancimhj33HpTTHq3
96H69vG78viZWpYE07Zl5IeHOGKKLp9l2ymxMNlew7/LkMfsbfy/mQ/t8IqUgUvk
Il3TKPT2j1oHgylM2CqsS/QmS/yQNdofSlWYpbPyJVctPv7nfd85kbLsP0OlzYZY
KpaqfUjF4KjE0mggDYxwCpzW/a0vG5cvXlz8oKLbDyRHRlyqV0XpOsDsbeugvLfJ
XgJmDjh/U9PKY6KDgIZ2IRQUzb+6I7ESw8sE4JQ5cy4OIJ8UQJGMbwIAR8j1zVIH
3Bcn+nEj/HPq32tNrm41rx/Cd9Rvx9WIJJMegP3f9jJCyLW+DAh7mEfgbnZsouXH
CvlngO4pH+hK3FsLAamafByjF2osJBzIeaVfMYhrDuiia/KzSDk33XqicMenUVc6
eOsTR1r+2ZvqCGa/9h4e/JXMBzsMXa0szdeGd4GjV1C27aKHFv8MOCyyb6lAArzT
OOW1uKAkA5GkgmE9OcwkNSJPZT5H6pdFD4urPUvdgKeo9Pi7HhHES2745zrxpoRZ
TVzcEcAaNecYW7zFYyzA0LJpxJlb5MS2hPJ6hJkjLYq1Xsn5oS7XcNhUMRACuRWf
yZMENiJVZDKBXow3R71CEasOeaLbksdvbG9a5yCzWT2lHQJ21kbtV+3LNlmiGqzg
eQmlMfynlSRfknz39I4ex5TjU5N2699cAMBnnsWayf8D43YXv3m5guo8FBI9ZNJl
foXmTUKexcJHiU8SNGqJRoaKEMgXVF43qSOmQR5wMCB6lA8TXyYkLGx/jT2MI5NH
DSP++jikcJULrEN2r7ZzgRHIe4DC2XmTv/0LqXtGcKF6xJLCE+49V0UmuMGpPUVx
7KD48+vCx/5IH4iDtWOTm40Wle9knRFjywvN1H5nFA6/ZTt5ySbmiPuHm4yfKTkj
Zi5X2sy6Cx2gSEa6Qs8+gqMJ72Pr0YHz5kqRBk8wlQjbWzhwFIj7F4NDVbrqZV9S
Gp0V+Ro6ja1oUq3771uiUEKEsNppat/bzVg+2wBbXlxOcGVWcOw4RIvLhs52yK6V
+4uELmoSfrcUGDqvLbvIatgp5HDNcF+CI6e837YiG36IaXz9UA8tMjxr31tZetrG
DdR3a9Trc30hBJpHtX9Y/E6CPQHPHi3VRMl+G9/aUQNj9v/8BmBpB30S6mCf95qR
fWXkcL9qN102OnTi/GpDhQi23Qioa3GCdgu9zCl+ETyfvR0k0ihxGe5Hqd75/GCX
VB3Vam+ecncIysvzxFU/c0rAKGszXtvMIMqeyVcDPsBQjBWn+1ZEyuiTFXQ4HiQ8
CxcJiINfb1exU6DeT991KydxKA+apFF/fPMBRSgqykW9L3HLc0d5uCGwMNX3iyqq
qv83vaxeuJumNGgh6uT1ulbcW8U+2hbKhp0D6Weec7mdin8q3RZSnspuvL2lifm+
WQbkX6lnSF6QafTLLeIoor+SQmiKlNBwY8NxlL/hcfQHI7XoWlT0Fsq4Xz404l1c
5x9kelz7Kri42sSnkYk+a1HmCYLoTWTCS03RyTOfCftjaR52dFZWX/3rM3T0JvC4
3zNmXYvmoCM445yrGuEz9j3WTwfbm7sT04kaclfEFjV5QjR/qV/jV9FScB1WaVXL
hbRZ+rAa2Bp173Spdq3PkmCaeeCocXyRkpcAqzqqwrqXQIApaP9nw4NNWTz+IsvZ
DGJBz2o+s8H77suu7AWM6jzm3pzX+v5yO+eWYRwvXKTThOmAB897dvH3d0h/ober
O9Uo1hLBBddOUT0kF3CBcXCJeqieTFQinU+AZI9WsboHm2jSyKZo7J7irSZIXz6c
Fasd4B702AxGAXj5YuGzjLJjvyW43ovlOMmxYqGDesnraYfQSI0edpE4KslJMyMN
PEdgUZWJCBILejNHl0nh4JncQSeW9TgFyNbm1f452Km8I++zUFvXkWWQa/yPqP4B
v469dypgLHdw702iCDTPzk0TwGhImMjB6b+cjbFLuCHhTsjfrDrmHDrmc184Fnta
f2pZoO3lXqcQsnS+4dj3WXp1WSIa764iZE6EvWUFjdYD6AJ2B6EkVygbQxsW9BSq
h+56JeG60v37oHoR+UCSuS+wkFfg6Eh2Var0Je3RJeusPPPKfnlB7oek6tSw+M/j
+aozz/nvn5Xl4TyW9pBpk9ojJ0Wc8oyNFniMrhSTlTYk6KUwJay7vG48Cf8qcnYg
qJc0zxr39b3O0jTIVO8zWWCsHNsEqsnD8S8yo2s9KFNpa9bS7vCiba8+pF4BpS/h
n7k1x3GuFoNWiVjCqpmsnaE33MjJ+4/FJ3rklgGAaYoEegEqK2ySgEIeDw7Pbi7I
DXdKRHVuRweX3h5JEZCaFHV40QLKinuO5UI0w69FLr9fL2Ow2zOfQ+hbE1VL0HjZ
2QRa3sD7Jh6l3KU+Y8GFOolRhLizJD3w/HzlWw9/3EwQGnJqwEIXMCIF64oCrQc1
nxD/vPq02PcI5mSCM4eDc2Mr9I3wq6oPU3hNloNKgJ+apklPRR6vBJ8PrSu/a5BH
1PjGThi/3kMJnS6I+3ibUEfYzgk9K8kJ/d3+7NcnKn2K8zHC49UGrpOBMaY/JP+i
gYLDNvNsC7JU1rHTSuSlJECbKqg38hVF2po75uQ8Es5TUjT/8c9ua9FlHAMLzMEp
iuXroLw9Uxw/uLWRWl7NDvs0sQcpz3AeZkkZRNM6j7pLnwlK7PunNb541WGYqIx8
PU8rRWJ9nnPF4g2fdJcWrpsIr0komuTWKRYvtChnUtBWiCzU+2GU+oAnLPrjra3I
QKSFFD4lvCHIK7dIOqXahJOYq1YJfB3P12FZLtgOwTVqkAangywJ4JNrYjAabfVq
tuP7sgjb3jzzaFMFN80NiOmC1gXXyBIbJkzlNhNGwC793SHjQtOBeNg4Y9kzC4L+
JQT4TkDL9OQM2oricC+n9ec0vuShwQB6SlIfizhO9G1yOnrwHGWTQnX8VgPcUjoh
gmqr1ZemeJfFOCSVzVCsYX78kwe9PvL9VZAiDnsx8+P3UQSjBeOcjazk5W3mn8I1
R4+QexRaQc2Fav3v6D8c8ddQlDHNJcOaoyhLcBoUy+v9g3Bd4jmXpi3Uv3Uo93DE
Uv5X2IGFYSravK6DCOEbfgUDVegEVI3kfUpzigj6UQhcc8Fn8DFSxSxHfab7EqgU
ZC8qExAJm7ZNvzUJ3kLD+mzOp19kCeXXV5zCgvE3+Y7dYP402Fi54PLSdCKmmE36
9dgMVHdwo1GCYfDfutLb5jPFYuQZSXSIF4uwuw5mJzPAGJs/q5g6k9SvQiakSiU1
fmXaF6cHbvkoBGaSs8aKobmvi6+z2uv9M84kybsuLT5qp10nBGAqu4gQ3oKy7+1O
+wlqFyF+YdcN6Ht3fI5Smk5caOu5WKuJqjWitznv2ufo0ROAFYklxR3G7XFDbrzc
N52j/lgy47GwYyXV0OX/izEDc60ZdJTHIe2mlav/LU2xsXrFlHeovk6Nux0s+r2a
3lZYYuWkWklVanBdj2iZvE3DerG0r7F7DGk3qKwxvBFev4k8y4FJ/fEbTCVIZ8Ru
bqYjkvJRRsj5ELBKdVsj8g7bJTJZoh5X2UTDSI4kfitFXgoKOQ0BjrFsCnFH5Up0
/Vkn0OukJStboF2lXrtfAvB2SKsAxCkifn7kVsKtNe9LAUnyvJEmYCKmWH4RBtnH
61wh/wLY8+sbEAaxVvjCDhYOifRsoLFPAgbWXrM4TZTEAUXaSXGA5ccExWE+QqPo
mWEAtsWU4rDyqwpw59hX0L1nRx55Ghv2HMrfEUdZnvVuySsnygPvKO8M++/0BOND
bljk/YssjrUdl0snDjHwWC0pG1RtHcmfj086emvEnKWtwX8KERa0dqnwzILxHMQN
JN6YRa4Qo7oy985b/8T/DdDDzQyp64Q8Oc90P5PL8SO/u+16v/CXFL9zEvEAfQJM
eawhGiAu850RW+YjwZSIOV8rjhtJW4NFM946Atd+BbuwjmLyxmG4TrIaevjDvxSY
UqGxr6g9ult4uCyST0um2R4x3jNkrms//JqT5PifV3fcr3cFjcKmnhWVTYbtRks8
RzZhNE7wOgoHfeZX+v6PqjpunV29qIeZuCeY+maS+lFK8FbxniODiYG5WfTK5VrL
y5FzcONTByx15I2YiZRFaiUPPNosIQ+x37gZzcIB7dMZmizWsyqV6WkbTKw6R32l
BI4o7eyLm+wEnVf8qPR9lcH3aJsl6tl3/5R3jDxaAKhgtAHcJNAAeqlOJ57uGyDP
NsoTACAsLGLIWp1Vv8zt7ndaZmWhmmlP2V+m+nZc3wOOTPQpk1b9zbwRl7J7C8tK
GBVMS+VKLWwbHFpAHjrQZ3k/jq72geMKX9Y3tOmgCTPyTFfJVdqXTItT62vt6WZX
RLipbyTnleLdkExhij9L9iz3Kd7Vet6DYmJZd8cUOxk1ylsI/J9JjOA9FqsGnjqn
EZ2Ul2rAe/iByYDWlb3WVRm6s2Rk8lPwShSL9Yb+tW/E08ksTacw8cVer51e3Vv9
9s/xFDJK8dUGs1bX8oP/D3gt86KIhaqvxhSIn7Rotw2p0AJXB4NgQFDaUXUO5PdR
+w25E70a8z6QyhDhZV5FjMJXJSVCZjTiHBHEYOBrcCRQKEXz1kAQtXxAGCLe9Nct
z5Nk8Y2C9wLVwthQYtOQrZw4SEb8xNri420P2BMtjcytUnvwD9GpNrK8VR0SC+Mg
xNX5RqzLQkNPGz01R0EPDAcxQ5WZ7JL4vOxpP08tPd/QVlDqhl5U93ZmKETz43qN
IgiRLbanBdgmONOyqqTn5ZkylURYJy/XIzqxbKLVnhPaDAz3bSHbMl3ZT1SzIHDY
m0+C7DOLmClJeGCkkHwKpFvtsP4eJ402BmjRN3mu/3af+vvVzJOuQcG4Uh4/dCnc
Xv6XEro9PthmUNJ5kViDtLWg6jjFy3Xt9mfYqSPuQboGawtGwHhS0WaDr0nV1Poe
BDypz5F1F7CNZM8IP3ivZsby6Lv/34jXPEx+qFWEvpn6YZqmziEIVQJux0gMthRQ
978ioJdWDHF6S9ebv0EhmueQfApDZ0gaS/y12/ikNybWN4fc0wp5UiaV+bcIzxSR
9a81ALdzaWtnufl1dplMmEUmQPQqy0P68+FnObq6lpbEV+7ZvT8LRJ0YLvFCKams
kLM9vwBeYkgOg8pgueDfv5ug1spCx9pC4Ld7NSgDdBiWOhimGRgV1fDg93wQvnV0
zkqNZ6y+6tdZltyIxE8DKghldV2eA/7fwr3i6oU29iuN1VXt0CTbn8ShUoDvamRV
Dq0Xp6nwOfWN2YS4vgk+OuYtliw2T1oyqvRELnnsfWsYEdWXLIFY1OPPnmHiQESn
zUMmtFcpLOpHua2L88MiYOEAL/Kjkxp8lkJ7XAZa/vPqOq+NywFrHXF9n1p+a20B
STfpfwUtvVOFremPlRfs/ujEHvYmCY5620PthoP6Y1m/hTgABPs6BCwAFdJF2dF0
NjXki+WqXwy6dx/w84uuCI+lWhFKnn4hpjmCOTKdRM7bE4Xq4W+omZbn8F38gTHv
9WKb0MIEeHbe52XmzEjHwSHrwrtBG1GnJAM0/9cVWPoLbulSneX7wA8Sw/p2mCXz
CkvWKyjq1qf24tV8yeG2auMnUprCeAbaLwMneIiG8cBdTf7eABWdbae3djwZnMuB
PhaTYn0gMt8h3wL9DYTjYJfEoGy3KlFqxUZjfueo90BEAtHAfeq2QFk2TatmljLk
Z7ErTdJRlC0f18jq/LgaO9AGKQSM5pSvYhFnAanm6mcuolABAvO/tBNHnfC8TwdO
EljhoAVL8QAynyIjpMpI6pEglSMMbRnRBPxNwueyYWBcxsIRRAk3UTw2++qwTaNN
430pomFAbrlWAzi0giBxfG1N9Dtyd/j6MUIL4vLfwYSa8bdSOjeBXtc4XBduuZj5
8fQ7heqCAet4VyeoALRaaD6pOF9myGFJt4l5QR147+Zd6rBuvZrBSxAKTMFe5+J6
ok0Wb8bVfNljr+TO0poWN/0HzsPhuucaYA4tOVzLBXrXOc9uxXYI2Jbg1n7V8o82
z0mwBgLUfRU/Q3XBtU2j36S+dEVIG7WciCbT5OYCoKJ8rVcMd+nlIXLdNC/SNlPy
rIxEdOGPNYImd1FYbI16YDjPS6SJ5B/OWpnzdy0q0vFMTiImp6cD6dPlOpzJruFQ
VcgL/2HqWgpEVTXUdia/ZvTG7YDv2WbuBRcMGW1CpEKixB9Fph6xcW4Lgq+yvtzi
EMkI1TsEqcwfSFOX2DG/n6c8piM/EyUiOwnalGlZdW6yNLeeW24CjootqqTBJIS8
Jc/o2WSABRIx7O5IpVDyOKI/mFgdObyGRv677HCNIKNeYS0MvzUCEecYVEHwkBBs
E/Wk2qrxdlkE+Mie6JWZKvn3oYmmizoxvY3n4DGgTzjCFb3HYynvYPS/bsuEiXp6
913+XIuYduE1iUais8H/64ZDqSi7zW8qrgFITXPF+h7MNm7FR7/Q56Gjcnn7DFvQ
8Pq9Vy3sR+W9fVP5iDNeX6OcuHxtv6UuCVMk9r4+s59wBokhTfvgdw42qGo1h/Gw
c9+qs5Q6f/Hd+/7l4nrt8ZdPNwXZ83raHKukc3jC7O6NUobAeyOhajmOlvBaXD21
XTBw8aRbIMQVIBNAXSeDxUIRvL2ZjkK7VOulbBlTlnAxSX2C6bQ468O1J2hfJc0Z
rYPyW7h/f3oq8g4f6iigCKHt7OeZaGXidUlKC4sitKQjt42f59i0Q80CFZyYtciZ
D1iQ0sU7OF7cERiwaX5y6z3mEWtUdcLCOC9N/e2USdHCDbNHt3LeNAQnkU9ZcO0J
wK33LAx63Cfers88xmJSb62JHJmDWTYtJsic2+XwtnkAhU5y/piyzjBOb2i0T3ok
XmQkq0pf550l4h+jh4SFWyG7RaoFTSNF0ckTssSbkSXxq604Fxw1XL8IzSKAS6TC
nuvtbSpsvrMqBsensa+JXxUid5+LM/PxW+mOTauCSmHRPWo2O8P/JtNAKEPIkO03
bZxC8WxhGKegANirlY1G21f8Buv5XxDIHa+159FIE8W9XgybPD9450Q9XJBUbc0c
f+qIISUK2s1AprR4cdCr+S4dNNR9N4aVJfDO72vp3x6+pynMq1TseeOsWzbgUSf6
zCqldFiHniDvXLwoPwLM02HSqkp4DVjWI2la1lvhrC6mJS2ZAun/TCQv15gy4vGO
iKsAQynY/4uSfuO6JJKws35ghiN/hvIcDuyfrqVcdkmqj1BV57nFqLYOzZx0V27h
yLw0iMx4426qC4N7aUF20BsuC/aL73FJSlFlMCfIU7cS2A9p+z8b+xic9BikI5JX
dGNPhwiIJflfvkck5LqqfiWgRwGu9eNk56v0FPT8iEXHlT/Msf/6LSpkJJZHh+8E
b4nNzCIYfU0GaYL/AbidqniGkNs1VU9wKcPLI7VD+m+HIcTV8uXDiXizBEQfx6IG
y4A5AXAE+OhuP1IKb6Lb74ZCIv/p8pwHaPfGwlMt7ZBe9DjGMxB0VyiGm6+Jyg7o
DivkIaiTyT463xHS01lcht+D8kt5DQ8dbQwv/H5JB/j3C78XRnXzRY34SAyukc86
TZcZNM0CySzy6p/nRLqkH3N1Of00qk00o0g+b+9JMwJ7Sad7Z08RkjWC3hAHXtSL
wa0dqfuMgqsPvePKA0LabMBjfwYNP+4OUYWMb8sq8/qlsb06L4Imv6wV56wB9dzQ
/B8iCjksnRHiC7UYoQBpxsJgMdiBBNeNNJba/+ODq3q0jjocAybLEzT8rUFASjQX
SNWv1c7VDMJ07S5rDfrFe2XzdSMHbQByl9q4TcOJDTT/Pk+M9IeZUnAsklGA81sx
ae65EyzhHgdM/cBOr8hd4CSxwX/IbwNDBmKCWXOTaFJIX5ZrxB+QB3dneKfN9yuS
RREmTaEv/wuHgepqXlrCH99+XxAAOToktyggWNEVMUnky3FcegefSCDHHdSRwXMP
SOr/0F3FYx7I+qozoMdhtmGLAE1tYFMsuzy6KFQfq9PbJfAjb+6rBEK9fQnyXb2f
xUdIUxsT7lIhfR9mtceOuozlCrBJMuwnvGIP/NDqe3bc6l8LFloOK6y5FWcWFh6h
UX97Ajsk69i7WSUXuiU2jWr4EZjWP1MwECXPTa0adxffp6MaknGPeNMxJEMFEpSS
GUci58pW5XNRtR+3FZgswrCBpfas3JGAyE2VqQhhZKrPgyJ/E+B5XuVy8Hj/RST9
pIw9sowzoBX4fXzO2jdUsVNgK685rk4I8raBCoRl5vzN94LFWhouj0P+cHebyNrm
2vuQIs/dzVEqq0Gk8hfo9yA1ArZwJgKMVwzCMPbu+0ZNvL/xsNOC8l4UJ28UMglM
c/vgOUlCks46u8dgH6YlIcNdrPeqVeXKcgFyrrpNdLN/es4yBhAsDXZJ7nuNW6+w
gsiWWKOQoG1ZabvsWAANtaWoG4clR9dG/bijndOl+xtVKFoUrLRhSVkQQpHqN2zI
eRmzOiGIahL5+FuS1Z3As9RU7Abdz7vc3JVAoDeJ/+UftOS+vTDZl0FxhRx+EsZZ
V5wkCZakt+nswz9v02ByN6nvd2h9KAQUGOVEL39WRTiV65JOsPtimiteeiTXRKzv
6BGY188kbzHCdAmLQ+LXchlVpQJaUx/yx8gL4WCo0n39Il3LyQABAo7mAAEUOU8j
k2bHaRP6Wy24xVgbgaL+mcKkGHoBoeQv9m99eqbR5I05VizXIhYhwynDG/cavjgr
+sb2OZSPkljOU1WmjAgSITYDvXTgrZLcDkcC+lGibGr2oN2O+5X4uWfRdML4HwUu
9HgWbbW3eHO9nrh/W755OurytZLxszVyDbOtl4BXp0Ps3awymxv2JKUS/Xg93QmM
eTZNxlnQTpTP+ZjNwZc4MY23EZ4XslIxZhvQKSjRkxW+osYHS6iNJNJk7pde4HO8
IvMZeeLoT5cgLke5YEKEqtTsOYAXXG/nm85IIAnDfGlTWLpqnIgIALPUmEV3Dbu7
MYaNmjh3NFbEi4W7sn/TIF6f16V8h0w/Het9SbMEpJxsjyhw7PO7CYcrpCgRLRVI
8P1z2qH7mykpW4fgcL3mcNyirJTh7jZBwhESQRnbeD0BOkccFDKu0orZJOUDuxZ0
IMi0276uPSe7zOAt7r0xe/xvJdxr6zE336g1OJ5t/SRN2Lu1NSmGQBlHrH0hRCo4
Z2FQ43H1G8a62Qy/eCl+QiEh6jjE+8KvibF/gxrIwJTRY5q81lEyREFQORWuo+TZ
hYtUP/paD06mhOytOh/LA62A9CuiYRWnaOlfhfDj20eqXV5XO7sqz1+p0fk8MUlw
6xyBnkT3XSuX4Sqv7DbW4rI4lu9nJlku6XQIsSLSfwq7bg4UTEYQb/NO52dSO2sB
ZR2RYMVsYOH+3keOF0Jw1OTrYOn2Yxyo9+Q8dGGtVCAYS3Bm0vk6DxhvBi/jgexo
tCNEDpoz7S08u5wOE4nqxHkEfs+HUmZxje2M7f9+l/V9IGqj2EnLMt6+3hOPQw6E
ly+H8glLC92pM0C5K4mOSwAuQCrpFnVRsndnIDSxxIQvNXeq+5ENQH2BmT3XOzox
PR7VEGpP54UiaWLG5R/uGH4ArYXm/dQ2oehu/sT2A4t2Z2u7WfAmz0NbEfV7By3L
TQbew5aZVrBddj3ytEuC2UNonExvRc4SzdS/+/VCHEfglczHXk/ng6v2rR2/2Dql
GyN3R8Mmc150BoXtF/N8cezSLvCVFDAklNJN5WZLnuFJnvILYt6tCg+yT9g0/wjk
mrCSSXBW6p16f/3/VWPbcO/9AsjXaOwvVucQav+FymhTlCOsMHDKiXJUhNXWOxBa
La6jUUZWCFJmolxHrLlbbFIeflvc3o3eoTgX9teKUrGdGl0uFIgdbBQQylWfYbtY
IDmFD/R+drepBXCzjQ/47xYFgGkwWpQWOk/5A2QhdgGnLSbr3NHXVI24gfT0eckt
+asFoywdTuaLzJNMYccKHAtmyFdOH5SBk+3aMdsAHnlLxoHdIwZfL+p1XRPaJd5V
/8s+PnQHf3+G5TmhDBngLOcF9hp/DLUntT22a9FziTGEd7vHcNy4OwhCvn5Wv5cS
qsFMr2W2WnJXx3Thrl/FKGgVLXhAifFvSHgyoorDpPlMdMfY3MayY3vUnd2lpmWo
84WDkZVTp13TOFrbTDTkhIBYPwTP0v0yb4sIsj9wQ4LP1i220fXiJCwMsATLO0Fu
Z0/XvuunBSifzunguyahXrpy2VD4z+79/VIxXYhpQJ5FaBN6c1W0bZT3EBMZh7nI
6pbyJ5w+WuRhtwJlFP4p3kdykbDl5amz42OLF1Pd9zVW2fA/pRRhkg7ZHQ5SuJQI
6JurjKr8NjgiSYHoOkB7rBV/Bjtsk+kTvfEFFc8aWB3iU13+uCjL6AAB1Da7LbqW
tmHAIqfNT41ZezjD1E6KD7nppBwYf1qWzfJ+EgfWiFaA3DvW5qn6K/wbGsOVPPMQ
ABkIF9qWloeZk382RmxZh/SU3CxlmUz1aBDKUgmaSFF+nbxU1B8LAtDktSmUzeEg
aA0xahDZnvn01iCzV6mqxdjJO5VFstM1MPJuhCLQ+jaA6B/5I7VK2cHWAwCd9hcs
7ElJ0sDZfR06vTRH5HwS+rdapPV2l5RJPcQpPoYfnNMj3JtC+HGHDnWZbDBEGKqT
TR6W7jBJqvhzmu25OXG+2l1XTfqt+pGh7NxnspiC53Uf5JaAhv/rUGnStsOygzVR
q7b+YLkYINj91egz4lrwvLLEyjeSrJH6RCy3k++UFsCIBMszB/hlx1wjEPItYUOy
tbEPytWURxaw7hZDil1P/qjLRgtoMiE6q7mgy7Jold0S1T/Yqgfty//NEC88fV8o
1jiSvRh8VPw5OzL3kN7JX6H/hknvC+0OGg8UgjUgfwoiGuvqjsceTwouiVKI216C
g+FDjr+3Zb+JljSHaU3Erc7ohGgJt4p9plFSJ5sP4m9YEe5tdp4lBsoF23Lijij3
jeVbMGEZLNEXCeverMIdBRzsvw5EjsubSLJ23OB9O7Z3O7FMwAabPSR+9hOAnOZx
xDnuFoqX3CaSLhLoLEymsKkHs5fr9y70rpxYUb25ZuMWQSFs8kRiiZcj9XyF+nIN
T08euWfIEn7zZCP7nc1l4ONm7YHT8s1u9TOYBW28FAe+/n1DwiVVIWKwAr7iOZZv
3ecbzlUrogkh/og7VTYON1HEdkuQc0tPz0uD/yQT7/6IIYi/WOCGwwMZr1beLxOS
6HlD/UMi0f5euoLwE8iuWrED72jSC+vqXt//yV06K1S+EZFWMn6HZs2Z+rpuaZz8
LJ+E7boJ5EEsZPoE97tpiR4UppJCNqomEGiqcKSGI+5Ku2GEwLIUM1wNkIv7l3KS
o6xnmcx+444oISDvOkFJXqUAdWByuwjElgOuvFC5AiWkRQMWOS0d2MsMHDt9jk8N
T7UDhr6Ff1Sj+5fWGJNHYynY5T/TFuMfxhlLt6TJXJfbwkFvLR2ljGBCyfmmrNKY
1P7WeBh8RovXHmtrxWc32mjn+Q3mAZnXqpLmUkDpHxag2u1o/3NC9fEE34zT4HtQ
LD8uyVn1U6LSW8FjHPKPKOjpi7giAb+Rvh3yppJ0IQOotak7N8UCFKCkd/2RP/kI
wDIae84pF3R2oFN2Uv88/2FisXR4kwzSdKU0YNbkGA8C9amXll9NY45X9A91xvI8
i5NyxsBA1X3imnstKeevzWsmkSdjAjr21xyAs0/Yg/Gd4dfsk91HiTk1e32w+Rcg
I7cCDETtcyZF7d8SYfo2nRxZyNnaxT2uVjsgZAJBPSrQswq02q4mWlDBwRFhYwgU
3xkmIYSo8McfrRqn83TvX/1q61rB+7SOoHLyimuzDwd7wbt+ERWizwrnV9bHzrek
mCHX+gnsLjmvrcngzNuGhBF4hM40qvAH5jy2eLT6AmEIDHukLbKYNy/rP+DczXLL
wfFT9eIE7EeXixKdKL5Lsw4RY2zU6kOSqXoE2mfrVQ6rKa/M1kVzGwV7GJB+Xcnl
w1VWcWW4HNw79cpGQmqMQLBoyjx4n6rEiCKHvreIzLWVLZAvuSM5lm2LPrzElU6T
WzC+R7mzt4pTwcQ1PNtISh8n5YgbAlpw4J4r9fPhphB/wlO5ln1Ez2E5g2YiUD7g
oQ6gI1jLWCMr8QeRuWCYY3AnFsIg69U0MFEW+iTm3XAS7Xqv3qJZADQt0zicn7VZ
6AKwJawP0LZ5DtkIyLRj4gE+yoPGyyYaCl5iBKkBs+rao12NtaqO7INew9B/6GX9
V8yTixg2bjywfWglL9D6c4+6YYCzn7pxpk3qlHTbyjIzWxg+d+bQ/eMGBTKpZe+T
zHQ7c8Wb1NWjCpfDNMd1yQ3HIB8y3N6ELuxq7s0OeQhn0TpesmQNlxnNBJRZ0AcD
JE471qo1FadA46e+5zKfh4b5WTTHsTx+akv93Cr0Z++ZHXJnLc39gUKUyKIEAAmi
JaslNxbDNijCb+CVzyNSK31kwY3n4mLvLYutvYfYjn7n3sLRHw6DKCI+BkwJfpDS
QSvawIfie3MR8RotE8yPgUPLBNKhyXJ3XyQORGq51Asom2ARoYXPziCnuCZTE3WW
vSamqTyNLozwJkedE/60Be+CKa/hdBP03kshWORzu08dUSHfdsN0vU4STWLlM/gF
yUZKlt2uXewHA3tFTgFlLw5Zic/2le3wJxndxeU/OWTC4755Jk0fSNj8TfGOSnG6
2p7mvAZ8KMzG9dgeqmg25hLZqI6PZ2xIm32LGL+JXVfarETZXufR8Gw/Ks5+/Jyg
rYc2UIUYyYCWYGldKGFEBJtNmkM9jbh3szO4MEokORCFzkN8wnQK+aqGEpWkBSDH
XWtgJzHDW4khbsP4m+fHyuc9NZRnS4pzrv3l6afNEu+BtbXNRpNfyqRUPDvcoTzD
qmdvOrWM9QdEB2QhgHE9dSQ3GOMR9+Ov7gkmRXE4RyuDvTAnp/Pq1bwAbwl2larD
dWGlG97YRhFZPlucdwkhtJwDYRvE3FjeajOz1mm/fu8r8Etb9XausV71KAOHGMtz
YnexGqS+eDrDBW4EiUn5wJt/nubtYQfGsaMHNgk7cf2cHCtarK3UEGfwjJh14uZf
b8BmnGizOh3eLgq/yNktN6TxjAAD4HZYPKdVKJYp5lYLAFkIfzsO8VypLjtQ+oBX
n6RC/Q9U3NnDkFh1AoVVUQQcewgIGPwYQncdC9ljICQsqPas/wry7TAfwdjt+T+o
yOIXlNVmi7wIHRdhVfsMOkrRTlKSGq/hoiKSZu9hRA04ZeG4c/mzG65xTBCILFtX
ZOnhUIFD5XI1veb/comaYGSj8aXHfgn6/2xeB+kcJTaicMDlE0UmJoEHuxtUlqSJ
jGgWNBbsG6uENKcKp+VgL6V1RuQ2wS+mQVCnsjQoWUBASVsztemsD5Qfau+OmNQk
U+hX1Hqf5TrJu4nklnGjOiqiuLDGOidx3NGAS79Mousx9bvRhCKVHuU8eEk9gZji
mDq8EGvcUnJ9V+8WXiFjLt4zkSO7yeqADKt7BOnWt1k3ARDptdufjxwEFdarPt5q
RULSQYgzLqLbj112YcsDThOBgMDc5valWIPiUqk9tlqTT6rL9XB5xkZ2frXYI+UT
AgI1nOeyPRj6tiXfMyYlfqW0QDuq8OUZl8aNi2MfiC/peSQFucVzbSOXMi0rflES
5f/gmJnHEIutVIXnulCT1SxXWkM5xtS6JL7tztuEwXg/XSzhfvbOXsNjCW8R74oT
E4Z3VAWZWbSENYtOlI+MzCNTqpvSo+H2YpqHRh9Ufc9C1sfnE4wjcX/NANo9PKrn
A9h6Ljndd2kiPz/9bUCbYSM+qASBp6K6BE4UNFxEtaLAVRo9jg/8zOJZmxX8LI5A
nREG1M1q+itYPOSGFi1tSrVYVfMoAmSSJIlAWwKXd5/jkJdsFwrlyEDiZ0sHbhdl
qrNsM4jkx70bgDP9+SvdXIZzt9eeTJcuWMrmRzYpNOlNrNlHqTpymXOksXUXJLWi
Ci23dD+ncdq4XcYtJpjiV3/HyqZnUBtpmAFSkXm7tSoGpBo4iIH5KtkP4/7Y8jKo
QvRzLfemsL+ONtxWV/Ubw+qogs1rs3YGFnPwR28T1DugK/5czOW2ZuexnToS+cB1
5Y2aLXMnBDQq0i7Nyn0eLOB2Y674bm4RxoyO6G4TjST10poxqO2VIy78A6ojc002
ofaLmNuE1xOwyrbz09nTX6iASRa8DWARqgtNuoBxG4PpWh9D1arCSH4ycZVHvdWb
5Cjp/mYccUiuOyLjA5wo1Al/eyhXqYauvK6/Fp7loWKhe0MVq6sAXDD68NZVgEDT
di6MPhJnjUS4+95Nzv+5HmfOnmbv4VdDvAfOmkjlrJdzoNcVlAj/ARCfYd5PqEf1
SDMh9AQbuINXiMgQhv4h0awN5Al0UymaHf7G89ZLekhllQX0uxd3hsfu029Oyuje
LPXCQ4N+IR2DpT7yIHKAGk4lA8hYL3LQWqoomdFLb9YEdhDnGFzp7gLjhU6LbJjD
Jy8zCdaIKcXuTFyAacNsa3hGdf/oPPvRDZLXQ7C8usf+a/xo6u1l2hgmrPgj9k+F
nNpwt53awCfDnSJFk23p6COvFcVvqJ31Ursoc3RdTwg3NGIj8qqMO3CjQbvhsH4Y
O7DCeGH6IkrVza4tJsngZxrIQyxzEg0R//syh+DqS77MEM6uJ7W+kYDT4EA61W5f
LXLYYtmoJjCzxBr9pSW1gnExd8pDK+wRx0DhZrBFERTDouXMpiXcc0JzcyfKf8B9
0RVC/oxzN3HlMZygBwWrwn9lSsqjOIjDSosLeUvfBzZGAQN3fKR1vB3uD0c+XJyt
bSoMvbCZPRHLyboerv1r+DxjHP6PD8bc9A+H3fwg+tC4Th5jF/Jopanc58Gd0guk
IcFXfa9Z6cDv/85xKlwtxuZwe91yFdcZ7SkbUUAwFjxb9fduPWEG0DbqSo/yfgEW
2LEkgW246Zs/gOripT26F0FV5JsaJAug7Z73U1zq0LSvhNDDpnxbqWZ/2O2E0v6v
lW0fDsDZskiJZ63NKsCWSFlzItg2/veTMYEEbP+r5K/5LuH52f4teFQiZAHRbEfe
wan3eBIAwXwxZBxQy4mczD0a/hpp/QyBsk1p/gJSqbtAjVE7ptszDoEOvASKnb86
1RezBgSEZD1JJvg5ovuxwg0JpP5F9plQcUDTaCDdy0tOQhfprmdMnMVdtycpo6Sd
y+dZPpRIJZDTDTpIXve7IMN9TBxN3hymgLy14ZoMUMfEUpD1OVEOkZRmYsWyWJ0I
ml8q9zbk9k7kt1pVcd+Gs+NsPlOTaHCtDmDwM1hAr1T0td9cdLKRKgPGvH0BOL6P
ksU8cIXbgk/5WlfNsRVftJlDBA9CbcinToEEx1zv9jNIpR22qq3XfMuJkw2Ev8wi
lhyQAxbj3sOnpGkoHRnRDFmDDZrVsZP8TTdjJeVjzEKww+kw2/UjvBcdYpLUCGUe
H3wVjSAsSctXwLU3bNF3mYsOFtbwN6A4EWddCVAWDr71kPOitkLTqynfLFM5fQ6J
c9N3BlvZ5E9VlCHEHFTEKkY4WfxFy6/Jyn7+1vBGGV+1LC3gu7JQhTfzpdrMXExU
rTcR4DLXyZ0ffee7m4KDxxHwPGXYikF0/qZwmWYHyOBkfY1YJfyh3kVJXQBcIKuc
ROpI9Kzuv4v8qHkeID+WY+2wWgNMT/WxYKg7gJL3+piiXAyyprr3mG6ntTtWHRbh
HBJDzFZKhREWME48ZldXaaeyxZOgeA97Xb0JkgRaYXr3NQMMcdb3t82am8JknNgn
xpCzWVRwg7yocdGPbjBX6mXfKSW2zyz0CCUDfYCqisEjn30QAQXpsE+wWIriycFr
PeZ6KTpHLBYUSNEg21lXcFd1nXfYPCs+sVfOR22BCVIWfP1I/Ettfsv+QZ8n0QBa
aJ9oQ9G6ZhPswFUZ4gVcniTLnvwHTe1rz26nNcMpgxPjTe0UrEXruMJ+Sv29icti
FfNzlidM2EIctxEcrsa9c882nT5kERe6PZFZxK3ICIRqSXb+UbaBzJ5YLlL5q9RJ
Mn7we2w78GmMWNHwHPiboviM3VytdlHsw2fMjNLLcZS7+wGdA1ITYwUhkzGPn04E
AgwESfGaaGvhhurwAmcOJIB6HsYvtwV4xN7v1A0p7bc952nglk3jMW/JTecQcqQG
62G8rhU7o1f5TmW3744YJMjVR7bHEmaPETUhwj8t/unAnWQJ0x2jpjpvYOsBCPs7
4g/sM0z28gLWE5o2fzhO5qtarjFheSjfHNYJAPLYf3GIw1xiH6s/pAg9qLO5F4S0
98FDT4yx4v/TJxlzzFZrwka9TRA6CMraE9W+2CDS/BkIQ6hDwuX23/M0gTW5ML/O
DkCch4wULpcTDfGt++ZKjY9lAX/C6+6bxPtgeTlT73G/3AB/n+15Fl2vZ6uQaiYN
qcxw96VQpDpiRiJS/g+73OMAHv/hCs6Aamv7udNqPqoS5h23leeGC/BxIAuqjETf
zHYGoB6uuBKN8olwsFA5xw8OBmA9oCmk2d6ZeGaYTwn7hTS/+e1zAopzm+BUjT13
j4SX2sCDGDkRMHm104mnedTfvGKdNAB4WoZl3gq7wvMZa1+p9QvPDbKlnRWhoica
w05Ea3i+iGhi6Y3gweWto2eXsX8jnFo7FjpGf1iBi++iJGWuxdgwkaPTYDMjs+K0
7g13AFBErL0ASzd5khpt7uZ8zNc7ejT5cuwMm6c3QDCX7UMCJjI7/NPotfOfaufx
tuy6BtUvlMV70tQYRQ3shcBQR75GzB8cyeS7OAY44hiVlDRvLZo5RNxGEBtexdWD
nPmiF73pXu9G5OvWDeY3ucgTIBm4otQNwUmfHPWXLWfgtlxJaGfSKccYYDmeiGjH
HfMcFHsm3T1PXSZM8EZQ/i32IWZ66Ye+C9aATPlzYZA8SvknxS6vMVy+yoC4/WpM
DaYLkTJfECXdS2MLRNuKhZiFSLLxLoO4x+U3vKDxChZoMiKpZP1Ukp2Fhgxirozk
DfkANUZLhhVD6XamB7maW8sdNAuSKRfk6Yg6PxQUI96xraJfkkRqtH4a3ufAgxRy
Y3LzQnpM4fdf+W8nn/zs/6dhw64ZGyYgzfJTIPwoIbRs5Pv8EknsCt+CL9xSNQuZ
2ISk0GRomNIpuefK8gQwLMTE+MvUdfUZUNFR830mumQrbNgE0O+M13HOya2x7Vq2
8oafsyCQkBiHLoIknEy9SKyMRH7X3HncD/2wtkNJ9MVNfuzx1cCwx6SKsSrpC6KS
Xhs+YQmeCUo6c3JCR7TmsgPwHlFLBevjo+oYPUrOO7xFO8YDC4ZW4lqahZQOMlkN
xBjht2IKrWSfWVTvsYEnR8SczSnqXEcoDsZqCYm9ZBFMTGBJi1igrHssX1agappF
geWi4zl/KEyMabn7pJoY0Mazzp4qwXrXx31z6phbJblpE2uLAArgskTKAU9Jh0Y+
/GCOZYzETRhg7IhIggJiAz2UniEMtT9l9MOfEUdbpF+dn7DDOkmNFBSAR9+w+bbi
R2nO0xlwI4E8pIbGVEHDAJdfRds1YdFrXuypJkPivmVgp3tz8g0D+lgbGC/veIC8
e4IpHBEXGaPfO6NFOi0skfYrQy9UgBf56T1fLiUA+DQkfyTLWYT2xewrDcw+v8Mw
pCNw+1UxrEF4RqfXMNTejXcZjzB1K4fTgI5UBo8dC8FX/XQ/EyUYkADPFXdPYQj2
biljdb4iQEWK7hHA+0w0AOwHbl8Rc87Um/vUSDKup6kNwtyG0gCKV7kiH9WBjY/8
AjNG10Mtt8vau6B0S4qU1/sk+XreVIKfmElrZLWmt9ugpFyG39wlO4xmgG+7rvnV
/bUjlzmfggC6xmqG3o8HExA6DWPuqG6b/Kexf5aYdrPIRyzqHyx8P8hVi6gTjGvb
KS+3mzS7VYMzvJbcKQmInsLZgImowtiQjt1rS2ZoGJYeKRzkEqNq7HuPUtfOWgFa
ToqDc6+q0gX3ifhLh3JfW9e2OF94dg2B7feQGmV2g4QGmvozACd29QMH+r1tCC6g
fZRzSc7Tm/NpM8Z7iNJwtkSrje6XtqChsr5YNyHbmMJ7Km6BrrHq1FjGX/dRgCg2
abfH8ILdCPh5nZaKeoFOkOn2TD3RAhKEffIjvedt5TjNlO3SEh4PD3zfn/WYhwSC
mNQYJrJusc5nhykJnI7/L7FxHtFauasv6xVOc2HMTa4rEluDy62fwEqVNc3z8CoV
npw6BjV00GbbOIH+Dnk4e6JvRdrF9Yy51z9WwRwwHY7+ULnAiynnUrIP96euKcbm
aDIOB3Kihp+fDqVsnPAr4q6ohLtvcBaSIRjF7+eBfoB99KPCmc2eShpOGYKjLMuu
jKHrGAsuG3GUc8uxr5HtNNkwg5VZBLLmXFagCFmjE2tOZ6Z9zdZUEAMSF+m8ta2v
fEHdK5+19AcQVB8sMHjqJmmyPCKNXqo/luu1CKayGCeJHzQ15bZnR09h8xqOS/F2
ztKwbyluIUE21kKtOTNsEBRkHLLabRshyDl4qQxlKQz6qC1ZZS37Iz5ob0RPuzCY
Xmih05uuOx5MV0NjzVcZE89MeOnnu/0uz9ZeSKvtTG3SD9ddEbWkNdl8pfkBTyAM
GeyQAHTCd3h8uZNwTW0/xO8yh6aPy0diiNqhwP1Rfkwbrsp9YXG0M/SNeWqJbeYf
FlKYmXB5ISL0PfHvpqfNZvY/0xD6un19v87XhFVwi1DC35vq3MAj5U0ZFSQ2SEXd
iN2SiurHzirB3ZATaXz6k/S/ORyu1Y1GgzdEl2ihqzsyfFX+YJkKA1scAVVXNnhR
T12H//erJIwALRR3YEUOTjdjaxhLIy6Jp17Y8hLBwPirwA330c8etcFCRjHT9mwM
6YZMSY9aaDqm1tqWIrUpcXYSFDGyP+e4HsNecy+NxBf76QTerQBplM69gO0lx15V
e7TTRVXN4pY9go0cDMkKYrFl6yt6tQAkZ2+B+ebtNVHu7Qtt715Kr2/RGNIzGHPa
+jl39hztPJ0c/WuGhhM1d4kXiW31pUr6kCXGK5b3jdiizJi4t7/U2+tE2ak5ZI30
OrnM+nXVoOFMioGBlEW7piyFv2k+ur4wazkeNmNLO1NWk6xLd6KR3/sHbcb1h/fI
wDGUDT4HR088Txo2CRvD5VhVCHC7oWHcGZozfeCHbSV1BaR5MbxgVUyXUYwSaWgE
YwWrJJaLpU6l6yQZch8lhfYls1xO8zl2J/UUvZ3IA8vqO9iyrutBuRsQF4TZ8gQL
0KNVWreDJb69XhFBPugCDSlslEO8aqDIKhtxtKn2sdXatBygv8J8LurQwzkbDNPd
roEfg3V6nMzanVXcuH4r5/LI/7ztNzRJt9WiiBMosSwNxg7QjwVspsfbNc3dn3ql
dfUJ8hXiyWLz8txJ25bu4IAVKzfR0uH20alL3Tpm/chrtPn77TUOh2HE00Cuvz/Z
3F/RdtlgrN39az5aJaJDtUuS2+uJp2at/AdtU+Wy5mFUduEtWUOrljtHUfLl9xaa
tSP0JtaftTGwEiG0GW6CJXdy7XsIugWFrp+uk41XZvK14LufrLMvFauw+H9VUZLe
G/QSMjBPYdMhYx5lotk37X6qpc+hRp6HMzHt2X4mHBG1cS/djHRCkSCbk6ihGWuL
2Ped7EdXrfQXX6xASwzHUOqu6v2d39n4v6EQfO/SNYFmInO5mAQivDereGeOF+K8
UXZgwkKEqsmFGUNYQNlQpo7MlmnRTUqGNB5xvr2TM2lNkTnkMk0TmGhQVkdzHQRQ
kVIFPVOxdcjuE/BwvET2LVv/48vHCL+AjbhdLhcni23474uGEMgjRjIcvinOqve5
UIg+SbAHrfCY+Bv/9D/B2ewgYdS3VroG/iDhQxdSmLmktfITlq5sykJEHxsXkS/p
bORMg+dffBgkOWNPK5TG9siiIC0c865TvcsZg9s25yJCthR34hD9A8OBfWZQ4s1k
p3bzL3K2zu+25Wrb67QcRBvjZeZbEZcE+Kn1f0jTNapMKHcZwGRZwgE+9622t73x
HJ/nENo9EkQGhDv6MILHSBjgMc5+bOutge+mWeRoTl3FyvIXKXdIjde5Xg9uD7oE
v8cokNfvgmTz6qLt4HQTOfcfMTyalgnY8N7zrxZckilaPJLMjVxA+Ba9EoO0+hYp
aNXeTPNoPYPf76o0yB2aq88R+PpggA/eY16srt0VQZSNhoyx3k1MULMFkaAx8O4c
lkYFS9g3Bbs3mlGwEReHcf4ktfoCK7BTKe0SToUdFQ/J9Hhbz7lOvxMFGa0fzlrc
a9feyRpNMRj64h0+o+l22NG7lu4h2Gl4sXZM8LRefVVWW6Kz7ngIRffmEW6WKjn6
saQjNrJXv8x/gZmQQXEk9FiCbUa8RH4tDnKWnb5/hfOAZ4PvRUpzAshQwaLjKfZH
yrAYozKR527fSK9IdGyGDK2XRCXeDbk+IdwLAFNQBDV1bmllk+UGnDZws89i82u0
prV0op5JOD4PU2a91hfRnclyn57COmb8xpoBopAUHhSOPxJIkDZ7eOYsvri7saOm
T0+JjjuU2800SOZlsTCJvCrGUXxg+/qZJ4sdI/r4Xe/IW+9md696lQjB95F9lFLi
Kq/RRXg7CsiP+iZorFHemvnveqvR0J2rc94CTDltlphfF2mWKEq0AOfiH4bOc7Yh
Eyi65yr70L+vYksE4tlMEjiDTQlsV4mW2k4gZltr0nJK9r9UXg9PErhxNNVmRj0s
fuBa6YiUsC9lqV4Ax/REpZ3zGBuJLTXMI29WkqQJgz9CRYt72oGf/Gd5myQvUI77
yV6Sy7sHcJw9aQoPCx8BaN34LBZnk2E0KJl3cO5zY1dPB2Dd3qMPjAwGLr5rT1Oe
Siroe+pF4P/2sj/qZJIxVqdUH+bdkQZrvzqxeUknN8b80khuYTzPN4xW11wqC0c7
dlyUFzhp15S7zQjBRqJArV+KoPyOag/Wn/Aiw6YtNUh2+S+T2PFViErgTyJcPYyG
1lPQFbbhu/vh7OQ2ACzILWHcbgyVFHmm1sJZ6WWv0W2InoxPqN1X5WqILIMNVnPU
06yk8IBVpk74j6M4E6U6FT1QoTjSfqG23kX3p6lsVLSmDMil3kQoRY6fOdNqf6Rx
nQMczDDYxbUeG5J4LN7GHOJcte1C25pxVnS+hl9MIQHyIhS7CbZWU/NJjiYuI0Jn
qIhfa/t/6wuQrdXpZ09TA2bIEjoGATDFOrCsEmxDyY19eQXOu+JAX0eUN0W/BF2+
IBJiMD/dv3jX1eo044wXZWMGtYQcy+n9PfjYWO+Cbqt4rb2ZNrPwV//nUEPS1pMt
nko+dhZTfEFIsoDhx4O1zrnQu/6wvFml8ve9EpvzL3fbKhRqZ+koYYNa8pTkLlo7
yMBNdwLQq9OBeX3w8tTG1ODzkXZD4hwU8LGtvEMEkn2DsEQlizBsFDoUx9OJwT92
ockgMMkuvG/dx5w1zh53/66BNlry6bzo2tlGAhz9r8fPElsYVzH1BwsezXyxQr9u
VTkzlNtg94+eUOaZPBtB646j1xG/Dojf/1tDT1Uf+UvuhZPFFPltdS63O+Fma47v
Q93mllnFlbxFkmvkHRJ8ND+RSlqUnolce3mRgpelnzn1yIi+pqCgzkAYmoaOhfmg
OjzLaMMzYQz/JSMCEV8zk7RD3XH/niHAb3VmxgK05oXFPEdZHpwvX4E55fkbKFli
lYUVns0N6qL5z9jz9rmqhvrNUaunyaRNCDAN2pdECcQknZRkvxNAQ79nWrXz9zZz
16/t1ViXpfWmmTq4a8e5mlKqvnlguhNa9QsBIqtN+sHVjKoAamqtlUdELmK5o/ur
6suOvy2fKyMA4LvjYYW8kxR8TMulpgInFNRkSKtuvQqH26ePr52nquYMmMN9YAQ2
PTeYOESK0/IGqDhgxjbsGVqkimXF1e55EFaxVYV/JolVzB1KvrhciCy46xBXROWR
FFNgQZ92TnKKJeeGGK/W8rsfnQu/1KxAnJDW7zphakISmjrbQyW3Ngiqg+40+Ism
w6CjQiHKAknVJJ1ZBLdxlCEpKQPwtxf5EOs/Gm/eYt3WkoXXTGt1z461Xz/KOGCc
1Imx7klPJzUP7sqxH1wOY0sNKz2CARaO/bLNwJfpq5mdG8VKTkif2TXc7NUHtsPu
a6R17Wl9ffK8sd7eoVpgApeuEgFJ/VeQJDw6ag/c17zDF8DF7YWu5clqCGbe+fGN
v+vMMiiix4IZbavedF/C+Cv0Hd47/seC/jw5UXTRyzDCccyatO5s4INTrtoSwjMu
MD9Kuwis+preOZcMxpVeW+PHvRZrKC9KTpta+p8fpDB+IF5ejYOZxKt5fKfyookn
fwKrQuM7Y9DnABgsbYeJstrIv96JaEQNpW9so8kepfKUM2KQNHxZ/iYCpe1AwEFz
sJXcySa2hxNA506pK5EgJ0LR7fVAO4HaMnP8veTp0lhNNEK9TEq2Fwz/hFjCUYL8
H9p0OAvCKoozdH6E/cTYdnF/DKqhP6jxbsUzaIAbUMzpJgy9mIdH5liMVHA/MqI+
euDm5mqehCe18ED8/JCICZ2ny/lowM6nyvEGCFv7jMtmYAglN/Yp8VKBM5+9crDt
ammxxGCNF0rcZjw5KMJloRjMONi1kfm6A/EkuM1inbV1SCGTNPlOAySYEtwHVlHy
t63LA+kSYuxQf7vEROC2FAqlcwL2ePg5zXrYfGz2F2667hNyIN8EteAX5n/VT/9P
84WLqEnoGvvUU7VCwg4uANowGnFaDkSjY1e41KNiJrJ7xdCFc3QzqmwJNHI9yHKC
Fh4F4llTTwoda28qftgtA9dG9dAGqLDgnOeHrmHvOK5Z1yUD7N/J0s24GRUVaFuv
SqdZd+HHnd6MvIm/A1SaDxyTELbvUTfDKJXiAK6czX/z9347RlA9xhSQB7UJKhCA
w9mcz8lP3dIDCFuXhhV6XlsADo7kzn9RglN9rx82kOeZtd6rnNUBMnZiYtln9dp7
XsIonWOtx0q4xKvVNF+oJvc5Hp6A/9tfSIAU0qe32xts+DH2OGesKNRy4sSXENlD
hDwSTpF2nugZE4XlDGccOuXQvg+a9NCMS0ckKTCRkNDNwrwZwnHCVDLiQ2D566P5
F0ODaDVMwQ36mpzKrnoT5etrxa8XHN4wLkSrhbhNW6xdIUp8TKJRlyS2DMEr5XiV
lIKa0t8ReBvuomgHKlii6dGyN0BUlU4TPKmvIsU/dviPjAaXytQ4d9Gn7GquRSyT
cfwrfxV7aXEsCOUeZcRv7T8ipiccCxJol1LHPw34FGWeB7fWSE+5I9ScG8/C+X3a
C2i+avReSggE+N6QCZMzw5g+hPOwWOJ/GaYQlc7bzF5FPJCx42Z1gteLv3wlgZPc
73Dpm9F0x79mv2kwFzlfWm/Kq0jKWJLEj6Kmu58LPAMwetXU30N5yTkh1uRJOEtK
PB4sUos5B/tD9/1xnaDtTA5PRKfzG0GSK7C5QoZIjFa3LJs+eYz1xGaVaj0nbaWO
A4ro+J5j1wvzMTlC0VwSpFPIx08xOQvGeKCXazxVVQJse7FQfuwqmToJ6RkeV0Wb
zktPz7UQ3ryWfJBBBPHEHqZhIQWB8kO/9mivhDUP9vcjboMSdhsCEsmoEVN3+sAM
a/wbVhNDes06m5hBHVOfR7Ukq1m18vuZhIMC66RCcSr1aAGNScVZJefzlsuHzRc4
2RHSGajlmgi2eM7EXpHWdTc0lDZ6vNsqySeJnytt2rNc4zk18GCUa/3wdU8o+9It
A7YOWWo1rVjuZZpSjzLrAjy8YHCXi8x0RlMFjoz72UeX7JwbBkn732BvNEmDjO3Q
uKxyfn0l3iZlv8xAzLXa1KVmMcnimkqKFxZbQgs+c9SX6YowygFtK4zb68pd/4q0
/qB4FeeQd9/DY1vNy6W0zfSk4CBxtbPe91rzZ2y04E+pPuoueLZSLBg53qa+WY/L
PsJhXgPu+GgHsJmjPVUGQZRRV0o5tJylSVquyZaglEedygWYSWQvrC2kM4JnaqbT
cYPezOHxEoThgb6fN2etyoCz7T8OVYyTJyFIcd90l/p8/N+L5wL/h3veZURbE8Eq
mdFMFA7/kO7Ubju1GVPosQzamgdwEHnEXSqpbyUOYpvvald93Y7NnXd1rOjaWR6F
YphtgK3uU4OkNIFZfFlw4TW+KQzziUzl95FKeJx9yIciCMepa/DReOn2IOe4Nc5+
6AA1WLSK6CEw8+liYxFHoQpdmfNa0EIUqC0DgoJVk/NEwx6434fKKIbMfEvwH92k
+7fT1SVO2vuOUNYCVEle5XNiLD+6oEMhGJ4XbexecaVDlxIpt2UCW6FzdzEDYOpX
vkPh58hXM5KcqgFOWavgyteIrb6MT1ciDOHagkFsi3cqVhLOjunMZVLzbMJLvvUX
7NJdQpwgiNUxhz//J5EC9MiwDjs1ApPS2atxLFBKJ/LFeWpufoHX9Fw/EM8i161Y
STABCfG34DM38sdV1rirem3uuP3dtqWMtmA9/L76Wp2AaHKwMNu9/mFtRw3klnuP
IKGn11geTazxFGJ+o1sPXSp8NHx+uhTNrZoOkwZ7SLPbflXCB9BmjLLufVgXvJW2
fbCSl5ahXJGE0a3cRv9PP98pSE7PnJ1YS+lnPTZx0RI3xbKavDuyoqyB+QLkLaiY
Jl+bGsDVVMklhtOz9whuUGA5eDZMS9MUjbGNCSx9ci48ZWSCw7Htrh2nBeYN/o6J
/5KLDBMsrfFj/VmWRU4gdbRAF0sMGXPunlYNz3Dek4jc59G+FARQVgfFS4liBBDc
mmIclOESETMF2JO15wiDFM9+2xVM1cd2S2l75U++bqC8PA9LOhgn+wwRkX2poPEP
XnI0WRqZUMuuEDTH6g1g/OKM+0NhwRnpBte+pqIk1gVaBv4o+uOHNSpULik9yjaB
yd7JseWL0YyrUDpjlfHhLAhG9BgKlEGPIXYlniWjc/fM0R761p4G45YOHuv5xsXk
FAPdPd/pjAf/GuBLwXqiblkQnkHRk9C3JzIWxp8QA1YjWBJyxepQCJKh9DeXszNA
x1UqSA+PFbJYZ6zdSCNeqBVLIZ70ejciMS2P/f7TvPwze1HoiJRKjZcJvQPILwrB
yUtV8bk9C2/DZPKTpUq82OBfOf3wWml2vG6dylSEpDv6/EAt+zHldxaP2TS+wXRj
lbBD63lGzEnNVXah7iSxxa2Nxx3z0xhbGknwTtq3+IX68fkAKLaO3FZIzVTtKGL+
XThO8JExgY+F5EMPZ4nXrReVr4nua7TQQ834dKR7YGmRaIDOI4dlLvsBvWdGH2AQ
M16lWdATisy+6EH09Hd3OXqJNyEIsvvpg5T7iOgkH6Eg1qeYEN/bgHuhZb8tqGIS
V2RMB9wMokG9Bz/+DI06GvNhwCc96LR0QzZq0QRQTWWV98WrzrPv9P6RWeX72UjL
lF7h6ptqKO2kKUdWqWrROl0Rpn/odl9TV8BJbeti+75J3lOBNKzH0sp0ov+yniKj
fBoSOHQgfsPrXyE5ZUpmE+mKQvdMX3NPVpLVkz+zdwHGjvY9A0QihGZAomxOK0Dk
nZ9F2NYVizNsK8oriHLjjcXDoNgpZjLOSQSXP/4orE+3arCgRTTPHpaVgN4WwZ62
2tiXvW9zAd5zivtOVqP1SGbf3RKYJFe4UnIg1hD2JYLRoDyZtalVi0ThMa/Yp+67
nTN1zG74onevVk0O3cRcIXHMLPms/8XeFpiZbceMpFlPs775f8r4xS2cUuYljJZI
zvyhNLTMxpIhYNYUabPdEOYVXtuPLY4tZatrRoV80pJNaBoZc0+VjPLVUg1+jFVv
iM4z5qcLlI0ULE1ZrE1ncpLDD955w81+EsK9+iSmE578roQ/gYd9KGB+KotBJRsv
1DEiCjJ4CXiZTgU80hUNQLVbHe2G76uOahsZ+J43QfWoz3883lxKp8f0YUnFffQk
7Rry0X9j7gksoEeq6xTIrjTdHvXVywnBQ+Fu3OWk83xHefplkHEAVT4KvWKxH4cI
Bi3m6zP/ujuE1PMZzH4JxM4mBBhhQjCGuuzjWkjC8W+PGSbQFb5YAwdBCrv7ptam
lfs1Lj5ZRxq7BkxE38WMpD+jnxUBJh5xpaFXXulDvjWaH+aqa4AzJ0qpVvvI4yfW
ekmyK3wbhSIIKtQWLVIduVAyxvLMqYNyEgBn6kK9UlwkMI3baNN5eC1Fx/IjhoKW
AGyFLqASQ0lkIr6iLMjsmXyrdSIV3ZzcusFlHqva8UuaJkYrqELzWRRJzmiZj3BJ
JpjA0qGsbjB+qiJ3KBPf14cRxxEaCd1zt2WYKy2wkq2A+XqIWQ4fkoAcX0CUAjQ0
Oy2Y8iwZhMdib+NVx93xj2Go7UfEXObSQ00rY0/6wd268Irevbsq5DSjQBU0qbN3
6Xj94GAK5eCmQX3YimChdqbWxaIRNqi3epENU9ZG50AeKb0YywTlV4TUvJDj6ZKE
dsvAartGbvhdw6UYPOzJtKt8PaaHv+B8X6BVeJPez99Ub0LMN61T5HJ6AuYR/STh
YTO3CKSIWTJU4/mM8xP3Qwqi+aqJIp9l86GRzgjMtQIolX56iNUYE/g5HWKXoj/j
fXAJxQYqDNfJjYIaIdLJvCa4H57xSiAccq5IBpCQVv2E3fayR92ZoXnVFpI3T4an
cu/Ov0zLJARUptF6w8pRvZZkALWFkgovgIwRhf4FvjMXXAR5GejKeL+59outfZn+
xKIdD2cV6vJPVOKOA6+dOQEQZJjeEeTHOUMih84CxLoFvSbDVGSKF1107iIip3BT
vzucdafMQHDW4MEnsNjVgBxC43BsYPhg8zndliG7ZUlEqFXkNwZkoLOwiHMOwHjM
EAQv1LLB45Sy8B82qCb1QtpUoID+PQZ3a/EEKU6YLnJbdJsWWc/VEU18SKrMYjlW
dqt63KY5SyStIzwTY9L5Fx6TsiSuY5lRMLPHqsViJfE7r20mKmDjXZQLfaW7RrtW
QV65SWbB0ghzz6SZjxqKJ7hEmBhnE3ikfk0CsduOVNRoctZuZeO867lHX7cptoA7
euRZRmDoSv4REXMRYh4R5Xfdv/YnzRnFXy0PEfpLw2/RDrww2cPrv0/ICfA1ZtLp
nla7r6C8a39sIHoIkJiWYbQl1PlSRYhIYfjGwSnW0vtvBzdjwgDv15HLxHpxg4Ad
Cr+C8/Ca9Nybs+tVv3OXcB1ShAtBREVvUgWn5/HFHqMc+HgXeCNK72gLGeya2QWC
CAbFUM14J1FQld0ruB0wpWBEl8aZ4TqplSbccjTBtBn8WxgPegkoLcQQaVoASFHd
YfCvDByGPjAnsYukixQqkRAUxdkqVXJX53EvJOnaFnLcfAWfqs4sAX1z2/y9l8CD
skHdGpN9BdfrrNG0SojmB97NIg1tIbJXgybEikfp2G9sS+d299/cboHuMaAQYmB3
F+kRaaqusmBmGuJpYlB/JTHBCxycSa1Qlv15Ygst8UC68+S7Y3cXRSL25mTmuntK
E+Xx+ZjejbuRe/dUp3l27tT2ReLXull1USmUme1ixYAgMsyD+S26wIPzFjflNP5g
LwXIqGY4Ie8XzjEohk5xJODGQbzEKSyGzXevjNV273llhMIVBBd3RGXIpwJiRi+o
WvSV/1r2uz4Fc72IFCUoHxITTwUkjv+71m46h+uVUDLJ7jis+0WdS/1ah2Zg79Jd
XTtJ4GPUoE+pi3gHUVWkNirJif/LNtUqNBC0lLOWdxVyi8IREHdnWmpmeAlbhfXr
PynmOR/95k+ZZfx84aW2QpLvtGKrm8fvhilU3m4rWKowKFUEZ82f0tDDF3Vj8CgS
QIu7HTYxrCJD6Mxw6JUI4s/cfKS7xW58qeXfUNZySA1lpzGYemYpVZXRLuBKQFkF
7oJhwQB9fg8YirIb+BL0ZzIDliOqVAmJzDowpSPz0o2vQMnv5eMhs0nwZapzyfX0
tG3QM03Vi7EYp2Vj1ZFo48McOiVd7gPsvkhdyWC4DPFl8hV/+ezNgB49L8zzeXZ2
WO/0MDdsk+8YjGa3GQupr85SgxbC7ekU1Arzy96TCG/vkAauayzqTg/88Yc87YYo
0I1fMjkIFyyY2+z+tANSE69J+zZLb0FWIRQxeKJaxxi95UwhxUEyYego8mgD6zcE
e7LeFiEMmWFQj3e1uUpiJZHzr305t+9JmFwGL2Gl20PwC+iomIQiRUIKP+mb981T
nVjkUGTJ5rtRn8gocHTGMO/60RFCoIYmZdx7QurXR5EXNNH+vSETpxQvokvkHjex
Dp1PDUNk2ojyeWITIchZp6ShdLmUDF6xH5NL5InKu9DdzlkdV/mcch/+mhQa65oI
x8KjQueumLEAgM1N3GjwqJR6dhDRaL7Z6ZrBir98Oi2vL6qOapikrliNC0F1/8Cq
J23Qkj5fU+ZxsibAawZGofK+qjL3497UdsnKAVunSXcKiqwTLDMSKr63G4hOERXd
ZWlWhmIoeITWzqlDHGFGjd8tuTS09UtcJRrjFzBRPa473YYhiYuWq1XTsrmsBFc+
5YkryZFYWPH46IOlfRRs/j+xMuBHGVPA6FcaEMizCNyxztLuEx70Lm16XTLD3LuD
bUXAjM/Vye52lYN6W0s4lkbBaLECdF5+UUX9yKrqA4aj8yUJyua3iXLd47T5wROI
g0Xlx9jL0OAAPTM3FRvrwsgcYiH99TVq74N8jyD53MRz6gFllSl917yQ+KWXMBqR
828+8bewSK9kpXqYpM4/9mPKv3VeVokAwO3nr60qyNqLEb/CguwVOLZ5bnVHYSoJ
2Apv9m5ijjCSIN6icynJiUXVjcbYJktb7tFDJjG5pguARfjLstWxJVLMBh0Jwi1y
lkf4xWWI8JFXth3g72xJ0CyrRQchygiJlQFHmPWZegsDYyoERnPMx7BxuTG/ns7w
wQ6Z976DC9SEBGmWXX3NDd9uNxiQmlsLXuTgzGiNGEcEZvLSDw2s4n4igXthl52y
tSFxTVdG8OipbS8wJBzBDp93y/icHkgAjkkY4hIkLj2TtnvlUGGuCCnYGVSB2hRO
hzUidraaWFptKfZzOyPds1c+/r6nXgnPmZnbRnraPnMMnxzUDsIBReKyK6KDGx8J
YGadEeg2ppcQswC/roC/SBr8eA1zzXS9Zsqh7xaDdD2u4ii5svL/+ZsE7VuEmFE+
s8opOd0dydTSBqthHwO1k+v6FRs/fPp64+lDXzblKLmnAnTcufa+99DB57KFf9HO
2nExpqMWiYmB5cMJALlDOXa376aZ5JFXxW9IvPvfL5NRvbaRZJJbKZwBg9wXS8xk
UYqTkvB0XJo8qZcGcOjhCwbB/ToTdvjTDyF/zpa1qfItPuHrw5X6EcY8g8fEfjGh
fli0MpQz0FtawLH9yP7txFVbRjfZGb1lSAxqClobAB3w891anm2cPUe5wuVzfxkd
/hxl1iNkcWwCnS93pRF2xXlwPZxOzNL+eLpliu5ydG6G35Qs5dlnOrrLqWdD6+Lp
q4UvIY73WKtlfmPtaBCdDpQbV5QB5juaG0dCfrEKvoWS9FCLj0abacjz63nDEXCP
nLull9wLTw0U9rHxW4cUBTTeU+xtmbE3g7cavmcSAF07FDfEdAPGytz8jLvKUxNS
z2ZEKvr3BdtURiEtyYXG68XPzkDEUkTDHbgTq71bp77ZyLAEWeHdwb4usaJJxuWT
pufhRp/0qsxhrhIHETnctJXxqIQp4NKL2YvVvKiQSOciOIWNGt9sSCMU/pO99lKF
Ers5jJB4IrX3/menKUi5+gxCOGZwK53b3i5Yf96ZldHnRwH7jJ2MbF1i+4z6KT0o
9I0gaOuyrSeMC8QNpmF1VYxHx4AHipixuK0AdV2sytnx/bw1IBuhg/zF+aIFawTG
v4OJx78Fma5A2yZ2qqPcuoRsppKQsZJSEKD9sGAjpAIYj5QIO6ksrao1jffcHI//
kS694YYpbFZGT8Z5J8wuyyXphWLW0VEg6yvJvrV8wVjzfUJEl7oiQHIX3fyhylSL
cuVEiFIdwSs5yxPRmOnEH3J8vGWdiVHLVEom/jNvwkwaef4WBnul/7IElkes9hbe
0gCPAFJIHFFgN7Hx8b4QLamPNWOZswAmIQujYI8lUg4464itJ82+CuW0TK3qaAys
6f4KxupHMuxx+b4SiGCs/Sgt6m4iDFKAD2XN3YZ/0QZ8J+e66tYDHqWYqO1vd+2E
4Aa1cjBOIdkwCXc81X4RjIjgjVLPBRDEV2YnLrwNSX31Dh/QchFcwEl5aPniawn+
NsJ1LAmx5rSZxVnZq/+6eaAKziSDvb1tSuodm0/05Jpt6YWiLnQwCXcYFzIDPbGP
eEY553uW265hDoj+ApX4Y8OW4BAqLUhraY0HMUuTkWXNFCy91JRmKpPx/lPmH3/p
JAiiIeMHiy4p17MsVqgt8gE5JJUgLBIRgGuh/flkDu5WJKtUpX4u6hAKgJyECsbt
5FpxwV6Cy6YwrJqHM2JDhxhaQcyTzU40r3vg2m5WbFnZmULdZ47AneerCmkxJRNH
leSig7RC+SxffipodtcVqsolr2j2nmuMD4Qnub8KDWcx5FDJz46+8wIaKsqXhxh1
VqJ72lvm45D8klKTPjT2mhoRszZr+NnDv9nxHFWu+HKmqZhd5CJh+t+VNXKpt2eJ
Qj7SkLn4jvzozBf/ceNOz3cA9AaOtFwO55dE5sh9PvZd0B9jHCjdxc5AKCp8H9Ca
5Z0TWNc219O3tm6A0XtxC4hPm4FRbcjDP915BH3gBBnpMywRJg1PycLLdCbCr201
fuULHi50W5Yfeqp1WKjgGr1ob2OuyH+UkC+YcujTReSXKp9ifbI/GuAzZx+UBf9m
sQy8DVjiUynYzmIscLjNJH1Q9wwNZVeOcHGRTRI0rPECqxmHWUxNszp7f8Gly/I0
zoXZfvTPB4yE/bQnfmugb4xvkc12gWb+WAFRXup0XkdojVaT+SVM3GM9rL7BvHwr
Jjk7uYEbVN6GAQH72lO8R99oFpWef7kLbq2Msj0Q4RhcOU6QXqsuzJWujcK/zSs9
vhicwB3bSOqwO8kfR16SFFAQQj307zlw+scQrBKv0umOiLtebSdaeOoAw4iWRlEJ
cLGX9UQ2a9g+ggPbwDcXzCWquU+ieycdqfPxtJjUTtg5A/5ozyIfcVjZCkaZ1/bk
2073NuAy8fdujiH1Rd5NyFF7L/izrQy1nT53vHathYdjZtrrJxIo0+aYyjMPfN6n
UB4SXAV7y9zdD9pw2pwuc8okRe7dUPjRcEt86XctEEXeuYUgzLKZTh28vRge4+el
xGDbUk5cHGce5dZP4BmclWHOa9JhwsgS0RS5zvUiizb2kHYydi+EXoRjTxz6rKX1
WM12wuvk2Xw4MSnzJfB7TkcssXCpPmArHCa9SZIgpvPOtScidBAHCHZy2SwllfYS
X7GQBst/o9p969Lewn8ZgHEJ6Hw1omkaM+uT0vH0zyU/KcT4wIaVBePVal9xxWP9
+OMdjYtSvCzpayf+IbC2HCPJs9bvzzCzWxzmnZkESNfiUsbno7T7aA89X26FJSze
WaoCOD6j6kzWndjcRisslo6UCywdxjeqziiWzcNtJqyL2DZOGyvwhDqS+gWFUXdG
q9FkxEJOExIECYcjRC1bRPEXNEcFTwScRMxV1207YRcolizCJoiAT1F3ddxwIU4S
GGnuDQqu9wacY1h+zMugnAcEj8u27fBB5dR2FxvWNPuYrfpUYwJtYaGuFVSZ2aq8
5zoAd5cFCkLUizPqFwM6QSNDChLt+RH445K7Lp+pwN1pkPVKYm8nHKvw+SQKSfpJ
qC2ToShrrRMMesjb7/sS+Ihvx+/80JqJvx5OuPlNG38GWYdRPV6p6qW/iKwj7u3b
0EJzdXO7jbX2vaBcltUDuxxeJ5pzWnLLQwcjjqW1AccX5KQj4HOyyHV25n4p+Nj3
0itUAolMs3IKMNYKfdQAdKFnKfco9OHR9JTSSX8XX2H3HO5+P8hL1ZRnOZJoItTk
+Ddv5r6uroVkkKST1MfudY3aWIpVcZmVdSHUmeCZ+6rxy93M8+Dc/VP4kcTCFGmf
IGL9VY3H4g8DbTIWC9negmc96rd3/6PT9uRP+bEjzBt7qJY9x/sN9KlIcn0od1hm
zFoM4bWBzHpJHu8JRTqD1++vje4rnV18EfumF37nxg7QjvnKS1LVTdMBE8lQJye9
WkcGra9uqcNTMSCaATyPyxlL8dcCPhu84I3T7HVFSfSo8QhUKYm2xAAhBPWkRVCl
urJee5+TGx70jKpsTNrD08OIYvji/NmKAqtad7fvOxwLeoDpYA8awFiVCkfdsPf2
a2IFUWsR5xRFNreUOjyPTKSiyKAxylCPVjYUOhpox7RHYJor/GLf9SvXGmhcQp2B
624ZVeQhcaLvWrVQKNrp5+IrD9WNsUftme0TfSMX5ATjulzxh5q/uakrijis/dw7
cprEDxalgoeI8HQSQEGx6dJKt1CKa/XaqtEJocd1g0SFUMvozt/DWwnLFd8t5aza
1I9BQeWYZCsVtyRmL4WRV0RDW2Yv5sm+q4xkhqGwVOGni/KlU7y5IkwEY+Q5NQD3
Bw3wIR2XK1WAQKWME76dv092h64YhgNhXDP6c+tUUTjOxWuJJZNfdsL448XqkQjY
yB3Ak0R3TAvAoRn7gHWSYUzyetzcRJjs7hhksCyfCdqdOdfeosyCRRyaEcN6XaTx
0izUAj3kK0d69rgKHRnsuiZ5q5ss9yBuXby1e4P+PxmK2jHyepFrVoLkRnwxmOCN
sCgtK5Rz3snwtViui5VWR9cRuXc5T22xyWVxpRcWpIwehbK9uT8UsdW1Ql83AXVu
zCNivwVdcYNZ73BmB+s2v5VmxyzMCiQM+6irXXTYwD4dX6Nx4+zqJ+7I/Cm5NcQg
PcuSDIfAvdquKcbzKMInrXly4YywqUU0SR1BGIaQgQfN51f6IakoK3ssrl+Da85z
sjdf5B9OFK3MrJvMNUfGgX7IAJbQDlNSmQ/2vRAbMG+Bsq1j7iBnEmWV5UeMandd
5wZv5Pn2DQyaDsb6j5YU/WgtjXiF85eCaPGdeDVxjGP8CwsApnJen+U+MX+V+iBS
7AfLN8v9dxjZcPQ1HWqhxwgDyzVlz7kS31J5PVG/h7OsIk4ueEny/yxUldmP+I2C
+wKe02u4YK7wDT9XWR1LoOSwB+GgAsBhsPKT5ZeV+vmQ4qp4/+ZwKKv7Z3znR4fe
gW8FgPF7oHmULXWOQQNsioHZtvj2ck/NxlZVz+80irWosRNAWzes9t3UcHCQ9BS3
q7XN0h3RbAEhWgo1BjolBfv27eksNRk6axuoqUIrFEcaDDUBfQhNYgKUajnOExqQ
Z/A9gPlbrhZApcTQ9Frr8x7XzC++r6L0cUvJj1b5WgCmHr+16vc/yZ8QKWF3w8zd
CRkYSN+JCme7H8qqplNOMpJouSQ8LbVlWDpKKq+YK88RmvqdJ+iUAhIlkimsNxcM
s/wMZUWWJ/mlZNoGViazziPTPXPPRkxzff6jIfJlhB56q70p3P0KiM3+vpWoZYeR
lsFOgPwUPN1akFgp0eJqCYkvVPEp1iugEVGKxlBiQ/POaS+h4ktBkcCiYJCc974+
/LfRU82ddZihhUAAx+RE4Mz57TDt1sT/2vQjgCVTSr27OTni70LX5r21SBGuYNpv
byY18qgqExFmjsb4znbGmZJNRa93jrgRQi/1UylR8uJ7XAKfd9NXrX4PlzVRRSSU
lXo7cPMN1nPLCdJ5zdYZ5A47w0YQCGcX4LNQ9fyIyiwrWlgZxG4RyxKdEaOSCwmq
cqLY/TUd/Pe3VqXQJsIA3r0FkiJCqqJSOEkjwb4y7c06SEx2Okz27Q384GTNRmwk
Fxm4sCRDRkGabowHi673ryKxtp/BsjBjORcrFYqmn2zPGb9TQEphTWbztOi3JtrT
dVdcVQroeEVvZBqXlMGsKbJRDwsEAcADfI1Yeqf8mP5vp9mWGJUK/fTfWeY3XiHK
d3flSw/CLUFrMqAmVvN9RoZoN5YE8QDUV3yE6UpblvRmE+o0WVPmydfO27Oahacu
Dgt5SxSJPmgU5pKgnm+SC22sYhdaEmfrTbf1ZoXYc2GfkenAvn+Ygky3c/ET5mCl
rHXbBTZNwt6r1LzlirIkaQWcMUMCafls6KktZkl9cZD77RyD00LAR0dBSKJRiHSb
blgwgPL1AtbkpxcpgM8aLywORJsIyy/Dop8bgBI6k+nWOs3DWXheSKNPE+r9os0C
rPmAaI0ENVnmlJVNnzIQuoxcQ5Do5N0K+VQfmZuZmnkRq/FeiXfhjg0AcmmJUGPO
zn9M8/WePv+CE+lc3nrprMXkVPY2TlQmGnfl1VyRxyUhoo0U3jr5BnRKzS+q5ny/
448uS9Kokr+MbwZ3RAL1BY70DRB3ow+VNWVcbWmx7mIrJZVCZ0bIejR4QgbV/384
jhVNlD9SwzFDM5A/7wNVw45ZpBLKkrjHidUf9m72gGjTQOb1UvJsq0rsNM0DwD7x
TFyvTXCpzxwm+XjvSRxxJElB1yKeF1AtU4wLTmtm+Ty5kThZDD18HTbyRgDdn9rm
RByQRDkhZrNu21/jII2PmSarkf3mZwiyNkyV/wdpIQeZ4zTG8vQg01dhiBpqH12Q
d7GkzVC0QvjKGorpwKpj+ldkBJuT6UYqcvCr5eXjlDr9V+x3WViKWVCLc5ZJtHUs
Ad9cLOV9WCS5tHrGW+pIca8rYeZ3cpHLaTblIGBqIdmABl6xFsTsyx6LcJQNq5PL
p4a2V5e/igG6bXzzFHe/ldoI59rhwdBInD0IRjd4eRfUVGBntokUUzTY6bbRwG7i
OpAg4YY2yLhmGVXB0JrIvd6gQbrfNnLpWs3iseCGTmsOUqq3IvOdwex6zgPmitmX
mpAW6bdi9mzG3/2KHFrfF9iWXqI6/PFhhDFPNLErxFm8hVkDzy9QfV1h42Fywdzj
A5Rlps8AHaTh/fiIg2t3aFzIvf0lnp2gT3KQ7O6CghnXzolgCcqI8JWA5Gm+xoCK
6wsvCaVCS2n5o1HKzrZV86vxqjeJabq5C+OQIp3/WTCC6USqIKenFXwnodZU6Dou
52smFv+JkiZM7ssxZ4vo+7yZyDUBEux98G2WMbWPjgHk+wro3VEKZrg1oSW253bC
n69jPvsFB7Lgv07tqNYrHu7NcwhpMW6N5D9fqTdUdx0uH3kZ8v5SseMjE5XmAeNe
YnXHEa+1AuHwQXwUtgKo5cDlRKidSRjT+QQyio9Uh3mj1x9Cafc2vqvYbxIWFhHr
X8r+GBSPWGT+7n3UCj+F/B2syX53wAPSXohp8ivH2lCkSA8r4RB0Th/S7qsA+uzV
/sbNQ2xPmFNZmts3CNH7hsPFinO7FLZMV3SDVnsfiTxz3ATqNbcVU82Wq4QJjvS4
8XOrqrmhau5BuiSazA0D6Yv+EWaMbfLHZnXk157C2XqCMXT9LLlftXXXCQV8jLTZ
FFWW0urzOtDDJnZ+W32JH+iYGg6XDd1EEtPJ59hzv0DYJwNcn/RffDssStyF3y6s
zYDp20s8/PL26aS+jw3BiGdIJCVEFJaFAnZmtiZxttiKosC27PeIRmhaeG5MkBBV
bk9ac2wCIeplIktghD4Q2E0MTuy7u/XDs02NdNton8pBX6/OalS61+RA7a6z1Jfe
fDU6p1uTSWp9pfJj+jy74ZaeAx36HubF5Kh4RlmghEi1MlvxZhODl4qq1ue7b6uq
EMAYTZLcClysotfwI8AFLpesLa+mU1qBoeWWP2O5mmMAEvux3HNMqHQrF8KxEAUT
UGXIRcMeOhHG3LiKht7EnSTgKpMtevF/u0CguW3YE0AYnQAepMtkbsU6dFvFPvy2
Bkwug8XDzm/ozaZPwO5FWDbLELt3+VHlAoek21yGRmORxCPjOa5r9knQytdlhwGG
Klus6WiaLnIy7JXsr2v/j8T4rqFQ8zSuGakzHRT6xW6eHHiK9Tk1MKJNK/2+TliT
AjtRNHCOlOpG2QMT7w51ln8k8EmMxjmvwct/5Nhm8sqE6G4RseW109tNZBAXuOdj
qB/z+FEDzrohV3j+6Lr61TviyxByHj8GRiEb/fc5LZyefXJedrIyyxDOXcIBf8aj
8ANjQHM5yUuWNoxa45qLJeSf7MuPMDk8VWynilieYvY09mzb+/Khol0+T136OYfo
OWwgUMpxqktGpdO3aGMbJTdU+klrZPjYnTxmAnN/RdrIRbvOJkyK0MV7J4F1zMqd
YLoNLV7rBD8bs/EFKZg1jdeTbKDCdSKcMLaZA5polJ4oyMHJ4bMUeBYCZMRQUo+t
5Umoa5UW1jIwJUSmk7PSFoGL8W/r+voaFOh1e/SYRWygLdZIaxK9g9O7gx5/pdXl
i5Hhz50pxiQZXLtwSwJX3GzPsfVfaBlqCak9TpW5Op7lr6eLyyjhhmdUbSboAmW6
+VaiIKRpxKsc0SI2SHlcopEFoPsnGjf0AxASiyZA88GFqt460VhsXC1RlzamoQd0
9UMyPk1SZzh5UjKWfxCI2rpBS1dnFHMBlvRN/B++k+dx08W27OtD7H+NqcQ8MNaJ
DqPiElXdViAvWe39qMHZzm+CtlfSCPKikMcNlSEMNZA8q+0X6vCWzvLD93Y5FOfL
DjGCOWUTbajX2rsb0iZ5J/L+OOBJMohKTSsqR950bJr3OEGkmbs6Lyegg860iL4+
jf0i5wFhKbHGq511hAeMn93qSBmuy3HCjYHMcC8vdSKR9wdgYIJuFdH38SFYtwlH
RaiEK24PW7DLf58rIbLIG6iHOfOt3mhNjKCaWaLdO/0p2Vh0hMt47sBTAZMwHazD
eORykTLM/WW3MaSrsYDpBMWb4eM3C/EeoRpNsrIjNwNlSyuMpM175E712vTtA8aN
0pTQzYtek8hWXRs/tzIurLVqw8C98I7pVrP+ZG0kgBnHsAYLzFqEEm2KeP7yED5U
WEE3SZdFNab6+nWBd/Zuw9o0mBg46wl76yijcCx88lOWjtg7Cd7T6BWjtDTUrFwA
YwQmjse7j5f/7gV2+/igSFlgy06UBiFWpk8H0xCsxEcpy5OEx4Diwmt0HafegpSP
SnjUpVKK7M8QLgWhOaNVWM7oPsvDVc4drFpfdpmLCHKTfhetFhiDj/pMGCPVQkyJ
kAva6klka5LN+OGXreF6MqOTF8VLAsA/SVmqnm9bZIeqUeYlpYr4g9AA9SV3LKU6
8FQMmlRHcxgtu1tXRReTV3am6sma6ZYVw1oh3E0LCOsTJaCSSl7r8mQJ7kQSqpIo
exWEUZEjX2CZ5cSM7mDLixxx83xlkaS1uzvJ+KXFBrUD9RYdvUMgrwpo0IEM5PT8
X3fDjgUkJUVZDpq3mrTv0GGBQAZ9jjUzgie1URzgFGnb47fhxmlwZePxlWBRMVDc
MAhKZ7VmUQPBWi7tNTzhM7WR4ed3JGE4TiVz6NfUU87TlJ/ZSRiXVG5+cZiV+N0l
j5zR9IYZwLrMjTmJLpzec1motAc3FSpgJl9WuoyWl15YbXpLI2cRpSxHX+YSQPET
TEJh1Vb0XDXebi3bexeKyqE9QR05688ofvMsr29Es0b6965CKRRB5jZgU+ukLko7
12SSMOo38w5uiMwygpe7ynS04nOrzwlIgDHekR4yb18y/x+hYSizICpXQnPh23k2
OOcWJturQBxkVPc76aTflaCRnaWyJEk8hegR+CgAPwu+x37AnHyk1NNpO9bTaPJC
SyjD8jDZMRwobl2G2yG29HvTZ4By6KSgffdgrwescm5Fy7lZWkvwK+0BcEzBYzml
vVbiFqUiZcjmNoxW3l7KRqEfzAzAiyAwfu/NkQFOuqQPKq3TQWBbHjvm8f/mMnAx
ewHLKEpu+ccQeUFC5O7v6qAiRhq6Fz/GPMrcAPwGvB94tMd7k3kDUrdyiYhSdd/R
w9QKqxZXJXQwRsUk6ORVmTBySs99x7OKNTIZ8gzNwxi/Nb4HbXIIRafvGAs5HFg8
EWepbchPt9O4hnZXHlI/EE/3s1SeRMTJxu9megHiEqZDehAleVQJfL5QnH/wa452
/Ix145nlacGBt6KqzO6YUJBMUsyU6iOiVoWKJ29fRcfbkbdVvZ0xajpfeiQolpBl
H4BYdg4S85Z0O1dIpQ7QPfjLEpLN4RlgtQ0lwvwhAoSgRbbDqMYj0h606uBwNAg0
JYnYj6uJF7RRF/VslqXYpyXNlF+zhVMoFPejPQweA6l2qZW630sJu9ni/a6bRKC5
CFzuUWIrBHkfPPtkRNMLZYn5AjPz3O5Iftk74KXQkyilTc0YdtgZ+hdBGiiR3zAf
cozLg/FQJd3tNFjKE1aIsNM4YDOrtjKNi3dzS24DRW/Tc4qOoiNxzL7ljZmisqGY
UwmWwCJVBG3ldGOC09iuhQuCEOOXlFY0e6qf4hYOcH89f8DUAML8H3fMlP7WWP9F
BKHoF+Gsh/IZLQZlFjMrrylYgVL9DHKjE5KxSF/RFMDr8dN0SpKGkNaZAiduBrTx
+qNvOO8zFBUX/8ChA1Lyr1S4rqAYyD0bfBkKwyUGDplADHLHSu4aCknIQxk/UBZi
ec5sxzeIeR+RYCdDewXkkq+myPJZBatZV1qA3dxgwqSHNp4KGDDsUImrOWQJd82G
ii9+DzGUZ5828Ya2jhLL5XOl+4ZfqoCswCxNmtzFfay04vKoPlrLZX2NPvuX1oY2
6S7aR78aWKvmokPjU2/Vp6vTtTlgn+hDvXr13WHiRugD6lKPyGUuIOhACbPHdgSk
qO7gCrkceBmyBcIk+nHGkoNnhs3lU9neodu9GsUY/T6OYTuqG6bJDC1yLBwIpDcM
xVyS242gPVuwmvX072xovT3/oZhX776hmVf6aAjK43aIHuUlqRIr+0GwXY+/oE5u
dj80fk8KCCFNChTtZH3llygzG26NIWOF55uTdOAWW97D2Rlk119qs96cR+fhUE1c
ixTwoBWwflc8vhIspsIH8S8nb5hOqOspDJJVzctzZPP3qWv153bTXAGsW/e1cqOb
cWZtSbd6gPPYVgOnTPw0ydWL4rd3BxJtxhkF3EiI1+Iqqh5bsByi5f5dEeSUYd/n
Novt8r/01emh6aTWycEvxEgrf0fK2G7k4z/oasZnNQu0eYWeeYaROk/tvzeNZM2K
XyXwzZAGiryF/C2gNrIYu8CBsP0lAPNHyhrr748YhILbfLVEY1k0gkNoZmvUg+hf
FEG3HxAedyQkjDQSYOSeK/sOfbiV7xecv0Mv7l3hMgS2gY5rmVvWRmHjgDORd4Ay
gSJaiWESbHfmi5Ew3KrNiEGLISW4gAJ9YnTuflWX7jHZfuQaE2R2l/k79fF3tKEZ
7ef2XlkuvzF2X/TfPl+v0soK5wAW/iZGxWymOhGRB0uUKEQcM8cy4HUJAh/ZVwRW
ujei5k1KXo5cSba8FWTV6qURRG3+WPJHztcfwpby6cBjeFJ2ODPcyUesV4CJDsmm
VZ5LlGYtQAtVcVcp6cpHmuM9QWG9Q45/pFXTwD0BZxbisE9plixq4z5ZOUyCDAHy
8U1KKClayhczHTZZuLig3vPloR2rg29W6kKa9ByrMVGc2AaweKN7U2pKW/09dYcj
eT5uyfGNfQhRa/GE2ijj7f9ZbR71mtt6gOlmDAVISYKbHMk9ucQUCbceYU/9uYOs
7EDRhc+XERtKQhRSJtD/Hkk0Cxm2V5N7+KSmTWnlFke3v0B8l7gHCfEU2cwzQWGT
XJ7ca1fioTRRr9g2wjkZAVcis5KrYkM9ZIohAqpe6l+Lzw6PJmR2M+fpAZeW5o+9
FVsI277W95cj+M1Dr/PcIBSmLuoQYSl+Wxc8EV9GYueKPRqKpScFWg39IzuXQMxd
4xsOO9NvaZJM3Lb3gXGW7WrLJ8M6U7d5Wfre1ZRp8K8f0OEy7P9lydIcJ5p7fD/e
/Gg5igEgbpHnjL4yELhxUIBVYKKyQeoGTmdbCrcuB6WpTzE+mRhvV4jKkirb59Ve
D6llx9a4s2evKfkMZwAq0ZOK4gwS1//PsmK8Wvp4VxrOkjEdM3XwMbm09a0PpOOO
WpThPSwonljni5AwZ18JfS8DatDlGjoxZXiJRM45cXpe1rdo1VZymsheefkTEgXb
gifqiEp3sqAKysMGcKcBfDIkXDv+Th7cf8WfS976f8SvJcijwtsVfX0nAcxEc8CN
NO/sogyl7B7rrn4d3bEIFBgeBzfk0JWSwXvshnHUCgbHkbT4IWqEyh5ypb4aYWSt
hnm4lI8mE60QFsJP5DaFSRJloPsIHz+2dj7VSxDPXqk3pbQWdiMQkSgLC3iPOkO4
QpxEqo8CTNJXjjdmwU8ijBrHPbMyshfP+eU5KKrw1L+Bmiff3SGwFHi8CufatTCB
gAQOBA0tz11+jced7Sq5/6VDUHk4FWoxcXAGLzxBNvSXwr6lw/YtvvYwpdx9N3+V
t7qh+mQEeJKOG9KbUKEXMvVYyjtebtX8rmXe2CEx1aCt0GzeDht7GzAisgXZJuPG
Vfi+RSbKX8Plu6WblfWGPf/e4vpH/V+WNZuV5ga0MPUqD2IAfQTlcpd1tN2H5gj6
zsGxSPUWHPvt/fUD2cvpWp0ZC3B07VRCcSEDtSNuBa4nWYwV/HkwJmOBIDZri4J8
usaSEMcK3hU3Qkqvfqn/SUYjILjhp9dkCcxVv2CKQw1rv4G57BBhOX+RkGJRn66X
CMswris7rC2SiDD4g+//PTve+NTLRw4bm4Duv/zBhMD/hXQwRoyFPew+vYXYFOfv
5dz7D0ZpWF6MW3Ta37m6g/tr0PKVzdiqFcdbucNa0CT6pag0F9o0cqhqQS0ac5i0
RUb9kkdML/VCLGAyeGhM6UtWvJmYrNx+UQBTSSlO0nq5VRziPXuscI788eWxc4e2
MlPEzWoUFximy/FteyIUu8YP9Qsw9FcYayZuCTPnebBxXk9wfTprqaJFAcPWPAoC
uGYG+rgjBp0L8eCBmetrqZrUrJlrt3Nt40QUK3lXlccH591molwYEDXbKI8S4W8S
Mzu1XW5eLDmLFr1Bls8vEi6aNNDig1EL/giBuBMx/y5ANMwiIH/qyupEiiqclbzl
NDfZiHkTrTg8BYUaZo1uEuHsxWztRuJTsrHpTIWS+h//1zalQ2Qqk6gfPWjvle3H
FtwAyz1gq7szOUzEtdBlyqiEIu6QoaXak5MbO6+ogHcsoyoy/gD97YJ+XaM1OfXC
MtYo3VqQ9aGNxmeVz3xmZOE5Mn1Sbdzoimj7ry2/fK018KgFePcShdITN0vNaFTI
2FWPJ8/CFUczPCUxrb0qFxf6PVp8n7Dz+MuZZ+oBhDJvYx9rm7KDfvvX/tUfRGQN
zTseG47S72Jp7ch54BEXB0iti/PuWm+aNJzCyXY7X+vERt9FEdS7UkoGK86lpxmm
411KaX/PYwejjjifh11USe8x1SIZ+NoS4BFsdxqGq6ltjEWBxDu808TsiWaHsmu5
EgHG94uYlvfqGPXzsY2iS+thspcflcFnhqI+7N4JQau9DmKyjTUv7Q4yJWKGIomX
qxNXSO/3Q1vpvynAr2xaASS1C5McxHZTLFE7bn029skhd6Ofy4AJ3CQmoCu3Cfga
yaEFTKQ3wHibiECSxDYoMt/KYvyoTLu1/alq3aN/MS1Y5LvN3Ej3Wmx4BVyOSEY8
P5O1Klk4xDPP1xNHSLMFDt7xYody6Oqn+0+93kp19BWaDl3o2hFQFiMlqocn4KM0
gWxgSjsaiXxzjTB3Ev0hxk9kiMVcVnuaeVcGy/ORMSoFzZrzm1Xfpvj9UCzBd0mD
1G0pyPxuiysf2NiBhwlItaRrIv5onTPbYWdvGHAaSHRv0I0ynq4DUex1hk+QKyyR
iyh9aBuJLJMuE8ESQr3ruyP+bzuREl9saTnFAhMZ/V+rHxwPCP2F46Oyx/7Z+IPM
alOzFonQzOiwZeV5vsZUZej3bKUM1KsAwk1glN/NWYdCsrSRMQkztHufmqpcFqdu
xiWpeGV+GKXehcSFNTIy38DAm94jdQiRaGgzqAypVFxC0VxlDVUwPGBxh7+dPEw3
6OQH+utdLrn2cpq5io1v8dPaN80fsgCTuq8JMSz9SldVFhEHNiVy9RO6PWHzBJO4
7YIvSN3dj8JTcd67gsSx3f1dKc5+ZGqNSEgKMj57/BpuQkV222G1Jcsva2HBb9hM
w3/JADpihg10M29kOn9EDT55JMyTmhor2Yp3S6JasDzNIaJBwLJpG8hMS2NR9PEy
qvqQZOYFdqpXPB8cLOz85JCCPlae6mr7PgppE0DvdxGfk4sMxjmejlAw5ZYUAehp
RY/dhtC6ARhd/5n92Hs6HYHGaLiSUG+fKa7k5c5/3FH1sW6CEgODDf+YkOTjPNjy
O+LhST84ikBK6tjFVJj2Ejlexm7ocjmv/KvV1ISl4NTv+8OdFmasWHISi2PgRCL6
MyOMy4vrgMswhdVYg2sqOOkIAmffS/Dwam0ooUouZz6MbE5cRqfLpJFoRxeZAbqo
e0F2G0UYuOoLr2BU8smOlDDxHQK1LV4p1XDGnGBgfgmc0MBfH6FYHs0dB6Zh4r1Y
Q2n9sVCwUXSw7R8x4l6pJjZIIFtCMbGBnnt3En/1b6V5yxy33hcwU5wk0rgPL+FU
cAi8xQGEK0jCrmb12vqIK8FwuMK6Udjn4pjyzXR/xpXVYzq8u0cVi/E+XP+wljuI
p7qkievpuR3kP5sVxxLEIMovvgIC0llvvjcv/gIad+AbL+rnpyrEJmIyBYLXYntA
jcXeZuKXgU6TVC02jXdTcY4AVTvReDaUTGorhiyqHWDVn2W3wzz2XcBqDqXsuDvC
pQ/vxcsXf/SytEz/lhTC9pY9S/Ug+LKFWz+1G8864EUEBQRfgu7nOu8GWJ5LYBdm
pyQ4tEF+sQ91/rXs6gpAL8LZnBaBiqSGOR6Md9kxH16pzKveulIqIPIT8M5wRYBP
w5eIJsuoDRwmLm7+cm5WBjnDqhSO98pMYAUBbTFudCB2g0w81NVUjxOKF2+WU1CX
CcJF+K+glv8YnpFfBWFLgtOpAXjnd+SairNUVgVYkdnPgS+h3CXsKIqjMwBHTwYc
9zqGfOaxWhl2xdurrNaE2Fh+JuKoRc3dZwpNtQjY6q3pqzJ82YrnyBYR10qb72N6
fD2WoLRzAsfdT+WCQFxjEa6lnCeHUOnJWpI+dbnhOsUh36zuCfV7TEF8yv3ZncGC
ONVIV9V/vzn6MMytr7kWvNgcRqaTvBwGhqUOym0ihKSZk/Ffu75jWzTJezOmNVnz
wSIH0trVtMxSPFfP3whNbSYS8yXK4Orqzo6sZmoQrvBzRYxckxg9J6erCuXcMetW
AoJ7Pp/w79/mSPL8aJw2UdvCRFmLPVsHx3ZTUruFYcajUnC4wUZIB/vMPIxojvVL
00RYfyUDp5pBVOkmQhplULX+O7Ofqtp3yiyK5j4E4iEWZ36OcoAIMcFDeueYqCoy
Zeqy4B/6r5RKBm1OJvzvAXaNk4JL9v22oxISIpT7KBQuI3UG2HDsKlYkhaIbCEJi
tO5/lbiXAYElOpkR5kFblOfGmIC66IlPIFlD1ytzW+6BFJQT9rZdiAEVgUElDhtE
8Mlpjn3GUChA5sJbXvQlW4P3+z2w4vtrB5dbpYTizAn4floiS5jM/EHPIByhH5AI
d37s3PbidvLswR6yZZyYLVdvTzfZcSd2qCvEhrJyeMxk/0o4Cx/xQSNzJrzI0kYM
my3uy56AvhagSkOXNbbUPZ+BtQV6mnezD6cOzc8ITaCFtANGrRNxeogObV7bkY7z
tIjDDZv2nNsxXkIjZVgmwp/L6MdLoliyOHo6VXz60VGZqlP4meMowIo3dQ9tiwES
2Roq+OUyUn1CPXPAoTLA/rTwoNMQfOJvJIE3ewgOh3JenfRSnJ6nlXNn/hHA901U
p+wMFpm6S6EQ04Bxp4gCznXFwEW0/vWP/j6YMRw1RYaC+JACpeognLEoVEWSVebj
b37CvheKRIvz30NSls8hZ0ktuwdxc4l96IlwWV44hHRkfaBYd2Mf+/nORn+iHRXn
s17+rZ/ApeUGh/LUrzm5e7iPmzy9tn0n7bb0FhgHtcptGLEMBy1j2rh4O4yzByZN
46zvXnvK1oLdYphtE0uYQvHLO4U/X0tTblDF4l+6sM8bLdPRKEFt/3+FRmocki21
W7IdDp1HoK08keyiJ2Q9ZvUXWeeFjxSc6oh5JFYWt31W012VJQy5kBPGicKLnJDz
OcBG1eKBePPfRPpnTjtXP9ZPJzoXFwiEUaBeOCkGJgQhBkd4+JojZK/++2EEyys9
bz5zU0H2KUFcU/mTlI7pUhkd2ty91fNeTRqJESKFarEb6NNOuUyl8QzacOh1OFlf
eWjXsQdBiwNoezpKRvoxlBsTsJOGIeVO5ytYx8X/SzxI59Nt0ywUPHQvm0z4hTss
PD+i527uNPfK08CMd7FGYzwk170pqyjaVqZ82sQ2splYhHDgMZ7qkShMzyPZNuGA
UHAfJJGIFHBmSZeKBkasOhWTm/UI8B3VmiVhEEEFvwg4hUcYOhuyCYIPtQjx/Nl+
SEP1mKaeaN++sQGxrYDM1hFKkKLHQJFPECpR+6c1APG2iDZY1iU+TqVm3yzC9PEK
f3mDozUVCeiYPWcnfE14OzZB8ji5PZboIXk7cpUUJI5SMPQP2E0/0XrYQREvb+1J
37s2PcN8E58OtYH41TVMevL+MgUV7YhsjhtsnwbbrfaX+MnhEbUe8EsrdsM/3XFH
bxdw+ukj28RssP9vJJYlc9lGMAa/HGyQ0/xOn35iTEgCNV7RojFlzHU1+cVMHuxf
wBaPL16e8J8Qzkl8uNySSWUZiStTVyrnHGo/IPzl7sUDS9/l6ZPFYyIrFbvWR7Nr
RhXh0Rv8gjyRPlNeNmkrPx79HjXUNKPVlXL4xUzRSE2lxnwyBQ8azWdM1Nw0vhHW
iYp+lN0yx81Y4oUhdvsxcpDTlr7NU7J8dGx0JXvm4GIwlU9foQHtMLeipc0gampq
Qs1MHIZdA7dvIlnJfkj5gUKJWV3rDToMdLTBXaiAD+VzUwnYEdGbJ/iHGDo9NIcX
W4d0/6HdOWt9eD5OG7yEhVxG6dUasT6c+XlTnyDOawsg54TQoJgBbCqFaGbZNl8W
ZIDmmI00dx1OHNtycz8oTal2VDiyzEEZHkd1xPYGJXCN9qQSLWgTDkkVniMRrLh7
vLvlCvSJNogpegE4ZFHMTwP7vz2FVR5uxtVgORC8pOk3LUWY4BUu9g1/SQoLe3t/
4SSopK4y6m4TI121ksmgGlzjyIVovRXbW2A59RVQmENukABqxOwFVC+IfvqwKax9
AhXAhZX3bxGfjCDNdhM1utkT1XWcTQ3xo/FbTSHisiHBDcHj46Tf2Y3X0WAJKN8v
B2r+zmmx89OTng64nfcdQ0NtIPvvBcEu0dumutnztiEULrSayvXnRuYgdcvp3qTI
O9M5c59gAt1kkzisLVNj+dc2sGLB3lyXqX1SJ6Blqir6PNWSygqAoQG0ULoqdSim
KIeddEgj0Txciq9P1rOdTtO9p6Azr6ys1NtJTjNTocj/bAfcM+rQ7t+wXNYNyQUr
SbkE5v4hp8B2cQzE3F500u5fD2tdJJw4eRs+lgzpXzQtlbo30GYy8GuFEBCU99VH
vJfgWA2Z5MDZ6Lde6a77bNNM1qvux7ULk4IY6BwqIZWzi3T6d9e0medefhZP3nBt
ve95LnJ/GTtkjnKfCRO7J3Cm4V2Nd+fDQk8jnBUP6/hKFSBy6HrF5pKm/GNGZNil
yBXNm3v7fX+T3XRUpB3L7r02M3Spc/KxlEpDhE1dtJAZJeUaybzrtgjC3zfZdSRt
T2Bb0hgRx019Y1Eyp1jpaQXHODluPd0X+Ly6MSXWOJmIzDozdOd7mICzSwJvs8QW
k0g7vDzsI/+CZbfT8cB2CwVmtivD0hzBeK3hpmbLZ/nHHAoHzgtj3NCDNksrI76b
sJJebJ24gd1LucQ6QxI80HuOabmugytru6QNanKOMCjrkuLq2oaAgRuFYSOJeQRG
JByfMGuM5KsLJf9+m4GiGGndF29esYjeqFJgB+WhBidCnyz0bTNBlVMqJ1Zb9qJ7
g/qMipECl+MY/9Sld4CuEZyuag261TwIY0bZ0QbKDgT1FCKOtAEbxtMjPDW++0jt
Ce3RfIJyHiyC6w2LuQVm3ECzU2wjM6hXSgbhzLmrOrkc3f7U4mYzsh8fJEswjSAE
h8nALPF2cXRUfVXO6/vptEWytuKoKGKrK3Sg+LFoK8oCs6Tyf6MwogQq8ElHKprS
blg9ioRlzNBLyW8QdKGbyFFsaGSJ+MqD8SySo6PgLo/kE8l2lQIAQVX5mEKoBiHr
l/Z1ztwfElS5OjdGr9SMVWE15SADy1B4bh+AJXED4PLLTR8kLI64v0hjNappn6pK
JVC8XeLezQRqdBmgwq0dY+AE8BVyacAI210jZJ6jOwiGyABhrHXp2FViw4/Xz40l
luAq5q7geGSUB79JpLzn1z0cnr0p0EZGTmoxdaq15GImk3g8wEi82cjzouUxgmhH
CRRKCY4PY9ixlEDX0F+WNfSgFgyUeN/LiPcrpwAw3A2hqarcqi5ZMzSTzi/35LwD
zQiN/qO1+2BZta9m62mluzMQSC/v3ZVIFjT1aznk+9nz+f4OjN6KZI/yR+KK9YjO
FHmIS1+oEHdwVuay85UWHx8MjDmo0X55u0S5H9gZJN/ebxbXnzsE+Bz+UkO0JnK+
3x1+Tm7VV6Ezrn27jT6M9NIB2BI6MMnrS8uhnhcD9LT/cZBtloA21xXkbQeAsyLN
jEZtPr+nm9J792iY5hSE+JZF0NeJ6v424n2ylx08EuN10pcBTuPbw13H7fjh48eZ
HO25QDCHwT09SRnfidBFnqBhBYIFrHUTBicm203x9sdaQRG/dzrMsTWpTRRD9jBy
2V7NJMWOpL0dnmuiqp+zsQFylaGR7XwWdd6ISNRUp9j0Hwg1A3bJGXjctZ5m8goE
AvQHWWx6SMNCHglJwsZ1EuBxs3MkNhYApxASc6/hGt84MeHHvcJkN1EYMqkacMpI
dK2K+vgfQG0EdbFWrGpWYqi/Hh1ERI9fPBD189t70em9bTbVCeXcgeJSj9J94Qg3
ZzPbwYD690bqULnz/2RukeeHOTi9qO1ArgywumbLd+hZPvyPWB6MbVJXVZCH0Fyr
pFXpOMdLMgmXpd5grE9ZBTzmQMfjsXP8ba008nJ1/leJpAIjYdj0pDI2ixIEvbu0
oJWuvK70c53MVFjo/JjKkkAMlnc/VbVcVPmXNaY4Ox8r1aMgZmewVX/Rjc2ych3h
0kX+xPCH/VoSX81W/YbwLJMU+YPnuC7XAjaJJp5oJ7wYn0bJgc//1ecwg8rL0O1Z
aWHEpKys1v6M0sF5RKHMYu5fmOPhei0ozW8ymr38pLvZeddkx9c957qxhiMWvQgU
DlEOniVU1NHxGWfVy+fzYGmFNFpo6Wg1ZwaBMh91RTbcYZ/g/qAx0hQLXWix+phJ
17e6HDnvkWcc77m22/DMUyoBW+CfTNlfZOlk+m1F2d9inLf0+pHHMpgQ0zm04BX1
ciy/iKV4/ILj7LblVv8B7/Pb+Ssj1vmNd/qLP11XyWTS1DsSGCwtYjEMM0/iLbIf
Xn1zz6jHRLW3BiaXHiKbqcvPFXTYVjIerGWByzPYVrtXPPWCF2DdeIRYhoogQ+uj
c55UE6hffQfRqvA4/w6AYcFRzC7VVnenWNR04m1D7pxoaI7ZKU8gyxhVzZGZShY8
3RS8ljyQX+QgZXp8bVcsrV7hieEs7KoVbB+ktSao1PH0RAc7MapJHCUob4Zn7yX1
bWQLcPh2yx3z6g8rD0CitNhb7PIBKEQ5HlCJnpjnyStN0qVEahv2WJ6A98VRZF/q
12jytMjYcIDG/LwiAICG9NRVF/bAGYD8p9JWt8Sg0lH87DAIogIbUcQGFFxIO7vx
fJbOj4fMLcsafOrtO1JGlGo6EyP2sGJ2XeMDkD3AlYpBCzMQFsCgjySQVwI7872O
5zE5Z7tQCmiLAAz3cXGc72ZBNVGZ6IkTj7lV3jNwreJYN4ZP5ZCTbpu6cOdzwzg5
gf93VYYuQ043UZEeIDVk7bEKXwa3cPnGcRqf1M8zOvb8laSSkIYm+LO+lH252vaX
HnXwjS6TKmqP7JlRcFLUNYkj7XXcQrj4YiaD/O2KIPS25XscG3XhRQWgh9Q/RcEV
CO/2vjjNjndxajILgZ+sQpFopMe0IhonDBr7TNwsbAXqsgAfnN0JR1zzALAU1pvs
yH/dkm5zIGmFRd6wEwjBSsxp1fBN17WU/YuF0+ayjsNFalkqt/X+eJj3/0b9p9gu
8Ry8A1bCON6GOlvQOfIKS2uwO9U1WgZTfVQzs7kYfsetvHbkXZQjwmceqSCiMqj/
78kUzaOGIe3b82+tBEppuUlY8qoPky8Nmd/k8Qmd9F86tOMgeijgnDFhH7rdaSJG
8aeelS9x1EYoxBSTBN6lc+Z1ldYqDtJy+IUE1LeamDCAZD18L8lGkmvuaED1U6Es
kBsH7ekLeG6FwJlJICXKjASy/vBLznD+WyXeRTh1//Kjw0pu0q9jwoRXmoYu/iL2
YiqjzDTqFGl5qJlstOIiQA==
`pragma protect end_protected
