// mac10g.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module mac10g (
		input  wire         pll_ref_clk,          //        pll_ref_clk.clk
		output wire         xgmii_rx_clk,         //       xgmii_rx_clk.clk
		output wire         tx_ready,             //           tx_ready.export
		input  wire         xgmii_tx_clk,         //       xgmii_tx_clk.clk
		output wire         rx_ready,             //           rx_ready.export
		output wire [3:0]   rx_data_ready,        //      rx_data_ready.export
		output wire [71:0]  xgmii_rx_dc_0,        //      xgmii_rx_dc_0.data
		input  wire         rx_serial_data_0,     //   rx_serial_data_0.export
		output wire [71:0]  xgmii_rx_dc_1,        //      xgmii_rx_dc_1.data
		input  wire         rx_serial_data_1,     //   rx_serial_data_1.export
		output wire [71:0]  xgmii_rx_dc_2,        //      xgmii_rx_dc_2.data
		input  wire         rx_serial_data_2,     //   rx_serial_data_2.export
		output wire [71:0]  xgmii_rx_dc_3,        //      xgmii_rx_dc_3.data
		input  wire         rx_serial_data_3,     //   rx_serial_data_3.export
		input  wire [71:0]  xgmii_tx_dc_0,        //      xgmii_tx_dc_0.data
		output wire [0:0]   tx_serial_data_0,     //   tx_serial_data_0.export
		input  wire [71:0]  xgmii_tx_dc_1,        //      xgmii_tx_dc_1.data
		output wire [0:0]   tx_serial_data_1,     //   tx_serial_data_1.export
		input  wire [71:0]  xgmii_tx_dc_2,        //      xgmii_tx_dc_2.data
		output wire [0:0]   tx_serial_data_2,     //   tx_serial_data_2.export
		input  wire [71:0]  xgmii_tx_dc_3,        //      xgmii_tx_dc_3.data
		output wire [0:0]   tx_serial_data_3,     //   tx_serial_data_3.export
		output wire [367:0] reconfig_from_xcvr,   // reconfig_from_xcvr.reconfig_from_xcvr
		input  wire [559:0] reconfig_to_xcvr,     //   reconfig_to_xcvr.reconfig_to_xcvr
		input  wire         phy_mgmt_clk,         //       phy_mgmt_clk.clk
		input  wire         phy_mgmt_clk_reset,   // phy_mgmt_clk_reset.reset
		input  wire [8:0]   phy_mgmt_address,     //           phy_mgmt.address
		input  wire         phy_mgmt_read,        //                   .read
		output wire [31:0]  phy_mgmt_readdata,    //                   .readdata
		input  wire         phy_mgmt_write,       //                   .write
		input  wire [31:0]  phy_mgmt_writedata,   //                   .writedata
		output wire         phy_mgmt_waitrequest  //                   .waitrequest
	);

	wire    [3:0] mac10g_inst_tx_serial_data; // port fragment
	wire  [287:0] mac10g_inst_xgmii_rx_dc;    // port fragment

	altera_xcvr_10gbaser #(
		.device_family            ("Stratix V"),
		.num_channels             (4),
		.operation_mode           ("duplex"),
		.external_pma_ctrl_config (0),
		.control_pin_out          (0),
		.recovered_clk_out        (0),
		.pll_locked_out           (0),
		.ref_clk_freq             ("644.53125 MHz"),
		.pma_mode                 (40),
		.pll_type                 ("CMU"),
		.starting_channel_number  (0),
		.reconfig_interfaces      (8),
		.rx_use_coreclk           (0),
		.embedded_reset           (1),
		.latadj                   (0),
		.high_precision_latadj    (1),
		.tx_termination           ("OCT_100_OHMS"),
		.tx_vod_selection         (7),
		.tx_preemp_pretap         (0),
		.tx_preemp_pretap_inv     (0),
		.tx_preemp_tap_1          (15),
		.tx_preemp_tap_2          (0),
		.tx_preemp_tap_2_inv      (0),
		.rx_common_mode           ("0.82v"),
		.rx_termination           ("OCT_100_OHMS"),
		.rx_eq_dc_gain            (0),
		.rx_eq_ctrl               (0),
		.mgmt_clk_in_mhz          (150)
	) mac10g_inst (
		.pll_ref_clk          (pll_ref_clk),                                                                                                                       //        pll_ref_clk.clk
		.xgmii_rx_clk         (xgmii_rx_clk),                                                                                                                      //       xgmii_rx_clk.clk
		.tx_ready             (tx_ready),                                                                                                                          //           tx_ready.export
		.xgmii_tx_clk         (xgmii_tx_clk),                                                                                                                      //       xgmii_tx_clk.clk
		.rx_ready             (rx_ready),                                                                                                                          //           rx_ready.export
		.rx_data_ready        (rx_data_ready),                                                                                                                     //      rx_data_ready.export
		.xgmii_rx_dc          ({mac10g_inst_xgmii_rx_dc[287:216],mac10g_inst_xgmii_rx_dc[215:144],mac10g_inst_xgmii_rx_dc[143:72],mac10g_inst_xgmii_rx_dc[71:0]}), //      xgmii_rx_dc_0.data
		.rx_serial_data       ({rx_serial_data_3,rx_serial_data_2,rx_serial_data_1,rx_serial_data_0}),                                                             //   rx_serial_data_0.export
		.xgmii_tx_dc          ({xgmii_tx_dc_3[71:0],xgmii_tx_dc_2[71:0],xgmii_tx_dc_1[71:0],xgmii_tx_dc_0[71:0]}),                                                 //      xgmii_tx_dc_0.data
		.tx_serial_data       ({mac10g_inst_tx_serial_data[3],mac10g_inst_tx_serial_data[2],mac10g_inst_tx_serial_data[1],mac10g_inst_tx_serial_data[0]}),         //   tx_serial_data_0.export
		.reconfig_from_xcvr   (reconfig_from_xcvr),                                                                                                                // reconfig_from_xcvr.reconfig_from_xcvr
		.reconfig_to_xcvr     (reconfig_to_xcvr),                                                                                                                  //   reconfig_to_xcvr.reconfig_to_xcvr
		.phy_mgmt_clk         (phy_mgmt_clk),                                                                                                                      //       phy_mgmt_clk.clk
		.phy_mgmt_clk_reset   (phy_mgmt_clk_reset),                                                                                                                // phy_mgmt_clk_reset.reset
		.phy_mgmt_address     (phy_mgmt_address),                                                                                                                  //           phy_mgmt.address
		.phy_mgmt_read        (phy_mgmt_read),                                                                                                                     //                   .read
		.phy_mgmt_readdata    (phy_mgmt_readdata),                                                                                                                 //                   .readdata
		.phy_mgmt_write       (phy_mgmt_write),                                                                                                                    //                   .write
		.phy_mgmt_writedata   (phy_mgmt_writedata),                                                                                                                //                   .writedata
		.phy_mgmt_waitrequest (phy_mgmt_waitrequest),                                                                                                              //                   .waitrequest
		.rx_block_lock        (),                                                                                                                                  //        (terminated)
		.rx_hi_ber            (),                                                                                                                                  //        (terminated)
		.rx_recovered_clk     (),                                                                                                                                  //        (terminated)
		.rx_coreclkin         (1'b0),                                                                                                                              //        (terminated)
		.pll_locked           (),                                                                                                                                  //        (terminated)
		.gxb_pdn              (1'b0),                                                                                                                              //        (terminated)
		.pll_pdn              (1'b0),                                                                                                                              //        (terminated)
		.cal_blk_pdn          (1'b0),                                                                                                                              //        (terminated)
		.cal_blk_clk          (1'b0),                                                                                                                              //        (terminated)
		.tx_digitalreset      (4'b0000),                                                                                                                           //        (terminated)
		.tx_analogreset       (4'b0000),                                                                                                                           //        (terminated)
		.tx_cal_busy          (),                                                                                                                                  //        (terminated)
		.pll_powerdown        (4'b0000),                                                                                                                           //        (terminated)
		.rx_digitalreset      (4'b0000),                                                                                                                           //        (terminated)
		.rx_analogreset       (4'b0000),                                                                                                                           //        (terminated)
		.rx_cal_busy          (),                                                                                                                                  //        (terminated)
		.rx_is_lockedtodata   (),                                                                                                                                  //        (terminated)
		.rx_latency_adj       (),                                                                                                                                  //        (terminated)
		.tx_latency_adj       ()                                                                                                                                   //        (terminated)
	);

	assign xgmii_rx_dc_1 = { mac10g_inst_xgmii_rx_dc[143:72] };

	assign tx_serial_data_0 = { mac10g_inst_tx_serial_data[0] };

	assign tx_serial_data_2 = { mac10g_inst_tx_serial_data[2] };

	assign xgmii_rx_dc_3 = { mac10g_inst_xgmii_rx_dc[287:216] };

	assign xgmii_rx_dc_0 = { mac10g_inst_xgmii_rx_dc[71:0] };

	assign tx_serial_data_1 = { mac10g_inst_tx_serial_data[1] };

	assign xgmii_rx_dc_2 = { mac10g_inst_xgmii_rx_dc[215:144] };

	assign tx_serial_data_3 = { mac10g_inst_tx_serial_data[3] };

endmodule
