// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:12 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RHrGhyKKxqrk7clZaDLJ8FCWMYLucxWVmqQzmD1M0dA3n/9XYAVD3PhS/L3awEdD
bx4fekZDE5Zq9R22tAyB59bvK8U6+yMN2diK75XtuwTLxZlzEdkY6PJdw1zychvZ
yL9o6hRELxVXK4UqsCLJRTu7AdC17ZzvI9Wu+GTUWqs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5408)
1I95hG+fmfzG1CX2x8fiBaKJXu3GsbyiXk7ErJUexpNjzBr8DZII7zkqW9g+3a2s
nPc886IZ7IqUiNkpjzAyakm2Lhd451uJjavcK9vPgPESqeWX0olcwGfe9dHNdI6Z
qadHUV4h3AU6lm2tfxsdpSHQ14AzYvxxzpUf49WzBTq4c/yJgP6zn5V2KSZZU22d
XA4BQ6e3oDGiczmaEIjN5B3TxZ4UhxXIENizrVkMD3WTxFeiKs5+U4vNhcdsutqd
EyBdkrnnF34HC+LbTdHAPU+BzOFetyqgl8xcIKt4zq2iQMYrl+0ed6A8i5soL2Em
UzF46TI1PrXc15RMu9Jfp385RYyCmokNoFCufrTRPAuuezQPRkVaTcDCpjgE5FeQ
H/r9UU0jLx/1zG3BxeUF+qAbseRrcyWSi7AcHyPxJX5WCkr2A1gztWf/8+wooy+q
4oa0CALfXlJvorthudy+xxlhjaIfI15xIZ8s6hQyo0fAS7w+aSkncQ08+H672pwz
tX1S3IM5Z+4vxDegKTkekIKsnvSxzk7FM3HmNFmB8iLsyc3scdh6lGneHe8+iDz9
LAwdVB4dbHL+Ywe+b6HRi/Y9rM2z9YKy+E9dgASjlda3hqrheYaAWQOsUguL1H89
832IJlcWE24x25q59SHB4ppHXqWwOthxEt5F9jzbCh+HQY6phutCIJ1aEHNgc9Xq
gjU843G7NF+qWT5Ao/vCwc8Nmg6DGey2YQA/00l+0Wc7JswkZokSzL3PcropTjXz
M+yju//HhhuzSbwrr6uNhbsQQNy9BR3RgRdctjKThFkcoktX1D8qPjfphQ6xoFp/
6xoxYXbRFjI61H9LCpbsXBpj9AGSaP/JOavMxgXLXaObrApDKi5YQSQk7cWcKA3M
ARyI5WGMHQEOmEOops3NKW5phMc2I0tEDOUsXgQfN5Jrl3BwOjw57bEdRbOL19Kr
Gx5p33ncULT96q7nieR3Hk439Cz+ho7kGCiRt/QCS9N1mhxZHi5YsIVCAIEL9LKv
PdHBtQMvvhDyEq3dzzJmGXxLVyt5wceKwkFV8cKglWvS+oZZ2L7D532Vywh+h1An
AfmbjWNkbE3pIQPefFUbm4jUN6Grd1Dq9Y4yXjU2dglcRTcqTNRK0s8gTkemobpz
ludKUvUNjwECzOjhnwknAUaNI2I8grrS+V71u+mW4XuVz9pBJfdN5+noKWLNonM+
/VhTr1bfX7+W2YaCk+HPWi38bhYHmVeoJVbDz+5siwSfYQGUelh4SCa1MhfsY5ST
WPrURhFqPSis0LZveoOaE5QFKXsI/Kw0jcBTqNLrgKxptiCF46LPmXUtBbpnewM9
3jCRC1ALwI9xnD1icgYw2GWOfSEzv56lf9AC41epEOJK5aEq0fCqmvJpStxQOGYA
P9rmAS6pGlaDONkK/G/xxpKFHpVPbfsnjxMKn4FFwb1GrFd3g5IewRyKtibCTbW7
08Xt8f8nJfXff9nMVEqRZKLZYFAZanKZXl/4iM7jQZoej56VewFpJdEg37zwHmVo
qrxJCy3O93FtHIgjKAXujeHs+GC2vqmVOtM2ktJL8BCHePmk0p9N2nwC1FA+cx6M
31dGpusfEyHMyIIbbz9PqkGBUGHjpQ3uukCFqicQ7habfjcDXnRjC8DoOMwXhLcd
goVgCeyeJOtZJBuhp2TMNn8gGS9NaOuK4JGe7IwgWCnfqJ+6o3sKWpYNOIcK2KB6
Sau/5BhmJYvjHR5xrT90eS4nyYBveVqIl2QzPUy/3RVimQNMort4GA39R9yB9EFi
zlEujciCMIaWRj3J/rjSJCkQeM4D7qTLlc4vvb0v62o+o+f0ZHCyPoKAylArCH3f
gULsIHoC8Y/xevTRfG/8PB9O0pPGasuBFxhPDMGINdi74jbmrv8lmB2Etypr07O5
mury0cJnCCqxFzd5QVEBNHwU52BdeAemud4BUhSIWGKyJ4DBUwYVbFzESFrNwBPm
PH/o5dRba2SFtWy1Hy+l8q0TVG4SXsW6DhaykKsYkq9rcQAgxVeq8I09cviRG+A2
ZyzT07e1puSqeHyOmtbZQPaDzr0m/jq/ywz54k3p2xat/lYP0EgKQvNWu4vgxJPX
OcKvAEqc666oJ9l8DU+KAe9w4OtK4SvXJ4uQezdXcvLkeL7X3nmmos0e6/v2DHgG
msh/eV5t0rSCSZRXyY++zni/mYZqUHYwLpVyjrhI9yEUc2OxPUcgvmY5/CkqYS2z
m9/o5GhR0/G2leBKrmhdmLuO8O6dvdsf9s5w6mK4dxpjfrreTvW9AmPbEpvx7ead
J9ce+sicCZ4QSCYzqoJ5i4LUqUFVW0oDVW9vGk90WBzmSMZvfJ9jyTQ5g5+12gYp
CvFx6EpaNf7HAi8xb5NZhCyXc3l8r4perS83y9IXV4U/EpfnujXFtZXcxIly1w+p
ObQsbqEssmnI6C01Nl7WtxMtjUoR/BOstg8W0mJRukJKATtN9zgGawi6R03vutnK
x63hgBUngPBBlMyMcAfmtXrUzORrsk+3DRCtuFGRK6U2V4Dnt6YESTDie4xY8JG8
lqlxdRKgiZ5IBJ41eX9oHC5HMh3Bonsugyr/uItxhqDaqA1WHPY0WIhlX/3jMuyo
/3aAirPYpTFwKHksc6Flb3nrWnxmfLhJz2jhXFoaPe1k0nhcBvprDtS9CLADtKT0
s8arcz6pIus2EEvFw2e898+St9pFdxWClJD2tHhqPdxN0SZbzZ+1EF8PDU1jwPbc
h/IUK1lzNsulyBUaiU8quJtnFNiFW6+9mZ4BXDWsJXkKe/WVPXNDQZZrQ1bqlNuG
lauXSQB6T3yjDlkMqUNR67lgZBNZi4omcovLHOsfakRsYqXdyYs1C0vsFByI5m2Y
qdsJFLT50w48mWspYQYsPJBuvf6x4U04dPMfWMkTkp8GX6K//shQm7fAgMp02zvA
+90EoByf1PtcwvCbGgDOc9FBcb4x6c01IXxXHoLP79FsCY2QSRfMjZIpIaJojJIq
k7yqyFm2xFR/N/PT6xK/fQv9JadjvnN6PvDGf+V7TGNlJvmtipgBiGSpJaVTimEU
XBPv+mN6nlJQm0qVEdT4sB3ELRWtO1Y87/ciQnV5POihovH+xw/Tq+hwwNUye+cK
keM0SoCbdrJqvKHH684caXefDnf5R58LFRplZTjF/gfPoiuxF0dRJqPzuTfZCHgx
5xL7fti8Y90Mo2jzS1eaLqaxnHZR8HvG7WgDsVH/LGl4tONHR7BBaXUbKVT1VzwB
AEu4GsMUdegigUo+TjHPxVy/g2pF7KIEj8F5hajcyMS8NHGgDv82SqnpBqO3wxXA
ZkJiXJxpZZytI8VflbpKDocFGLhZ38tmwFuCNI9F+zzW2Od6NGOB5rxO4BfOLo2e
zsjyPSn6RZbLgFvWZHSKyC3p+J88TCxX1jXCu6AyUTbzSLTjIAeBP6BHYop7DmpB
sqDoVbHLINzh9kIDQwcSK+t5JSqMm+JA/kcheoNjFakvhYi48/S84opa38x/ni1H
c2RWVhV6wDJkaj70KYnAn/L1NNLC21+AjHyPoUKIEdG4F5+EE5CBjyr26RroYvRQ
cGeGtwf+PX2SamJESzwLUCMC2Xb7/CXHqYMB3FQFjDlWj/rEY5iETqEAcQov2JWb
me12nUtryFDqh8Ar53/KmeNRWmRo9XnYCXVvZmIo1D8UBaN0wuVdd5JK6qQzmkrJ
UXjGog1OLy6dfz+PFu9ts1ZsFgV6QKj3tv+xFsn7+KQZ0oaLlbns7mqVBOUWs1SZ
zmDY3sbSmjCQ9gDanOi0X0HDRJo7ouOUIgixrF/uTSw524MvvJCL6/yfTiv09X2B
y8LTpZuZpbjtWTXFTchRl57oovyD2JHuqw5oizMIb3R3r6mKTV86lmjxN+QdiSBP
Dm8ap5Ap0s/BjfFxc8/9m3sMJKaTqR6HXCd4d20O95reT0LzKIhG8XVO+Md4STM+
M12mt8H0O4GeDK48khFKmZkkiYvIPutprISpbPckHdkexBvUPCwKA8vKC3V+Zvoy
lMgp3GhJid0McQ4UAUKTVfHntvauVCVhZbFfTyLgxYFwc1OwA8XY9fKK08fc+5T3
+pj0fcTd/SanANK22oUEXq++Wah9q/MpOa7apYYPzFNaj1g+rIxNJWBOQ4he1OyW
sqvXyoy+AREJiD8ldFvB10VLdntUhPzhDZ6oi5q8sexgRzoj2GataetgrfGjxMlv
9oNETDENHwwD0+CIejHaAEuWhoWEuanXOc+hFNP23Qwr+ssJ4+cg1P13g4EYirD5
ElTEE9etuSVkz1kojvLXR/Lr/hiBxncnGheUcYe7ACv/lnmQha9D1Ox2Ihl/L4Y5
3oRxViwd4PZpvBFhwluCIoRuJSX4ZVXuzs2ukJOvvBSlnKNGC1X68Br+kY1RfEm7
ZnL3d/OGqoo/uqHPXV57WkFGinGprv7kJaj0luSNtDowKSs2WpbY+V8K1WWvMgVw
0V33oIEnflTqKdVHe4FxIXH4Bz9jpMhNIMdMCJ1/2Mz786aU12Fr4iMhDd2OSGva
QmGTJOZe/7ePa5koY/f3AWtirTzYqwnc14G3Y5+VLDp4gwpqnGbpiE9bfXpXkYjt
EGB36mx0yWX3XtJyKD+O0QG9K9/kfPoftXwwBh7TYXRLqA7qCI/JYfOJ3xUBA404
vzEL2ifv6BCJhVS+2kzPiUzongsA2SBLW2tzKwJwzk5KuhGMKa409/RGXiHPJeu7
l5nOhNtyqJg9RIl3gsTcMPmFgUubU7G+M08kTMi/SslQzqkNxvhjiM7mtcHBpY+t
i3ljE0VYvksSWf9/MkqjtDFq2IEgddvqjiBaUuoXN55PKEbQGkWCKAWPFGVU45k4
GatIsp5YVBGplDvbZWieWxhQrQpftrXfW+2Qs2ulkNh79NgiW2926nJ9/oA6NuIk
DThq0W0Wa6t++0RGbi709IACofi7HiDGbRCCxArnS9ZczyDgcXvoVHUqv91W7gCU
nPzvU6vZn1XBa+cN1zTuF+tetel6C7v4kFfq1TP+vxWo45yKhsYkgg5NxfYzurDX
+BlW3OhDTkMNnOlOkHi5tkflDOXvS4e5ocAYLi/17fj7hzXup9bSJEgR6mQiZQ19
idBXyJaZdRaSSjxaPE1StniMWvn9J0SmCgqvJV1QU5QlvYrErisM4Pkul1oUtOBn
sAkzfFe/fu6jMPS5xvmYbZcvwyV6cj0Co/Cg0TM5P63jQq7ZEMWp47SZRTwMg1Zx
irvi37N5rQ0qNoGbOfK4j+Q78DVkpLAbrT/RtAY3Pg7WSTlGHOfDGLFlHwE+KXsk
a7ep51nkCgB63LmJA/Si+Ap9zoav89sSyMk4DiSagCPPF0vA5Tlq0zmIM4HyUqTk
P9Y/rXFrNnhzl4rsyI0dDpFfvDU9rdf5ctfxsft4AgKWEyj5F6K5TWv2Qcqr14gL
jwnO68kms29luSxSr8y4sNdIJY9g3GyNvcUl7TfNu4gpc/Sgn950g5kl4eG37cAx
84Mo2fh05kF6Z/JUgCOx65tYHkoS01mZoy9ZHtxPxSLaFUA8HzauA8fkydRWSjHp
mM/CDKqR+MLfxcj9degf3IrRH6+Djx5cSEgbPZS2gmsPNzJ2TZ2SHR31X14x6dpy
FzSxTEV8COwZ2mk+3jryp/79IXSFX4GW1mhtk6j+qqzrX/R+LsFtI5cNNGhmUBKf
ocmMR0oX5aT0mowmnnuBhSN7kmzO7tAf81/VGW0scBodqlIn9OaGcw4E57eqzdee
fOE4YElXUSdOolklVI8V+kL70EYmiYoYC80ZdFxPlwARki2RU+nRiGpEPpZOpnYG
H5czs/aEkTVQcOBqNqc1KOHIdayvwZSJ+WslrnaGxiPT68RHJCy4iS1JP2a2O3d7
A1PSsWc+7KCI+AE7pgNVPsxh3o2QHk7sWoDwh9ewByXp4ZQKZ6Zmx5lsT2A9BIgZ
0URVoyHoyk3iUGQeQblS5sYz/8EiJX9PJI5pHFnfuf01Pxt0RijsdtXNN360/sIe
s7rYVEIl1phAdGpLTZ5XfmmE7ODu5nqc0vf4i5jF54MudsMz5j8Xmbg4aJf0VRwd
yuR8W7InuL4r8RfmPr3+0V+6Qw2VfV7F6NVKziw7kNRqfC7kZgG+HV7kzVUJOQZU
dgJecI893qjdVgF0wHiqW7a6bvUCdyBj8Q122H0Vq7oyYZAugLGyDPzZZIg+Hbo9
ZpjuF49mILlG4+t6X7ufY4Gyq3kBWXtnjN2bE56RQO373VewQ8hC78+3j2Bo76Hw
zusUefVdxRNJuXLHRHuljb3zGGnxSARAvsrHElbqj3/nF59p98YTOu8sMtyay7ky
kfqYdgdilfgW1KDN1iac2GR4ge/jbPV8jLfHv5y64WjJh+sJZ+iOPmAfZdVwQX8q
OUwMFET1eLfk1fWrgi6mg83HTuqc/0QKUgqCN0QpSCZIbxp0QIphPqrCWt3xZLOA
b127r1/RmM8UjnzPbywMlQcYNpJ/biHWwW0V9/CRY5PA6YT5xHganG+6WvpFRkKN
VcWvM8bfCCfOgo3uwCLRUd0j1HjJiqLv6UJVA3rvraTSSF9jZrj/ul9e1gr3xjI7
eqH0jSZg0ePMtsj64LHgI79PE7BIAyH+/FqcenZ8E6UFNi5jkbJWABcKQT3U8PNr
3+nhHZ99bDG6yk9wVZBdbvYHp+VNO3jBYfREcS0CPglBCgEgKVjKVetFRZvwJZCu
nf3zTbHqtRzLFmfOMrznuxIEqjVI2bfkbGjVveByscBYReNCIRL21UbRAS+rRCRC
vJNhUhI+xZsXgVjb8LuU8U0OZcLWBrqBOLb9fL9WMeAvOCArEKFVMxVACn7qvj+u
zZbYbkQLsYONc5O15aI3yMSdzEqsUM6tQB4Wr5TzNyvdq62gah/0wE3BdijgVS/b
/is8MrQQM6UnySpbRce0bJ2OhO72i15RdiOHL6mpC/S2jqMgzCN+mPARdxEXtG0Z
fpBFh8gMZHtQqyPdFSmpyiv/t6x1VPnGCKiw8XI5Dz3VLd0B9pVSxVkcsVrl8f7q
h966Jff7ONhqIFdGPEoG28NYtsMHV2GK3wRmUK/3BvySmp7yolarSyHp8+jBUfd2
FDbFKq8y/XdiSHVs5aZAy7w0lWaPE5+f1IIpVcrRrQtLJAex4rpVHrrKI7xo9Fvd
WXAybwTeGtWyCk3utujEP2ueWlMXJypffbQTjbho948=
`pragma protect end_protected
