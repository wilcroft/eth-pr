// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:14 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KgilAtnFmy0nSXashD2SM6L/nyI6JvLzyYmkV/UH3bCEc0SmZgIy/DQDXLEbQNqP
AWU0Nh1F96bsfuvouatArmte2j+1P0ZgBeMqscGusuqqOIDrWX+zoRY8MwB1lIew
l/HeaDzFw2yfUOVfETS/zenEaYCON1r+BVaPUZMqbzQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20352)
EdFK1D2bY5b29/jeflpgQZjBcKHnS15xG5wdqhCwM3tmD66D+wIQTk26W3qRqmR9
DeQ3P7b6OCI5Lp7SJBHBQ9s6vcu4m012ebZo6UjzfZgQiPQTzdn2FYIW4LoJ588G
j8NlYTYhCZOAAYuKhObrAqKsYa/JZgfRIxteOg+KrtecjtGc+CdyWpmPYmmjWAxL
N+KN1GBjaiiPthrvg9Y1gpJUxkCB2S+YgxaHEAau1vViD4WhRq26JjpWapJO2qEG
CMmwMfkggpG1BFsH2qzZ2blXJJcWUpE6Ni+gaSuat1Ae3EGi6MQTmj86AlDwf5uv
DmLdzT4sPWCCF9IHzv4swODxtOKw/o0/Hm7rn7qKJueVZ6IxsXC7Xn4AWMZt1Lxq
8iBEBF030pAO3VAijAHoyrYd7aZMSNvjImqayLyXD4x0jP8YkNFUtBkHYdEYbdd3
kZwI4Ex/fQpzbsKnEmsljRJt9PI0uMBQRtiwNSBsQV3TX4AAERu9YZqBHyCU+mzz
uWQmu+VxC5M9BV2R2WsVE0jB+BR3gOZ1X2Eaj/zRQsVSUVVH/t8xFl0FUQkcwbWc
9ajdYDewU0itks3lABQHdDY77t7Dz56VPk4OIP3JbdoWfTYEVVSKg6KMGDMO/8R3
iDJDtLDVJi2jNV2NNsEJe8SgP+V9XtGTX1Ss6s+zrCXpD7IubSzUQ7Tpv/OTYmhJ
LbqV7hblyRhwZN2dDTkG3fzv0QEdn8gZrdPmxFE6TvMla0j/IOsBB0ueIiYpC+5N
sa3NXnvUH8iJYrXyniu3Nc7/bICHjF4Zar/hicshFJv0uXOxwEhVZVIDkLqLtZgT
NBFh69fITK1U1PsMShZYawoMappdRAA1O0JtGMazapnXlRQloZ0Samni8nV1ZF81
LXnVY9XzCpZQD0fAs9CcgeptU7gwXaUJLCTESt9Ahroxzv2ktKqTLBJCNJeghlJv
SYvUlPavSuvP8DdsxyHo2zajP3eHG/GCT7SJYe0p/B4PA3sK7bcKC3f7tH2JYJH/
gxyzwu0Q0FvfSJ0QXMIOdeltuTSzYZqpcSvgBzv+sx48KlR1xD6LeoQxg/SGxhia
8zI1bApkKiyWEBNlTMMxs8XNWw0b1QH3s7Eo8HYOggNCoFOY2wSDkzuTrRzJTrrs
F4TjKJHnhg6/iRPiZV5qRQzHXgcbhYYsSK24W+G/SaZQ9v4SOO+VGv+M/0HXHSXS
IrBH3wzZF4IZ+3eS5HJdnVp/p3H1FiKdVfCNUdGA2+JsPq03pBcw0/1oZ5l3K7BQ
xPJ/oaUlduMWKpg1kjxi5doJ2cZTkdu6dbCFt3nZB+W5ZAuAsLon09WrCgciQkvD
PfmPbGUxLDHCbEM5E+UPSX4CpHN5j/mZBKMgLKxazPQSny1xFBQeTnEmn2oe9/0R
jCzTn09TQo1+iNavN9kOCEf8xZYOeJsfmx9Mc9PcAP/nAqYyNfXCS6cA3wDJe92E
B1E3kz9AGVPuvtB1G04jv6JUJjGCXy2vOsHHdcSb5uLM5R3uBeMTZvaUfmrHcfgh
8qt6lHxwT8TR9hn2U1S2jNcfrY2vgJtVhDr9e/olrQuzfrvE3NbrBqG+uz+tXmHI
LAEl2z8XJunZfxO1rLg4wQogerViQ//d9CT2hxz0GZD/5zgOUOuL625jEvEqoiyG
Jgrj2ac9BVWjh80TRlZJ+m8CnY3+eIAzA/f1Rov6FtkjYcATYxNR6QTItL19dboB
Tv6gxTGiRigDhu1/L8U9BwH6WlvmR/a2ejQEJeWYxnF5iS80XjOo273dEZJ8HvPQ
44gsqGtWkxeso5pk8A35KO12mWBmPQCuuuZ2mrk73OlU69L7aW7Lxjnc2stc44Yi
Q1/5ykPyGczzoYwxFpu0cwh9g0lajQ8Ydnw/7jAYnkVMgi7HmbuRh2I5SqrCK2pu
y99mH8YZXw9b4p0S44pbruBFx0e6kR2/Litf9UVGS5By854cVfPiam7y7TJuaNks
cha0WDwTnDrCMg2o2v+VUiRLvRdImxPdQ+pnvwtKzYijo59sPHAMHhbW3tu3/HGR
rzfToQvY4VVq5FmSSqrvGdkO8H1UeysN7Fg6U6uTjVvZovu0wkxo8KksxrNCYWEL
KO+stMcPE/hj/ljFck5o2Ntb3IZ7+to4DirJ3OxwI2ICRGAZgKeFK5TIVW5EGW3v
5Ko6msKr06A1e8pNumCrGFMyhsNOe5j2Inw233avxJ9PmOAlU8P+XqKg2F0wJhUn
SCzakQN0ciR/E1HZ605VvlanJrQ7oizcGPF8OJHOU26/NiXyBEjI84xczWietBx+
K6qeOkICbIo6G2q9uNZQKKeQlItt07CXZa+PkNOQ3hQdvgyO/ubeqqi8pCCfIRHx
IOWl+HV6Zq5e8ECADiaOWhm+Q2d67tHhZVa3jL9A+Cc25m1voXEGXqZ96hujAGzr
MnogOUVGOUa+oANyMOj+4W6SnPh8vln8BomwMWpyFypXJAmz3FW+Fa/ZH8hAtRVD
ObzyIOmVZhiS+kN1UI3Hnphm8BkY5UfbW/zM6IsBbXiiH8Bcg1oMCntcg+IJ0Siw
cOt3az3eK4a3WRgx0r69f3hYB/wnvuelW+lk058O920qT58DqmnabAMI1nRWGYiQ
n458v9hPZYneNcLpHEMeCvtYPl9bHwNnRPy83JLpL/Vf8ToKLHuc2bNLTbgl2Rii
PEhW6ZUJcQdF61fnaUfuKSsqPBh7s48wCp57+l4IVYZAg2m7dqdFeYhT5mOp+ygP
cdZxlkfdX3EZESnKgyX6+bA/N2tOYawxKzdWq5uUGmISJWD+WVZ0sf1h0LlTyXmn
ahPAL53MzE7iBZpiDM1wKejqyr3LKOWqw9oXF8e3QbcFTcS0ueGFbQOl9lG8Ng1K
B3pn7c7Rc1yQPPbEmCa4DqGjJ0+cMnBBXisYYKY+7d7M/JEfVVfmhuFX2UwpA+ml
brLHGim1SEsBUf1z1rNRqK8yZ4V2+ka89K6OWjYgTYkJUvUVUijQgEk0qnlugF2q
QhNYdeDJfZY8pAaT3Uj/gwRsaBXhK3aAptLALdieYmdtu+uyzc7MKKwCKnBXbzg6
yt+aZIjIKkUFy3WqX5Psd5lhr9HFv+MBMO4KtwXnpiQTkQiciYBepBySmKztykyb
kv6XcZnMzb0j+N6IsNDEhNyYEWbn/CES1u3rfP5LC3d06zhzSB8Yt2Nv8DwsEiy3
6G1ukNWjWl75R5Z/vhtHuzc29MhXvtX1vQ4Klc+2UhlCFBAhLUaLeuE+EmRptLUM
sXDXWtwxF12wNQcrI53sj34/XpK11Khqelj+66VXwX4cQm8xDB6TDVgitmv44iRC
dna4KojPYFbBsQFjcrlcmDJ3zCepHYrdauoLRd77Iw/EpnSg5Gwklv2MuxtuBaFt
NDImSUWRfNSYkjtjQTitZiebR5CEm+RZ6AJkp64faqnfKnMakTiPgbrkNn8EZ5bc
/ONmWa/REQhxrWR9HuncNhQKYBrD2Mwq561q7WTQg8YU3uZXTwIswB03YCJ3iykl
v0y5qj2nODAUKPipEnF/N01Pos+0xShVoGEUVCrtt/U7GqSQpmPqiEDTQ2Rdng0O
bj5XeLjyy+1jtT2LHeISCAbVD0nzh4/PdS7lqXJm41U4xptyoxJcDMnM5ZaWSz4h
JpoYc1c0p06QoOFtGEjupxtH/SF7wn4ZVHQnAF1n/EHiVZjefQmoNLaLg7dimrrp
auXTyFQwOcVVeVh2d2FjxYXa1i6IP7AJ4+D/Hro8nJqqmSdgHk51MJ8uo56JFbxD
84TAYZ6yGTe8LYBOBbM834H94RYcVlyiljNiFoftadNscVdX3Bk/aBmuX9ZDVNwj
sN0iCoFiZ/vgoCXOoNOYUlCGK/B7eujkpOL2Kju8p85Z9Gk2aBvk/V4NHDNJfXoP
5dxTtyQEmPalD9c+cIxiviIOxK8beePsQk7fD97BNeIO9wNB36cu/asPuzqPUfIL
EtZvUr5i8dcCXkI7FVZZ85VSJziZc5ry3MFgspnCO53Zq5a/2t1kZXRAiIgFHlle
7cPGBxK7S6KbFOvCtlx2iUETRjC+ba9QVjkuX+mfatLPrCOcRPAohmHDiGeRupFa
vynqGFk5ZDlQgQSeq60lILEqKoq3SIKNcCMUspn0dNXoci9p3m009REGUharDN8Z
Fs17Y9Olxyud4Y5Ng8AwK/jfv0zI7wEky1blp3ZBJ8+Jg+b3u/7N5/Fx4OMi4yZc
7n+Ht69Eqi6R447qBK4KtVDCuiAuMTUkJD/F55QCRDIiIOROZ1Hx1GJgGq4WNHO1
BkjN1kBK1wYXa56ErTVVF4cJcaZEUURIn6EL1619ILFFmf4QCb8znOKkNO/WMZg1
PgpFiPA/fRe767H6J1k1ZUquje2G0Vu+b7uMUeQnN6E/aeqCbWvY6/4saMEK8TRt
6/azfoOOpxw8PwGL1Ff9D+5jGbLo8HXBYqduPBfx4/FRbeXsxC/cNqepnvchRe/g
VeGndJfNwQe9bofC2v7WXV1TKzKMJzEblOpXmnjU7g1RZWu0n3zyD+HvD3wMCoA0
vUH9p7AakGLK8Zkp2CstOLFPdgU57cZ939BJxpj+rtN+5HdqCzg6a1AfEi/7VI1X
AQ1ioBacbUCuifUrRUu7NwyQV2kb4qruf7EPE+AIpyE0vHvl7cpRBGQfe3G2Hv+a
eFoUVpTs1pvXZtDNv6OQAqPas0sLStZP+piMSaO/aYGpsG6uO7hKrksfxsGlMQIr
W6Ve+Q14tlBjdQxRlYgO5PO3ecUGHyB4EOhxcrlnySJ4h7+W2Qh81JntM2+Q12x7
xCk/aWwvQf67A+PjAQUXNqs4XtZMBYwRg4oCXyus/8IEmHnXl6ne4sGeSmy55YdZ
N4m9nG7GJIrchhpGZ+OsUFEfxL+vw5KTur9e459FTgipuujW+qSeK3xt8Fk3LLMC
AM8NdSOXagqZS8/tAWl0vrQrQGC34EbKQHv5r7Vwd4LtyC1p5zVUFSStopL2cSP6
9IrFQw3+NtTYI00nXk7Tpm5V+yya3FgECK3d5a0h+CvQ4uDarplsaX2w670+iLOH
wzWnE6AIThe7icqmSHf3rZcMF81uhmKwHh1kPvp4Std424OVbVkgmcQevn/KNX38
wNJB+avEJc0Ipnpv8JYaIJbBf979DL5cCNjGuicNtgAtySj/QCIzzsOv7mvmIdCz
zhqt+2eXaXQtnNIorZxukCmbnmd+1fSFofsVeHexDBWNw/Zw/O7AUUTD7bq+AE8T
3DXGkEQZ169ZyTfCCHvUFyBBaN/XZ572JNHGhWRJS14eJQ4UkRppWD4NkuML9Ajg
BmQ1w+jZ+LnqWejpwlSy09rM1u19rBGAYNPpAz7kq5RaS0k6d2yg677CbhuKvu0O
jFPHMjyUFTMEpsBhuRrHpiPSl/PZykeFziqztmZTGVpPnmO2+bjNyEjbhDgDpVIm
972r8+SOsDh2BO6xdit2yBLF09Y2XYakQg4DqViWWZuQMFzUzYAUaUvKFMtL5RGx
a4d5YgtLcI4CwhU8JwgRV92eX3NsVyK01yMjZsH9B9BFE2iXkE9/6gDycaeG1V95
GiqZ4TpzayXTioamYujnS6Z+0cjdHqICE5n5TWZqFtuAM7nZfGu5Y0yU/hk1S5Qc
qnBlHUxhUQRBODxg3xVZ3CblV88oX2M883RW4qbz+84o+o9/oJk04LbMnEdAtRcQ
q/KmPk+iSxziw8SAIKjIz/A3RdOnqjY4F6sBE9730lCJ8k4DFoDm4Gc048uADZfi
m3xUGRyX3CsUPR0Gepb8uv1Ct6kfweQVmKEZIxuK+sD5uV1z3ava11g865Y9+LKK
8sdDMSuQfG3M+0uNXTq2Ongp5zSqEqtN1ztg5/Sa0fsfmnnh2BUvakTLy+p8rz80
RAxg+Wz6FhdXK21+Iw86C+0gMCE9JLxGNRZwDruLQrE7yoSkG4W8u7QiGEnXLwlO
+6p6GdSrmr3uP1wmtf9ZwhirgM//LyEaVKfzfRhIEovfZzjSHpfQP5RPFknLmWvz
57qQzli24oBPkf9yvh313U7GR9qh1QFEpYUD8jJhjKjxYhybogFsSxhdiCSBWHxY
UCSSblkGY4/VbkqWj82W0wByvKjpd74BGPXsC+rOqUp04Vvx7Fvsgh5G5+CTvVDx
pyLPgR5ZmfcrobYpHyyUaV0LOxA8mFTW+bsQquEhv7tTGkDXIFjqnWuwi1jilwnj
mgfso5mym+ESqL0/YJ40h5yqxlnshsOmuDo3fhWoDBnA4pSypQZMNdBkJnAJfr52
XsnyDqhgbhypI5zfxol1IvUT1LOlLcU6RYlfzn0Y8QpobJqchBGkAJU8O7pXq9w2
OgLVMpWPKDXjjotGs/pQOlBRjZtS2AIxElSpXsR0kUmhDIILLMLUi3WrAPzCam/G
qWW5MT7CjNEuWZDtr1d4T2nsvxYZ9IV6IulDwYZndTeinuBuAuWqjVUtLzzZht1d
CghhV4C7wdYCIDRAXjAEI+q4zEPkx/8yksut9KD0t2nCXBMShq17UjlMMeFd+MCV
KG2yjxpUE/tXY+Ut0aBpPzL/ZuL7Rj35m37V9Ef18cKVx8E7LEtSmiBvUGFWmjXb
gAvaa0uzJPx+jqjCFEIv1arSlw5vaSjczWp7jKOpFbPCP3Pf9nMCRpgFxRsvS/XF
loHpKHujd9nMFn77oiGDYcTTtgnkCB0xAx30QZxBesnw4VTNbraUpDcCMEWKR/kE
VNCxHYXrvGNydyaBiIzyUn2MQlxMTA8JAHA1r1hDf9uOuH7Gcn2YlAdccelM4KXJ
dMEC5PkjjFzvCVKWchzkJ06WBcBgEv8cLXjUPktQ49kF6XaYg7GPRl0gvHyNhhiC
GYGn4+R8iRo3mAdt6WpssHn95iqPxDszGNCSIH6Q2AKACZvsgXwWrNkoPx7DY7Dr
AK3T7IsVJGETF8pgLejlZPGD0Ep2wgfz+FIItdwzbmfKO0DE3482MCA7QqSOcq77
17d8VkC6x7vBYqLEr9rRWcKY7HTurMxvgufrf4QXn6gc0SchCIzKESeyL7zzY/jL
NgOb4asGSHqtpN/a7hKuAXHB+Zpb4uVHUPxYILmHxoNN8RLqODCDDu9b2bDR790Y
Y0DAXf4c7rt0YQGlwUMlpobPcYUFUrF6asoR5jCrtwzpihMZt+VMeMAd44T99RXb
s/u9owL+3IlKqeH4xfGDF7x9JnOBLAuXb+ipeh8SQwyEJ2/0txSs0XFhI+KmG7uN
Hp2n1k07F4lseodnE25EjIudyKW+g9LtNyehedbIPAkH5cvHCBJwC86axR8i3oc7
Rf2b6kIK1PNKAr2fkAnNvv6FgbJia1OmEb9NVGKZuTIEnhqopzYqm4V0C2hMp9Jk
7/hMsEQJxy0w4oFUQmWb3HDEafOAxX2xTwbR4JJg3kfjlA0Z9jGf9ayBDPnIdZ1r
gm2hOkvPtYJJXnwvgTa7u+Oo8Dn7Ty0TKOOVK7kX+QcZoBevwMX0Zd3kt3f5WGyj
SZuv97o/GM/gmgo1dkdBaySd801z2+ifljr9/aCr6apvXQ0Xy/EVBHkmDN2QQ/cG
R6nNilcaIZVFhsokYDtSq5/yjKI7jvBBl7Tg+j9SNWyP0xd6XLSj8GayisN6s4Sf
FsmjyPnJl1ljA1p7ath2oXmp8d36hXBc1uiBBCvAM5+SdIjao2SNXU3S9lwPQ2+u
BuzU+KWDfxVPP+ib1OQ9Ov54Ebphkl6SiUmb6F4dvwKAQ1i4Uevkm2YuSKun8XHY
/BcPBnKbOGC0Vl1sFM7002ncfBp3jx9Bzk+RpkXVVDes2KPtOH90vHguzlRCkLCR
sDQ7YCVZk4R62C0Y/6LpVsZyvBHcZkaNjZMMI7Un8lGJ3O8Gxa8l6mRdJqv37o/a
pC5gNvCq0VhZcybaM20KWGmtg8s0/Srl1awSGqRdSmIvm3R7CuBACqh3HRg8jgNu
vyddq6cMFLqhY/NOBlS1eAqIuvHFV92W8sBO40K+YlNZvOj8+EJ0t1zWyeoVNlzl
rHCaP2y1GM8yys/b+eBtjYlvjnNLNEX9cp38iFt1N9GAzcOXgdTeEBCBaFXIi97N
J5lk9C+ksHYCfNYNS+W1sNqvd6/MewOHZzdo+gaXg+eZFCLWeggx5DuH1oEk7oZ3
dZcr8je2c8b4+DhICdPB7giHehpu4+MJejj1AWMct8uy0t1Wx1gv64PKChk7GKdo
p/yRmgMQxUNdBIy0gn+K+7akGUmON2CmpY7o2qCGP3oZhiVawyuNul0RcBXfeG0q
eMW50f8fnXWR28RXnT/JDz0HMdUXBrwEyHq/GCHi6OFcOdVXJovB4VdVpaJgU8eB
ajykfNMbIqIZbVgAJgDxui1KLdCleubbnq24LF5xFAnc91lBgkEby4xio5C9MAu3
9doYXGMR7F5DlwflgjTcTo3VlmPKIaIfZOaHFMnrGOpXD/sheGdLLUbf6Gyhx+51
s7mqKa8hfqHduS+d3yq5IFA7T/enx36rV2Ps0YuzceJb9iNAAHSogdx9ydWA0D3A
Zp66U05D742zEP+Tk+k4I5EO6cMR5N+CRa90uRKf2hzKPjlxbBCNmzK8tHTR98xH
55f/Ca4t/XP6Beov/Zh6LWFCq5G7w+Ia/LcwjPbTK91spIDYGOVPUhoasNqIB4Te
E+DzVDp7oXo0V+KFEMDJIvW+w/0+iE+cOc2yptn7b0bPUSjLhqsizSA7VK+Mkm4v
dy+HDJBnwvKB0Ys6Q8YDv2vQTlHkSfZ3g04xqGye/lANYDypmGEK9o+KIZRjVigo
i9kKJF86VbBv+q629cJTd9WUGSL2JWOZbBoPinpf6pw0631w6pYjRpeM+ta++Xgy
cmwhC3oQwVY5vps1KFx63ubFwPiGjHfbGDWAVotj9+j1+Mm+klt3XsoRw+z70P6X
D2b3gJHS7MV/ISPjyTwJhIQcdgP1+w16PBNz6X8FcwjELJb7F9+nOGINRkyA9t2x
gLO358zRsFbXzUZupTrgc9+8gvmqmsWfEdztQYAsLv3QfFyUYi843ZC/eJogEFsY
41xm0V3Iey9DgqZ09GRMQqBSTR5RoD5/H/mR8ddWhXEs1FVQn9P+gx0inZrIKk5I
RRsNz9gHSk6DBDA0ewzTTLZHTlDs9a921xEpyIJ3wN5YteQrns9WdwUa2Ah+1gLH
HZZE6Ers0LW2PO1GKA5/UeTVVvfpRstxtd8sy/XnM7N6DzLM5LGOIbfsuu6cKLcQ
To7qHX7XquRSMumNgglvoV5YH8KQJc6SYFDCUEfpB2leFuCd0Rn7PDBoc1lvGAD/
LDvqncSdwZhge9eJomhhanzL7oO5wE16EMhFysAd962iYmVVsK7V8VjX7O8FOQYL
Mta3DWsW+Axh0WQVTaRTXjR1e8U4lvSKh0sak/WfEN4fZh097xl93/swYZk5NxS+
llqJHhZoCfxMeucqmN7fd13+xUK2ZvFw/lciozLJO/bXaHoV2v1922XHNcmVwJ97
o+nVUYQH0UvLTbjeUlEKTBdUqg/MAEV29W5QDgeGuhYGXLuU5S9J9uvW8Jnp5U+P
UeNVHEhZVLwq5o8ts2TCdDFuGV8TMpEsSQ8BPmEbDi6hrVZrWN3z6Gz7uz548vKQ
iidwsoK23C+tWWDivk3p8GDeJAMYb6VYj8kGMgKFUGkB3yEkJE5Oyo0NIB8Fte2/
3w31unrXqlyWsZJwcQiyDR2/xC4ll+8YBhdVjc8aHD+YYJctGSYz2ja041epI6jT
3u57q7A+XND0RiIGlJ7qLiWL85MmLL41dkNhrqniNjqRI8D54kXjYwtUHKVgl7Ku
gXwt2Y82NifgrID7c5V8LQd3o8J7Og0w9uEnb05FnEkCOESWHn9/THMR6jSxNZz+
DGPVQSNKe3MYprxlY+88ejPPc7CJmV/60c1BCyHbCTYELMgyweynV6A15A8+bz28
gw/IBrPXmbooS68OcaC/uN11ycH/+P3hKKHDFcSFCBqWjEexofhAZQo8me6z8nQZ
hFKiCTosSJMvy9xe5kzqxehhAK4x/ADXEOQTtH43obApDcfpaKciV2//USSxir1H
jjYDvZTvPctisCT0DwQPzWNpLl0PMHjVtNq68dJ0p7ULHeOBLHNzoPZESI6sL3hy
68OJMG7CXVaA1BJfmoh6A9C56uJtpO+8in1JE+BPkGQaYJDOkglhgJLQB6DporpP
HCrl9iuBXbri+/IYgSLqnnI03BIssGYSLRtSoTvAcLvT3kkOkZOC2Se8EPszQpj5
AjKbX/hrwHuIkvWX1IWYgS7fmaP2lfcjs4TMG+GSFA6ZfaovMQkLojjGyx68r+X8
aJxG5JNqGhPUGnMzhes4/naePMJYmUtgL1Z8p518WY6DNfR2S9NWPMNn98YzcNjM
4Qy4oBhG20y+BeIiqf9xMMP6Bo5sAgXDzMYRD6bzrHHatd+wON34x8Zghb6XcgrE
9sQRBKDgLk7knwsVOTT6GnyWp0qsbNmMXIe0nDrj6F1WNp4ldrQoo0q4Sfn1rmAh
TDMmxT5XRivnNR5QEjp3xz3rJ9XmTIk/6PWUmrnQJgPk6BwM622m1n0+/mQsuySb
NP3nDY5kjGHMJh0aRQCf3WXgOkZ9yjkZg6Uipyj5oazCg6CAfWPoZMIsYnCmgsHz
CC4X1/FFZVOTcUEHEFOhN7+eowagD+dDJe1zFDx1tOeYSv1d2HcFBlE10cBPunch
2IWRtr3qsuSB3SVaV/tNzFIEksJHt7NM/fCP/r/lnFIoQtAcdgSAHhbDXCESeYEV
EjkBQU6xmyQuoNmpLzIiHNMsmnan0qFrsfpiOX0w9kbpoY1Cx0f70HyKF108nPgX
9bIoAnTloBsbumahkj4jFcqxTVyBleH+cp/LYRaNHYSOsLGj88QK1tm9YpU/0aAO
IoedXomzCXwi4VrNbcSJRkihPbse59QAP/JfDb+qFPZYqbYwQu70vZLHz6KAdzpP
Hezersgq+ny4mpLjcZ6juYtS5hgrVXbre5xQXUPznwRpguK1BhlbwWU3tMcCQvHa
KoWDT61aPRZXFsJv0aKu2PP111KdyJsvxnDRXt6WxAoCqZ2Qp73sR6cY4JQPYFdF
xN9QViSbHJkv7J68yI2W70MOPuEvPimzn58wCbbDCY2cKKQJQ8GPMpq1vdlbehSK
5gfFSeEEiwSgB/Nsv+Qju5qBh9WN0seLrHZ0LjSfBhm60zdMj6KmPW83frqfFHvI
nu3Kg04oG2SSPEpaK8tecyf7pmfReUO0iehg8K9Vi9hQw5U2+sVMrevrTqcV7VD0
x37PdrInu8aINjrMNUR+f89QC+LG7EoxV0Djm6gt7eCXbMiMQqIleZmTHBuqJYDx
zrG87QicV7Ae9+VgVqlgXATs+TNpVUqn4SyEzYFDw8hBup0zQaK5hiPNqrW9BVE7
yYDScXWBgpSfHoNJQ2gk2x84F+9aos4wj3aIHsmKZ2RkQgjLGsXWB6AFm6wKAIQZ
eoRS8OvWof3UBs89NWcN8w7IvwMlbjqWboBm3FKP6sV126WlsUUeOP+OgqbQYpQH
xj3BPTg37Y8xuYO48Oan/X85VkzJe8ThxdA+1zKWQOvZOnFSavheXUoL9ppBtWy+
FrpSTj+ZaEKCgMA6H52znR3Zuj1F5ZRSOa7FWMG0rbM0N8JEyu/3rPd1USvyzhmQ
e+BvH0iBf5RI8xwIOcLABSpSQFpF8aRC+8bHMUhYu5Nn4AV2T1hCQi5J6TIRQYm4
pYUaaKdtUoDgW7OT4eR9i8H+tKLBn3220RwdDzN73rrEzqI1WATAZpHlJU9z1xht
V3vbl5vODEKixxn5sX1pnSi1AwAXj7lGnqVuAXcieMmNrxuoD+376NsuB66lff+/
pUhJdZCUxu0o18xdyd2FlHsYPXtAyErVhKu45GJORLVt0NmsnhEXzdQCyyYmqHC5
N58R/agxWQFFwvPGTMJlq3HYJJUVOCtOUWVSyn6vAOo4MbWp5wu/tTgJRigmOeAP
sOieQSDI82k2q2BG2RfBf63nY+BA41xtd+oQb+Kk//OWkVzm9whOrAiM/HEjQMTn
5SOdPkqFeoPPtEqkKTJHSNGEMQF2YOpfeKEAk4gvTY8qJ3/jYLIMhW3D2UTtqHn8
G7iLRucpPciK8faYas9NI2ISHCibWI3kYnfr1s6r92KIkj0ROO05Of+ORe9eDHRp
dAI0oPCH1wDpP5qT7OR17sMcwv5Y+tObEnt5s36kCQyFjtT5yt6LVAmOveDiXcRN
ASRCgCOoNZLMtvEmEqZlP2MmJOGhZjlj8usvhvCQduvdBQRhxcUd2+vi7iCiinz5
ChJ+moWPbLK0P/pLIbo/371A0BZ9B8FqoJmhuKGRgkSUySIVL5a9KDJnG5NRKTjU
9pCc0PGsmld+HRJYXGSfTfIn1MSX76eqwdvIeqLgK4nmMK9MyQWudDegVW2SWg7k
BbsJSGdXIROghFBrnI3xUMn8CrWEnWHJO2hCV1YWhLNx5l2nOVwP2rqe47QhL28r
L0E+nqTZuM45t9gjeWFprQHXGDpTa3e5XjxeMLtlKNI2MUSY6FLpjhZJtR9JkdoO
imj9j/XfqMKCAxKPAqhem86ANZnU8ugfn1hn5E5nENHQhTsfaHTvHU+7WznyueTU
00aPaO+ggKnMrMgAAWPEct7TUnVwUhY6EeNqA49vKuTlioinLvkR6ihn83sJ01ll
iRLq/Rh1ltR4VHNANytqIPz5VRxjynCO9gtBcUrr3Res1eSHRZePMirEs1s8xyGP
xZleBeUEONwW9UCdagxcyokOagVfqRdI4Yv3v6GoWbN2c2ttyDmFptmACkAYaV40
qS/hmLeDNQ2HkFaQEp6N+YVkXEoDKE2Xa3fWSk9vzFjWg+3qhTCtdWFrroeWrrYC
E2KPJYumNgVOGhCaQee+EsJ0D1BqiOB4A2cLNqs0dL9MisrlZ8gt2HrtGcKkmOaX
J619e+XnxFRQq1prc0z4sm72e+EjCJFXbPMqoi1Sm/38hwEqggc29/aM+d+QFq77
+Bpuy8OE11hm/2pYqBQoPWb2qCM0d6pwMGKlj10b7ceakO64AS2n/R1rYUyt0B/M
cUcYBVpi9Bf4+n8nYdS0Gia6IhRUD8QrHvYquwX20aU5Lr9sdEnG4muLx4C5uoxx
m9tP2gBtfJPe0oU+MiwY69ef/AWUz/hlP+XE5MTI1fL5PbRGqcLbHn6DprauSa93
pGxyHJdAf9Ms0W3JwtPXMRa/hle2Xc+QWuqVr51rfqF51xMcd7eJ7VZqzFJxZYc9
8SqD/YKf7sicjmNcpkTdOHKnH2ovkcZGEJ8Oe15fiRqfJkdbOmzjdQqO3AUBKGtq
A7MtACT/zwVM4NECW1ffa78vN7xoAFfBDROdhL0S5B5HFPwrgPEYPGTtLaRAaNp2
vicvrMYek76Ns+7HeHlq1beCMyhweShz+yzgwL3yrL0T0y1QLhFdQ+ZrNRhuoz8O
kYR/X4RyblonRZdd6P5279OPuYOn3NYOyxRQa4EhOyBos6+LJw2AjCtWCAf2+o7U
24rsiyb67EN8JAZ9+l8FVQNoGhFq5Wl3oUeYjwVgAcodrnrTnANbuolh7jCKy877
77edV0LR0ldkwHPw6TTlDg0ZV3OUfmPNtCSEn16fvSaK/dKZGBxEHXOiNMT8JUwO
7CBih4fqCX9JEsUZdPNy4CHOKJZ0YTgznm493HZ4Oxx06nAwV9bQTQWS5Jecj78Q
4yNu79p4iqPvUiXZxtUG3VZVs6cYRHof5oEtR8bsEUlID9zizc7jgOl0xkKV6LYq
Oa7rSoNlEmAt4zwUPcKm3Sgk4AZbEzf6hXc1u3BDhVpSbm3rdhWKfqE8u1YrCvp3
MrxOnjawsvtfuZidOAIujsGhpTL06bt+HIobpOQJ+haJZb899gy4YLiZS7IJ8Jkv
8sA3t6b9srtwYiakYVHK1b2JsdwChzN0w08rdHAhQC1U+Yrbe3HFO/fdE+vsZA7m
t3EDIab6+U4sN9Ac28BKnB3IX6oTtgYRb6KSNaFUzdO1KounnPYasJjsKwu5UbME
Yypc1K3q8esAcoU5swDIWoxPrTTaYI9KZ8NUbRmlR3E38c6NbMcJ06hcJvnXgLsb
1IsL3vp84mCNHY0U3Ns6uhQpbEPu4l34HoL924/ylRAWibtXwDboEz6bdDY/tmbH
vBWJG+6dyOxvodL/vWbrbhsM8VCBiGZrfwvNJoYxtf2rRXDKqg8BpZWupfEmGS5V
1JHqJvGFrllFWPIH11gm/1vQIAQ60wq6fWlNAB+04Bwv21gtMWPPW8mQUNVydWng
bpLc5v/h3t4y9/g8IpOgj3w61juG6sPdKNkIqikjWIXMuC1z1N/tSrSwNSlaqYTR
mE0siOpCLOaBMp+5nnjpPsbIW7ifsh6Q81IPtUElP1BZOzk6IA7LUkJSUQFRwjHp
576vGrYcFKYoxvmk71MejqAPFDfEAHxnsI71dG7bRRMgX74kdy/90+3oDhOcNcfD
LpEeWWIEikqb7H2Bns3tK8c3ceyYXwfpQgKi65RMCXPV8XcS/UcgZo4C6gtd9TfU
kbJpYhWNBSqwvTG0PoN95qjRQ+FDTSWzGtcs7Iw2VTTAZO4W2p6k6f9cSK1C6r3C
Zl97vuUxr4wWfhEizCaQCVW+upUokfvQ8iaUe3a5Rmrph+xoVSsj1kcp7Enrijzg
t8nEJu4ZoOCeAeglJSvj6SK1I+OM07MUbEFsdqN5TvOFaBHh9jUIgNzRBjt9reOX
jOhM3kbEUR4jhgm0MGhxRxGiRz3GRdNt7XispsoeBDrPIh97fgvp6RCiqX42N4gu
esdaaKExR+WUrew2ANuzMv0eVCeBPvqsOKpafKrFSEDKolv88heh21PdEYLf+x5t
Y5iu80yZfLX+SrnJikCFyel7tQ1oHTD4LdpsD7Lhy/CAB1HW5Ux1ragbjhEKgir4
UdlgW2P357pBXMHNL0fbdiPMK2spm0xnOUji+msFIJxRZJiby+4sp2w1/k5UJwi3
jlCrrdSic80/MFKYGRKYbo1JbAE3E9q6NJYNPTR3hoGq7fkxnOzfLeZLorEfp9si
y8O467s4eVXmwNX1sDP238x/L+Yu2AfHEKpX3jjCrHuBYXtVrD6Pk90N2t0ROxbO
h83ifY6uT4fX9aNWLh7Gr5wyrUKVFLs0YaCe1qTuBmXCZI9jO3yt0iysWwddBDhE
VNX2oCjzATqmVTJFXoZT0IRw1S7Xo3MaxEn1N3j7fQLnpo6noIj24hyCO8dV0Cu5
eB/yzkHtZjNlBKkj6gmcDfCtsmorwnSZc3kShitsxrvOX1wZhiIuaPyS6wL0uMEP
EvFBt8xr8bFypu9/UZWMTPao7yG1r7vyAZ1VbRNFQRC+D5Aa6pJVVJ2oN4+mrRat
SOzeJa2x7MdMBVvVTiA/iwhOy82G6e7ijelKlFNcO5iawCQZjEkvoEd/qxES+5Wz
h9RS33DLrTy9u+hgPdE5FHBjOkzMO9V8B7OEmwDd22QfWfjH9xezkCHufi1rKFf1
N64w3EmxTR0X8hVXTJUeaBxeHJPcTCHDuWpDMqgSm8s8Tp1N7ewE7v5G4txy5kMq
TwYXb6IIXpUBWJK2ymHY4BGlWw6ykcIyQO6lA08kCEQ6CJsVCutLDXgPqaDQxM79
YOJh6MOr6zZeTJ4sCeTxoeYa0LfVYYYpIF1aNEVqOI5xozbNThtZ/eNKHfOjHXaC
vNkMmboXuauIJHv5tpAnevU04AVM2LD5Ms/21h7amNwQcd34/xj2vVsiBo2cagPQ
Lw4qhiOuq8UaKnHpxtfgawoK+q3NuSGSbTC3aWW2Asm9uSM8paGvwwgdcEWC+48B
lkWtk5qauiUuu2IR0Y+c1P01sCL5EO8NRqr9culMwFWcPvKQVSXV/TRxvBw9kfrg
hlfEn86yYwIuqcC2z97dX5esuJe+KH6SGowF3oTve3qhXLOUX+h6j1cbbWRZSwdd
Rq+gFOSmo9sbeixYs1YRM+L7yP8P3jei5p+x/5Owu2WgOryaaf3wsoCCuCCPSBIw
LSEN2dQXN9VNhiVAVrDqLKQaW84ccjKSQgHO7WnQOtajq23x1NJTQ645hc/V67gY
htKVCQcjUGfn5GoDLbOgbZ80AO6H92D+iU7UxPBdDZl9VwQcs9ZBlqfnLDbuVAWz
EfzROEeINa2V23JfhktZrATdooqnbhJQZg4qrl9JE28jmk0UeScnVZuNklTimgWy
KC6EtVXMdfDEDKHwZbInUhBYAXn5Bh87e4Hn8Y5Y/yCEa6Zcki9TgagLp6FsFTrh
U3IkQ7t/UITMlYLht9vLsKkRX4dzuEjJqTUiiovHV47fRuSuiBh94guup+UFTqAf
AFPLahWgQFB59STJ4hNmvZ2HpHQ84SnfQIl1lmkRs7rWYX+n8+MGYYLyFD+s0uGT
bqAXHtbUDuJsol1o3FbgSS+B06XM/VhZufsunKOvFf9mcrJkSkq7oI5SYC2cj9Bw
t1jCigJV1aFbg4cFf6kUwJEZlv47PZzIoF71UtlyNAeKBakCg/ysdxViKcw1Aei5
4MrjAGG4X/8aQ5luzzx2OwEb8SIThjn7qH83/xnJdsL7WS/QLBctIB4dfAJcxBKq
ByaS9kRbNFnQBsMLOMd9sLIDXl4A1/ObvnM7CD11JukIyJuatQPvx0bSmim2NwPT
sPX/e+4rq5sDaN5N0inc/I7aj6oV7+3Lg3xnJ4RJkFFyw93lY46dfQRrTWEU0/I0
VREUukOOuVHyNuJdGTV+yKEa/ikDa/rMK46mPGPDArf3bHMB4Pc8Drzbvm7N5SF3
alDdJOPSKE3W80BQEHWyjFa0i6EZwOlCzZTSe2uNvTcPJt3IEfotC7+nmVm/6PEZ
qjS+OUrVWVHYLDDVaHZgUZ2kZbTj/b2NCAJWThD1SWkug7qcUq3g2b0kWaaC5irv
oAb3oMwY0ubL9mLL0P3Szh+VLnZeICIh90HkU3rYPrgIyUyUwvT/G46qvg4M50JD
YWzJrAZQj4JmpE55dNGv0LSj/DtdKmUfLGTbTXhc0A1N9sfAx79B1tTuttbcPx72
F6TPRYJ4oTu7ysrUf/5/Qy9PExYWFhNbJAJBFM4zcwuNakliJq0uizIUODsiEcWO
oRvXcUSSdcXji3rNnvZxF5yJDx5l7noyTs3ZOHlgM62Fg3vLeE2HqMTdAlpfOq/S
dggW7paeq7ZKZTtg0PaBiS3GTZsB9mB/f0n/upcTjdccucVAyXiuk0IUZ5EVKbcG
HIRiyHj9KO1LIDnDIn+vyHyTyYK353MTsUN4w0K+FVkjXDN4ECZVALhvCrhdEm/s
FhRQGNc6nr+Zie0MBruvdQdIByN79tCB8vK0+thGvMZtfIBYYlNaNxoaw6cU1Q6S
dvZiknoB53z4rhhVU1uR/8ZfIjzPJiCc21B2HtO1uOdX5MmWt5gZZnK4O1mwYEJP
/v5rZguS6h1zTP40RRszQ4Z7YEoFXTSYeAFO70Vzdxd8fOp6xWfU2LNQ2hkHHBS2
BI1I4LGHB4qqa+qlX9I86XE//Sw81DzNGBo2FQURHtSdbhsVGgqGba2pEKOLsIL4
uYuoiApd3MKC4Kvia6ILNgajC8NP+5vurfgf5tL05cvk6EakNiBElP3BkMYmisLW
r5YIXcwED9YLnCKoyIMhvXldKUwhODNWzWcwRDEFmdIMjKuMljHTWDRjJbv2WhA6
+SFBh02BbF94IpFXucIbP06q7bzv2fCwzuUNLMdYderHrdriHIoG28SN3p7HXe/C
/CtLm5b2HtQSWo920siWvqigRbEStDRieVQuISMU5GWR3wP+u15f1WqljovFkHgm
xnTSiYK2Rl9J6/s3aZWBVbmDgbiM/iaKhOzBbDaKngkxRkYMUMS2WCgfv1nKzdbh
FLkc+M6Wo2p1Jo24DbVVBQsKoj4YVX5pEaUdFDQ0xjGbwi0QYLHYEYMPdq8Ow1i3
dXcMWSr5TK5K3uQ5H9gCfX5Pper0gGhRjMM8mTYR1n57UbaeRzMX345bzZEOO1eE
zhPRIu/w5I0DurZ/n8mX4Q5WYgIpdrfzZPhN6/OW/3GumibLTRDKduqthlX1K0Mn
yxr9yOcJ7sV1pZ+pZjmJKZwURvmyvpjCV0yoHwimi9Q9wPhrbccFda34iBU+4Oe1
yZolLz2EUlK7ZFctzuXzPIQdpteJ9GIq4Wu1p6JQ7omQkq64x1Yhx1xXiEIB5NxB
Z2sSB0mD7CUrQbvKKLxncipq/MErsBKJAdqVWot4KQWvLMjefK0XwcilqAk6EK4g
xyljLt5aSzmUzKu8fXg/IvQNAvGOvL+O5JEusr7RcDB+QXKy0j1my37ytvIGdNnf
f73Nk8dmnQzmbiYZQ/WUAg7vDdfb4zQNDS7qkTYvAbliCdgbzatu0DE3Shm29p2n
3cpbYVHqiTs2AUdUekJvW0FKYViUPcdk9xYdVCi5UXrWmj6M7tFUqaQU0LQvma8b
Fn0ZtGwaarQpobaXvpDtf2+9a7k6Nd4Jrn4O8Bt7dIawsLfC8kdwhB4VvYn8SB/F
JnDM/su0bnHyXs6EqLgJHsTHsdgGBQOuQJYzDbz4+1sLySSk6MtcssU7i59on6Gp
wLIKqKWjp0KqrrIXLBU7t0YKdH84kWX8dxRjvJjrGoERKwM+VvMlQkD8u6CJuHMm
/bOiXHlSMXoObuWhpmXIsjtDxdqvuxmFL1kVHsRMUFfk140DBmb7Ib7iGVYEdEkB
9z2EunFUp8ZWLYaCMJN1B089PnSNvWX2GyEli46hSVSCrq6ZyGpjSM2ewho7GyB7
i3OTUcqi/58Xh7UlYEyvekl9z9i+ls4n+AMYk9bNyeDkokBXtd8Fh4s9hAgVFeil
uOR8gIEgBLaVDNqEXBBuPxec17guTZzgsKq4iJB4Nt1Se0KvLTaYcPKF7DQCUBe8
V9m3llFgpjlm/MFI2/FR+LPMSTrbAgY1+en1bwMgWvwdf7P/ZOGt7PFwiBxQefMR
NV4Ur6XjiTaTGA0lJUFFSas8KYMDFmwXBPB08c8eUhOKTp+qbQuOAs/XE6STdXvE
83Yr/W786rW8loUAhEs9vw4HZYAWPsRO8b64MKGP6ujWN7Hjk3RA2zjzQbyG3+mV
PQ1y4K1B4T8QWKDxz152TFeXURqaoGNJnsBvxVrN4eUjXOU1WbbfLnY5SHdZ+1Ng
0v5a1A6kGfj8TnQcqWNzb0N0aypXarJLf5xrfEXBIBdBTMmYUkvVvVANROdkdo+L
l/i752/BsCo5j5j5RKkmNpTOhBYbdS9V1ucTl9r7zwXv15buwiC2YrX6Fp7pyoDM
miH9+iqu576/dYTRZ31LAlFlOJENyrRNBv9TvRN9iOZJ142jJoh6D0SdlI64tOit
QuBry0qcRcfE04VJNyAlK0DZBhPzl9WfYkw8fu9YafjM9Il3TuTL83oa53moKUnn
1GjJu3zHHXsy9IpYPfG4O/sMpvDU7+5UdU5z97KjNmvx7bmO7IH8epsXZGm2j6YT
QAqqVef7+FR+hKeeqkLJLMUuG50pHn15OstatSicEFW/xusXW/jeTh1OuO2/XQN9
4aYTlaPxF0aPbL+26Z46WdcSfXmW4eHIKKQt29uAChYw/wVh0bFy/dKDkSkQdnim
siilA5rZt+9umeY9l/8zK5LdW3MLh+QeENms1ek0SPujgYOW4qwE+fjrstFEFn6K
+bBjd24IHtrxOh1mjAc/G2jmOME2QbAH5naOuPoe+SqRiU6WlW/1p0VBVqbiVfBI
QR+kqSkaoY+bngP+B5C12o2H79RLLNWDhPNB6xrISz3Ul50YrepnrzpkcocDn93k
coFJI2skJMh0akiXoJ29dhCMQTD993DvglSg+DBa8OgCGInXgBGDa4E1LZvNgto1
H+P564pJlrE5Q2BHCcTEX1YjZ2rcdwlQIoRjis7UQOpUkmSZjJnB1FxCUcVYZdni
4Lf61HZ2x3qcOeDi2c6mrUsccQtJhRz+BJv9rdOiwLEhaLv//0p+gFbIwndO/PiD
05Z35n+XCTN6Z/Wgxikn5syT3hJzSjlVEBTFgqRxyOciUr/hQh0SeyAhxmWAi+Od
EzvOcugDTc0NeU4bokXzpJNH+M+OKpbCHbcgj2v49liXmCypn1pPJaBb+Hk/O+M1
VRSZIytlfs2aByjSLrLITzupRFWitLaZ1t4q2mqVZLGXfmvJveX13Kf/gQU6wKQQ
mVrGg9a7bXE+v1uCD4ixudAAR/w9qJKz+l3M2IIAvsq55pW2PcANaZzs8sFu34w3
XnTTYg2jgFQNOV00PqMFaoLIIiXDplE3fgZjEMcuthx4HMWmQ4hiQT42VKGruXUN
YqGElIvT/b4A2ubR0r8jUhdmMKubUQxSB4befGtkBbk+ZBooviiiyMyIw3IO70lz
Fk6I78p/alFRg5LDw4RC5resEN7JmBOTTKqQYWwPBZjqJF6hyVvjTMI4H3nXN/4i
XIUBjKfW/maM+Az+2NOtl8xO2wcPzg79R0Y4Vvx4sz8I8CbBPU6G1pTqM0oYoRRd
e4mHdZHooSOYUVPrMDye1EiX/IizLOXdR2qQcshCmw+42tApkZUMLv7bspJLgnce
3opFqhiLJXKGy0kEqiVrDFY6dW1MKKBBMp/dImLANkD4IV47wO50HEZ8RChME3ea
Y6KX9q9FxYwf7a2GyuBkz7QzeEq85WqKTXPltmcydFqLCKWUw6ptp6j6bPGaZUnj
ZT3DpMpHiecnxzfnMI6IAtw/rXB7ZhekE4e/KtjoIAV0z86o4OP47A+ABLDFQC+U
F3Z65jOzynjGhWHA5E+vWi1IqrQ548h9XynBWN5rQ5a9nXH6ySzjqsahmAtgvAjK
2o2SzbBe2oWzY3FTtIxg602iinwwIMFXdtwXv/zUgkZL0LWe99bNCaUK5aMhdxoS
RZlrciedZpKmJ7KlKdFJa7K2eArgE0E6lbeWITGvyPRtPBx8c7smnogexp7yJ1Xl
AJnUovhw82EiLBzcwlYmS5sPiv6lUfnDZx29Pt1u7qMOnt96mLdfPLLvQiF2DEmV
caRfQvrQjma4Lr+um91lTaKBNfX3Hie5NWvB91HWCarV1qOn+nEDR1W8acscmNNP
mHYM1lkifVZOrzujmNUGZVJ/i4x9mAXgYWqL+okUUC3iPNy/xN3eFyyGW6F/E5oR
i0hgrhfQAmUYocQrCCVP+GwQ8IuS4dbQbcGwY8Adm6E45RQyHMGijeJmJJLuTWU3
Esw504R1d/YSJTLTKAdIPBGAyFuB0fbax/GAO7xc2kSWVTH7ScQzvI7q1HH3GChy
IiP/ip/gxz6TZKCiug2qXeGDUGHrpbWY+YdgH6ER4Wbeqfef76nv7UpszSVUmUrH
qfavABBSwikS1Fe/eitlJ2eEvurXrkOoTWpXUvNHYR5RrsN7odfUjLD6ZBjNp102
SjIuB0/TUICd7c5bD073tRRqldljA4Orx8N+ACjYOv9FyBAJ9TnyhPYxTJdaWEac
xpo4qJD4pDGhK3PSa4gxPB9oYUQKd2rUHfTR3L8sFlPXkFzJ67AT3hdDwBANuSlj
i9JgsSkuv+GN5AMQ/LRXGJRHlgZ9Uj4iKgozvvn3p7b4Rs4oua8dzJ8Ztk1FD7Xw
YcdCGL6VaNPb+chOgGp8mQBq29OqpEaDSiHRPBt0tG+wM21+2PKYz8haUVitM9VZ
R+9EHS1Ldl1OpaiX9UcocmHz3IHjlb5mo/f+xMkf9jGFT06n0L0gGISxQbgIcN0I
h8b+19QVtWnD37bwRbjYKcR/nDSeXXdq13NtoVkUjXSpSEIuqG5ZFmGuxtQu3ngh
hUMrmwB4nQ+PGYMFDnDbN7kRriVNSRYwR+brPvA0jRUYz0L9RJaTkX4KQm0XH0a1
dWTzxRgYNA9aCAOv5Hxes5EWM/42xXpSGUVxIGrh+SVI3P9R0cPVv+sDSOHyiEVn
jxsw1+JP29SU6svtwlolTsYrTjNOfXHjEJ7fy0FmPPbqNrul6zznxnACQgi/o2JK
9ChHNywIDMyf1Z1bYuccIA3EEHvyaZJN9S8vVGClN69Eh6PMsbWMo4g1rM4Qr7sJ
FnSxOTdgh6i4/8eYLovAfarrE7U4ZDkg1Hgxof6Ghg4NWFN27HsYPMpAeo45s1G7
f6UAHzUyWzNRzKcSXncji0KHwube9t6jY3QVkM3oYAVhUWh7v4MGExnBpoQU9PgO
cALH/9k8k/1107qzJ+jvqoSAc6XX+mQEJ7tNgHN75v44PjdeecsriGuLGwWzDWtY
WtCzOCdKymCa5PDKutiMrn67rHImZFXaDNhV4nnSxneUHH8laRrJ9b8vCz6wBgEm
njuOTAsoTIlhadXAP30swkbZQtKTk8yZA7Xe5HmUEmFVCx+SeFN1Lonnks18dW1I
z7qfN4T5sKuu96yEyRKO2whKwr1LOR+lF4oDR00kN+xunfu5vni3vLuBjcjVxzhd
Zxj6EF3sBeXaUdMCZZBodwSJVC3I4NxB8XZnJwNHBRoYS/h2llAppbDpYFWrkcih
tR+BFfRjHiTUBIW/5bz6CsvkJgXtvHixOnJS2FSIItM/3iqs/kuTdDmO9elUPtuW
HObq3c+m+pgi9auMIw8IhU9GIkDQSWO3tJftxhOVN44TpV1V6dgiMipXWzfrBWoq
wPPOp8BftTuG9azShGv2VkryJDujP37hSALn565dPU66rU4PZhOxSBgEq3xIMUOE
UycbS0diOvCkHDYvC95vif0oZCCd7exqnIcFpsQnAo2wrIz7LR6LUGYda8Y2cokc
MZanbXI5AxICgQhV/B0HG2Pg73DHO24WXUtc/RDGXnWLXTV2Fx5ECiSuCCAvJyWk
ke6XDOI03fNL+I88fkQ0dU/CzzYI9464KddLce5Va36mKwJl3TDflDAnyhdqi9LW
xtgfvHxuMDBCmk54ywxe8Msy2DeWHUtP3NkxuVQlO3zBJm/sMF5Bp+n6KOnIZiTZ
xvBWYxinWGo0JdVLa9+fn4mKAvnvG/datSWYgsdusvAktgIVuULVZ0JXAN1IbAyC
6iDqzi1DHPqYAGDczK9uSOeNI7Db0P+jDuomBMcUp6uPJPQPgH511eH2BYlAd+9N
juLH6KfYKuV53ElQwoJcsqPre2RDEuwQebELmNPh7uUxo+3LdF03YRatgR/2+ibs
L4m2WDV9Mc/JMD2E0zrN290TtphqY2dnMtuAO8VYT8OXw1mykJob7cyAZ2rX2ThQ
4xHLQ9mx78guWQMmN1KoZwQQdFgAqrbLCQIDvLxhc8svIjDjhEWnfYGkfNeiCMVD
Tmt/Hrs1OHPIZLuVU9mcUxsganIRdMprTrU7KbfxP2OoCds4zuoleDbgSw99NnEp
hHJjYAwVQHIKZDtXtPMd8JEBbgZru1yPYDD9sAtJ0pZQpV93lSdEkvivcdrSSR0K
qFcvp/y922oGSuAnWsfZ+9+dGMHybraFl7N87zu8fgQKl3OZaIz1RvbwTVrZ0PYt
8kqUtpQLzRsqjmowT14gtpHrB0DLSOTf0OwXzL1Q2i23+w8ST4JhX1Fx/DpGv3/S
5QJ9Q1f6q3fAL7Ir0A/UNqPLVGabNTm7ivmnXc1BitHQgUpUUIVBJ2iFubp/fA8/
EZTjCTgZhskVZXyG1mD+KZKuoRsxCuzTwpRN9tOHDPIW2bGRSDMOEu81lzqnVMi8
jfZGZULYTfz4Nh2UNQ+jEmzX5Y4ap2b2ruonFqhAUOLhbJPdgrB0utU1do+L6ETf
2c3Y8dY67AeJgE03nutrTV+TIBJdnNqECpUma/IpCyf3RSRquw1a8CHxDtKL8U01
VuV/whvCsJhSYNZP8XPk1qgIbuWkLcSft2XXfUALkF2om7EKfJac5o+vV8YPrggb
wgleQYwR8z74JqfI30G+lqpIQ2ggMmk+ylyAv3hOvUPKFPQ0LkL2Qak49GhnsdV/
XTqzZNoonbDfKwXMm0mvf5ajRxBIuhTK7WRD3G8AMCPWMc76riTp02kv22N6B56b
icnn47CpEjdGIDralhY5to17Yw86tc8k33jMHDZAXeuEGlTHzyxb6T+JKp+S0NzK
CydRTxDkOzAG1XeoBBzg8nY1P/N1zkFToxTu77mtJYE+OIOStD7OmuM8pXG6IBBK
fE1NlCWqN9w3c/7enGC6MQ+4awgqGN3p2Bvum6ogBmB6rT2xdhFeGkobUPLmrxNw
1udDKiblz+Bge7VU4cMCY4WUoY/2dQzzzEaI6Jd0vTstjspju5pF15K4s++r16jr
sEksNnJ9CXzjBQFe7pp/LqrfKY1rYPvjNQkabp67T2kRx1yf1DNEAe0wGaTKzVpO
NaP/1K4+rU/LfIO4aokPv8ALWie+vpWGzyjkyg4y9+KXSRnxW11skuNPCkgJT2/N
G6XPUSALR+Dnyl+API1U6YhE2JA51wNo4uGDESFGBYOn6XGoV/OJ20i0x1iT7E/F
520ZfenwIjR33Rtq5jl+7Uop4z87qgTiDggaFOwJ40cNoEuUEBAZvB2mjPAcAmHz
sbD/fb+bNNKhBLxwgABwhZ05lnB+qaZHp8dyfQlWX5w1PdOQZlVLKPBE6J8q7Klp
zrCsFqMvuJ7HPdBG3J+8SZruwlsTxNwGH3DPPnawYaPGFAWlxYIIHrN3AMWT/dr7
Zlda4FpxkiRl9oZ3filBHDG7d3Ppvm5Un7uPgd5WcmolEVVxoviw0XM202tFXHl6
xzknz/mHjd3DIffN6tGTwECk2NGMtqrYrk80VmtNceIdj76c9ODMjIMAGR5romkt
OMeMKehQiDWYmOWHt4kROg44Tm4CYcUeNLDf4LZvSficvfAB8J+go5KIKlJkkW8q
kgXcHP8nPwLOIfw7hN5YNu6Z9YLZvaRJCJQJ7XK63ZKj2+kcJgZcIJZ+yp9NMxrN
BngHLPcHmlMpw9c4jRDKmNeyAdJxqfSNqqqTj3nBSEQXn/4+UupMbe/GBRs2GQzx
nWneBjI7LGIZRNRsZLsHZ4OV+0sDIj/vWsHYfIzFMUpZUfzFzz4oRt5IAeBtpIb/
DVIzsrQRtjLarX761Tb90ArsyfJnKQU4YWseNnOY9r+zaUlGeOWbYkUKXNhDlHOm
moDlyWC3x52C7FIN5EJ2LbCwXOSc0653mGTRR0cQ8F45a02tW+3TPOchJW8shQfb
M7qTl+vyvQjeuAyN6QQBT/QAobV/3Lyy23IjlJmN+g9CDL5sdgtkhw5BHuXelUM0
lq6K+bATdmUODKj9ajNk6xXHs1I/kvH8eME7T442lt/XdQxGI4Opte8kYzOMfQib
EDpQx7YFKx04+Sjehoj4DAJZKu79pQx+cJ7xhSjb1Vtew8dd8Q1DzShyBDkPo93+
44pQnkFi3FElbj8APEXuNd6yM5uQeuLqPjD37wjagMSA1597cHQ625k5ZdkWTDyF
hHRHOiQeGCVBI4L0i2AWtIf/saO3CQGh9rsnIfeQ5IfsXYmURAssN1ZrmwD8TtTv
gXNytQQHcHnHSvQBAbylrVVkmbIw1J0T4usVl9qUzbtvTyTlQrptuWhYaWj7K8k/
zisTe4Lu4qLfBm/NjYiw71O+7Vw+vbpcMH94xS/XFINKhhFN8xrKmUVaJRY1T0zx
PagAMlUZV9aHLASIGy5dN6gAygJrYXij9/WGZaZZJntCT0h4IHxs1Mpj2OzPXeAg
xP0uSmtRCJYtOuNcLoRizoEq4gUGICGZtuq7jpbddXpJGD2ASYeT0cmW+A34/VFe
Od8YuFsxei5D0WEgi5BpEpYmsCZxnsM8/AudjRMN+GHrsksmcRziok/A2t7z8UTw
DJQBv0tTaFdWxriHlcmyB0Bz/ekpM91jjiew7VyoYw18C5WdE9CR1SrkznX3Co9N
BP1z/9xUnvmSXIuIegCDty/i90bzAWbb/OBZu/o+dwc/pNSuCHzo/gaun6HnIbN9
l4YTQbRuaRDos/NHffDjkM8VHYHz6RZLmRqO3FuLCoziuCwYqrwp+nr8Zm5+KyXn
ccUfLcr2gWsaRLy2158UMtK41t/XrQ4UmFiGvahT/0O/vnEhbCI/7zCFiNT9pGPZ
SWpl34XSZKNsm2oSmqPZX5P09p1LBdE6QTeAgeuvHUzQK7bSWl3/Q4VFGVJ/5X7o
LKbe7P9uQCiBWR6Ole8v03PWCeUWUELpxpAH/P5sb/tKvMxLKWz0UosiRaa68Y1o
FdCGMIs0YF10mjPiWWXX4Mwa1yrYmFv3RPYg1u8KIpVb0kISJ60qmYUPBE3VY+zm
zEwMNzGsNWEDAlN1sbhC20Po6+NE/XjakHq44PYXWJOFq+d3KPZ4amh8HTFSvDUR
GjgNSx9AKu3vYuuqyEkizroJ7U6PNt1BX2iiNs5iC5y2ddzNltngXipgoaEmdBuk
s5tk921dAW2iTqfl1BxRegGcUFqiCFhlDiLAhmty49YdbKEQanch/mIJpgmnfqad
cYA2ZbKnBJkyGAD+qGk5nWKd65gb7tVeN6NSnWQ1eBgj+gULoeeg1JKyjTnc5cM3
NLTpK+nX6hIqt5LOQPN9gLS+IOXOw9w61Jg3dIuEMdT5Ja5B/4tsYyaagAxQsJln
1RQNUOcQtJXLsgkLROqNjk2ge8S1R/aEVOvT+7lWwMw7wuUKsTvJHOsl+EwqFhNC
BTNqekoGt0gNOoxwPy/UnhNF1PrLU0F/ysBd2yWi4eMNqYZ1ZgZhPMJiqZS9LImt
8h50C9fYH7Y+8ZyhTr89nHnoB/0Oc66iXP+MCbi/2YmglUEgMezIoCOFcfpzW7gN
Q0ec2NWUdNUdHVKPyFd6tBXymNSC5FZMdCr795HOGqG0Ei5pfFt5rhcrhEj2AHEM
5gof0poxfr1KOJ5W4LXtiUtr1WdjlbhoLd5jnYL5GctvrHGYLtsoWvqqetX7kq2T
TpikG/HxE/ICvSq1ZHfnmc5AY2IRkBiU/+ToW6fNvP4F33mLclBlsOCTPln81Mnf
QCVB5bTWAb41F7NqKhZ5x9jZN4C4q+csstbGcxewRZ1If9psfnPn30LK42tvV00R
0ggL+cKO73hxsyIpS4uxAPQ5Y+5Ti8MEL8sM49PLkEf40+MJTLaghhwqEMDks3gq
Mpbe4dP6Ubb5EoBKwJoM5qC4jKpEWCuGMrkA/Ihs8sLg+6sp9LzX2pL9LW9Nw5kz
Dt9P0TlNfjPSrhEuzR//AaG0fvYdAZucP+fQ57n14cQ2YrmR7aOJd4w/ET2TXF4/
`pragma protect end_protected
