// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:35:06 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pfYHNZpGTEfU1Sw25r/mTlRx6JR1nHwuyVyuSqhzWBRmTTTpTVOYz3qQMbMf54eg
/Kbv1eYut4+ZTinhqrcssOuEYsjWp+v5KxCiBO9LzY1Ue5y2u6GbD4GrM/fjJtYl
p8FUolUkQr0X9ZZqzPsuOtX/aZY0ulUYv8deWIODP8c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 34720)
g6uqdiA3eD3Bl/omnIqiy6N5k5JdYWa2Mkd6+Fvh/cI99Daxp32IDW/Hb6xnq94F
PKMWZPlTlLHiwLIlZgyan3uy5tzPrrml32MY/+3WLzeGkt0KXL16ZkXvAIODcAgN
8K1lgzGYpb5/vyKcP0cA+WVFIGX4c7KrcOImArV7okcs9mAgIitA10VWZ9mrgbyG
v3xZsxWIPNSB68AtGfFYyHeCpH3vJk7HJdaJziU14U+05QM6HGAhW7w9UGGwNXgA
jYCHjjNce7rEHFkdXrPFDf2WBhCtS8h5IeYeyeewvLW/gX+GtmAnBlk/jH/88hK9
aZM34F+UC3eJfBssKRUOQusc6ecA3I0/QreFAv9bUxQHfGC0ZutdrTuVwSuGmeD9
bxyrQ19KUFuEoac1IubWs1/hrXgAStT5VIMHsJHByYhM38++canHj/+jtfw516E4
l1D8LvEf3f7Gt3J8XW+RV97hfSFvqq0VxB5TeaioeRvvkTh6kg5TLYBmw9WDsntx
fMbw01wTDvEtBL7ZOe1iqwedjnYvJo4XhgnG3q1leaXd8bbADHpJG+adzJDz/LEE
8JkO0ADSy9HQXogT1xNLuxCC3El/ScTMT57JGIZIrizCLJE+RZ6tJatKfzVexWXp
oNay+gdD7WCSrhHkB2vCvhitHUwg8cWMLmVqB1Oogk305CyvhkGqTln2rdfO5xlt
IYkn839yHxSyn6BkR6wuA6Diw7XdiHV1YHa2dNwEKQuH7KyAMd6lqBXeRKYjl9hu
h9+kQdxoVNfULIqATV/ui5D9eFwFzh8nbP7sNHILCpX3eA0B2gle/z7mOFCvRiGM
HdOuli+IXPGx75zXkCXbASLMBHP/mRgo2cmoY3qcrPJADSESDyhlIx5JXZO6ntNL
ORjLN6x0mPq7/OmIdNQ2BfFi1aBss/9sqzVX5Lem+SEN+/C+0WWtxI7d+HQg7bkU
gkNTraMniRSob9TvBVknwCjqowlwDj3UIDzsqi/kplFswft20fkmLbhZh/1nobqH
WiXe0V7NsKHy2/VOtbgmYDYN5MPCyhTVLnZR1eUMkosJUACGH6xS6PjAbH8vdNMV
e5u2wlLqAnJ8KrdE+BllagQ/qOwovf7y0zLg76VT715nQ6TFXfD/8MEIX8AGR/u4
Gydoh5tKDKU80eMyclPLd6WOnm/31a7uYp3Y3InBNgrfhdqaiuBifLMVDGGstiQD
mQbKu01N3QfpNl4U0J8GV2FGOcr2XQKlprKh6XX3tJtjYXXp8b/+QdfZHtFMMl05
JBdLQ0ezzKRtkVI1C56HrDy8ejwNPHTThKq3WkonrSFO+yM5xXQfXxCD6p0Msflg
sKy233bTi6XIbzABXpgVszyeked0gZWUV8BU7kezQdfwwDMe1FR76h1t9B3hqSDH
ELw/E1xO6ocOtkJut0YW2PFV3cpAeVOCrMRAdd40AE3KLLDeuDGB1prraC6AQ1Rx
vwBQaC96yWAmuyQ4APmQ/B5+RKxJ7TBbdBDSSLQ8XLlUDK8rPZ8F6pWuFoQBGmO0
8OuF5ZVMzOV6dY/4tLLBMgLjjYmo7XJL0GG4B9lBge3rbs1PeSXcdbT2urE5vuXL
8ntXpQ5IoE1yCiZh9hRA/vooVfNyBAuBspvXWx0NvaoyBrr/caN1d6hBgCTKZfbI
NJ/Gmo18Hfk78w/2ZFLrYwupHMyducQeOM//FHNrc+dw1WmsBqTIHjFXbgLPPOCO
TCfQ9uHUYoLh6HV2PH5VFsMQ93WYpla65+Ca+4GImHoceQPqgDdF011TPxrZ1xOw
kFrhR7j7YwMB/SgYHgiri6BK6ewovFRHWAqps9nlwLWHyd+jcb0mB075aeciaaIE
UasXF8MmpwV6IDul8ycaVb1pizOZG0NEmh7A0hQUyo0Gu6iP1lg3IhzpRE1Jjkfp
BVqX3iLQjRSnYgkQhW0bbg4k5BOzQXibD4jAvx66/4d51KYaAcV7t0wBMrE7H2Xu
D/fyspPZxgvNQAaXa/7RikgF8ALmO45mmH0Yo7sdOKGuH7974+zI1d/QhFuupjHV
+B4lyukRR1YwHokp92oLtaSDQuF3nZQ0ZNK9xaNI4e2vaKi+Q4dZVxIvYWFdtK7K
48m0q1qP8YA+sEBQf/fxGy6XNhtqAnE4Q5uHbDCTNE6mxMDe2q+OhJfVUW78iwLs
/gvaxkHJwFAf8rQqtamjJSx6KHYa2I6P+ofnTi3CNKiRDWXfE13eJWaQ1HSRG4BJ
OOZGw1+bLTIm8g6n8o7xWX4Kgtb0WoxNXZ2Xon4URByW7yPvUEB/MbYo9kQgKOkO
M4YRS7efkF9kbV6d1faDPC1z4H12ZkerHB4O5riPKfFlVQn52xTWNcdTXhoa79t+
lWlLpgyGSrn+DW8sL3rqDMOULIZMf4S1nhAT5bqznJd6Uo9T6TJ1SJzwYPKLxy98
eXN7VrKv0pnR55RfLGRJBpTffgGZHofC+E8vG4pbN704QRU2HjeoY3JewPB5xb5S
upK6vUOL7I1J/BzbXCtjpP42EBwpIOqqWZIGRiPwhW5I7Y4oHvlEplw55CBuPlUX
916HwjEg11jBrO8VTJFPi1R6NcRkBqMvMQUXWQ98W9BFM+K/PwK9OeE0TGN0tUWP
Mr6lumOPouUborKrLL0R+YAN1YPLjqHaqi/k6ZsY2Yceazn2ntQi08DdMYd0mGmI
RgGA8n+LmTyWv6HgSKnwPxjOVL2LmcZa7peQFe7iTirOMD2RHGbzUSiszZtFhjRV
CHNwcMmsWkxLnp6IbKe+Vp16AJxyy/4MwVUX7Je549TkqUpcanEOhPoKWn5+rBjn
wurM1OwSPNsb3qBS+yYSInl+9G9ozfQ2fKkLnI5d2j3zPoGtATDg7Y2ajdRqvZQ8
rCgqTr+SNQbk2skr27CHxYIGNyIydDlscugfFX0mE/YKiNLMa+tbpvW1xEqicpxg
lVVFxHvahHqeR+yRZ2g+Y2mlOlqVJsjZ4zhf5N+jZ5IUctW7JCKEMXdCq3LTplU2
Fgc6s2H+5Js7zb/zYV7GLtjXKFFczdaQqNj119p5lH2JizR3iHwGF4m4KUUTu2Oa
q7yXQDoTwdTNrIjgf3otl3cJPuaC6kkwJSGejWVO5rVsZG4gCsl0kvjkisU1BFw3
iknJFmjcBsd2D5+yor3t43n9IE7MD2ED/2ot6u4fA9O3KEvOBzMpOQ5gmxEtUXJa
Y45AvoSHDdyRTTGqYqeflnJsoIe7Ul5T9Q1Mx2nd/2WXYUybkdBY8FMJGRGGjH8w
mAux1cyMtg0Nz8Jy5b28/RId0/cdjRByH7mKJJv8lf7gplBAckDH7qgPatoPqLta
rVkXjNzu6h1bYme1Dh8X81GWDwyQrHXvMoNJ6nL7A+/6RafVt1OVWMhxm61qMfGx
MetU0xW7RrQWgQ4ZYLauxgUNtF4dJpFLFleCIqDAjxgP/OqE+aVX16u1tZtaRxqe
OYRz2caKKc4TlpGDiL51/MVp3dxg6YdMml76aA0R9zIluaPftVmhEavSUFWxGumm
kxIyt/VwG6AzYOcXsKiTF5Aw7LFyJx03rf1gZO8LvBNe/O51EZPCFh+6hY0/nkrI
MtMuA7t6kLRZVLo8F5uGV3Adc/oP+f6o02MpCr9FqngX9LXBOaQFI0ftdAmk322A
CFSZXwGhVPVLvWr+7LPAEccT+DBdo2Oiym+CQCet9Qn25DSHnTLmdZD8IcY5c8/z
eARQTbDogt4jOKYtjEl9ck1fJNtWZzUoAXudTFNrwGS5TYmWr4du1sCcEHfYjmqZ
MhYoI7IqlGZoY9vIJ8kVqZUFDY5GkJLkLE6cfImiGY2Me1565EX/JrhKaP5iPqAx
3yB/ASF3fsHCpMiYm9zPBi49+DdAGvdVBNiUMKutlQnzuxjAjsKWKM19QPQGQi6b
1LsANaQUmlltT4LKDOgxF3CnrdioeFwfRl+8HOMRdKUuPVnVvTgMPRuoF6u6U7cC
cPioWMzwSKJMnzMMcLLGZ9Dup84uxaf4AblSl7N0GX3eViwddf2bw/qQtU87h8Sy
phYSzH/2D2oy06z5hVpoLH41szgCeEK6yH5T5oDv5f77ElO7K4FDL0mL6PJ9Z22q
iYs3uDx8An7GXfZNMUQGZsEQb8aI8oKz/UN8cuEFH6TNzWvBgsr5WDg5kJ6eifIh
CkBY/kK/yIJs1UOHKbCk4ClrtDl7v6uM6hpDz/u+p9dkhZsJPtFUmCT/MgTmconu
1TKy3FQ+prhFahtJgcngKODkFErHPuer8EDJwPk0L4Fuv+cRo4bLrgseCnq33pf9
lQq9wXxtHpS+DiFnwNv7u19Wt2YjA/roQcsq7sv2SIHlygZJYMdbWp057WnMAR3t
c5qrpK3nhzv4OdWzoDKkWOuTqjdlzpmMt72jVWJVjuIkeoBIHr94QCnYHkgS6Nbf
v66rCeXa+/wHXmQ87+tfZnSgjZ0v+J4tBUab1tcGXTrZtUnmoAb/MKruWRxfoMPW
6O65jdacLYIW+bgWUwy+zA22plvVrig+4PhiymS8zS6jzMcgY1XbeVHBkyS10VrM
QjBWDDPhtrCUD6O8G63njeuGSmVCL4vj06u4R2zQc9OT0ilb2v2c5j+hahFp0axH
nvqS4Qml8xKhbxUGC58XV/hfjDJMDToIsv03cXZ6bpaS0pIuuI6Q4GgUPwevVFuo
rPR2nV5tJ6f1t59YOriIeAB2hy7fpr3T5MJm44Yf7oWSupC0loji4GTbi4XC1/4X
o/UBYxAurQNIKLj55QmTdnPWKpQyXxE2km897l4WX0UgvIUVuy07jR3BDOFiY95w
W1Z/gx2i0C18gZCSJCnRSlVRxb/taWktFcGVGWVJ4nLA0BCRvOtO+u2BOQLQUFlw
anM/yNt7fR47p0aTA+8iQ7wsakaPOY41dAblqA102sx9TZ92Fj2E2zmUdqNMaqoV
MK96SxYNWkwM7t41UNyKrziA+ZaHxRgbWV2cqpSdytnqvqatVwSOCPBFKkIls1Lm
BJRT6j409tHogMSbe2oLyeTho3tKqrFIHvJaNBLt969jS/JZLPS2am6D3fZ1m1LA
IpzhJgokCy35LGMPc+zxDy3ckQwuKQdnSA2uMW5UUskUvPq6q3j4/nYwowz2XLIT
bi8PZ10dFHqEsvYge2TQqz3VKi7BAt8k70tIMVUOSJ2xP7dQy3KsssPY4kcFgD6C
9e5q7aP+c7szLuoCWO+MBgqlgM5J+lRM8JH1Lse/QLku2PWn0IJ2bMNOASqNwhe3
sU4ZE5BOKRdz/IdvgpPzkyQ4gtZvh+3eyT+1DZQAlPaB/zMfkCGmaMNjeN79/1n/
/GfSfy3QpOu5ALUmdWjUQJwDS0YF7CloEphLNqNt59IBnl3GEHMHe0vYpjpihGDx
IF/PCDjzn1OBOznIFdO+RLVH7EHs/Se/C8E8EAI5d3uKnbgaWiyz0KQzAcV/LQqU
ZMVjx9JtfzxsPupvb45Uv4FL/5GyRcRwCmVeOYlxydj0B0LF5goyQmYmjxdVw8Tc
Xvlclhg6e0rhV2LnFWAhn4nQ8UGmtRDynL2iWvVeuPALOzC3fcKpcNm7eZCnhdw4
4SxrdXKbQ7NC58JyzU4BC99ajXFUnSBooxqFaTM4cDlHX6Kj/5T0OggqcaQynn4C
H+CmlFDJgwelVrOGb3sYKpldsXNlJ27YCPfYVHsnRcuWWpJnH2bcJTeeuQ4hCmJG
B3YmB+O36ZRIxz+IFCFNCyrJf6iYBIfLvohNQJdR166NBVZLDVC8GBVM7sA/+9Z9
oyENopUQWKKVvqnHU2gdF4eJX0mylmVwqzaHGdYzEH7ZAkqaTkha3vVZu4IHR0vh
5jeXNQF++HRx80wGQC1vN/1k/yB4MVDajyYjNtQWQb4HrhSNg9fmsN/aqHf57kNZ
z8eYp2V14mQFbmN/SIPPPrZjuHpm3N8XGaQ1eJyZq+E4drp5X4mlopSJdTiJ5dBH
4RiWBrZmCyYzv3DRBLR8e3YSWETurmm6zEqcQNms/k7cvK8S5RL8b21PbQnjRPIs
PVi3X6574fE1wuFQkoQZR7D+oUD503Svvb6rXJRLrhM/ijqgFrLHMF4UzVIUdIVZ
tCbXsXrKNjvEKmL6VwgrMRWbyiZJl4DMpIwP+KBGut42wc10kr7A54Nd4WzlvjcJ
0ak8wmvirmReo0hjjsPfSZXRJb/CRz47wgGXboqoC62YCmhfFedEbRER6HIDP8G8
8Y8vmrMo4cqi1TrQKY5kgtymZ9rnXZW37yjGxG/EtBSPMkxCelYdy6YLDAF6PZxz
dXd7n5K8pQ0tzUx4Cq9oZCUbcyVW+jwpeLgw01Svy8MynkMqGm5wmoYLgwnbbCEw
tDbx9Fp+hgeSmxhvHSWLxnuo1p5G0mVAjZZhTlP+gMbjV/Z27iK/UWRIOzV9ddHx
HMVl6wVDTIgZ858//bKZRn+zxauPqUsbzK57wxo+zBpo3bAM7SMChituKyM65ydy
tWYLDFDipY+WF+bGjjIx+QN8cblWdkFpEjX/e9DX1ocE5siaU7ijpjs8oQ/JHA2f
Ax7kL7h+7Ern+B4AGQjwonSQVDIj0zPjcEABBabmjFfmbd1VY+bWG36Xt3YSNhQp
CSplJBFIOG2DtTXeshiafGtJtq9xlqRaom2TKWpZIxt4iCmMknWMmye8xEFaLpGH
0tFG3mexCkWUcAV20rlIn/BVhPCCXeQLM25YJrocyA/DQLGSWZu8fhiiP1d+kFSp
XMTnzxTyZFEPOm3lMijztlMy1cLOynuK9Cos94MUhvgP4gyFExBELVGBXp9TqI/1
cVTgNV8Eyd0FhGzsEZvKlMspzIxY2yk/7ZljpxM986n0p7x64+W3GeyvaCOf2dOD
36YBaXdVER6+hW1hsUxFIobbYthnXstLr0/2cc5+PPoGZA0LyQJH6vqNY7zwm6uH
+6SyUi2KsdwWuIU9vHdx+mlDTsT7EP3nspVm9xw3/2OP1AATGFEPOkzSd8oAQR8S
7jS5dOQsokhxuksK2oDYaSYbXef095+edMQfhK15c4ppvdRiwYvq9dsMohT4oT8k
RwkSZBzEnBvWdo7+X/uOZkRXBxtwhEKXAaGFOEg+J3VGcN9xwnTv71ULjLOdTyrT
nJBp0aySG3FfVixmIVWglDkB+yWxGtZEAue2w+jDzJa7qySa3wzUcK0rZxlzWwWf
/NuxTZvX7Ejd0Bp8p+5lx8c56IrxtcwWejP88scYm4ivdNaJ1gOSUmntmjh6/JQO
H3dd0Vuvv2oFzQeVal1mMzZ3Xi6zd5uLqPOm1b71GV/iC6CYTDPcRgcMsZBYnnGG
88xFQ2PdlhZh3/3MIL2hG7yrRTffVNG/T78VjNv2I67pwbgT3G45oWFQ8Gggm8N4
Yrp0BeAd8fPB3HUxqhpfu+Jww9w4/WPyZOJWDdigMAZUugnk6a0ahHNT6bb6G4Q9
T6dl1k85BjbvTvuXAa7jkMyS4OCb1MQbgRrzj3KGg5zlsBDEqZLZwBFengQdndIX
XBwkYStmleHp6JA0oR6OoG/caDW2XmI1k7OJGWmA/6TjD+WR5zHcNFjO/jIdvF8Y
q0bgC68AhhmoEHVV6JkCC4z44Ik+tt0FmHhUYR55bwSOOxcifLBX5Db1kPYmG8Ja
swgW5+qhoRSqGRDsF7btrU2ElSrxM5FFDm9BKzlJFXBQyuh+7iiGDCLEWlNXU9Xx
58zJCePfhH3MSj2E60YVEJJCxfd75zMUx/A+bMIRFnfbOI27x8B9KE9A34+tGnl5
7R5wtPHih5EiR8Nmj+51WWqWJ4OW6819w4TeR33NyLoDsLof3/AXQtRf9Jgo021k
0dEmu2YYj1k+4zHqnS+dWqYVk7LWJBC9c2psejlVrkJFmaMD0Vxob340SItRIv/p
KVbbAB9DIEYlddJLenYYx7EKzdxFEBtEdINyIJkcf2uRH+W+KCy8+ku7JeRhBYfU
6s8+w7Tfy+fOzri+Tza1xCI2WVT/4/xhb0phfqznlW8qgCC3+cEBV2TrtcHXPgix
qU9BlZjKQcXZzQh8nyxcHo8dojwxSv161KYJ19wKmnazyb3x4kRs5Ll3919bl2cv
zwDK31uItCzZY0r5SokH+5juGQp8m922nIsMskQehgfv6nw9GettRj6burLFoJrE
pB1xuQCCOiqmUFXemiiZmO/WOp4fw5jgEb9hYCE0v49kl4WKNPWYqHy3eUGMwd2g
uYFJhOGXrgsowas5ofptemed58DQxr7Um1DKN0nllY4wZBQfn9xGc3+l6u4JO9YW
U3E4RR+Han0JBNZBGPkAGpKTkVJw9M/faA0NfDsPzB3/y1nB6X/gRdnCgLGsuUGT
f32MUGZZkPyStS0vRqR466pulFVeqyMdKiP0n+riub9kEBfGA0ZnpBzAJGwLNz9j
oZMjzGJhseU1XtBqWgwtlSMkyPPOiuLRF7gCQX0KucA82Ign8EXYpyhK5pv9Il1f
i7XdfnSG1a4H6uP6QrHbqW4ehloBcGJ79Pug/cOLJI+HizhhdFkfLcEiVLDY9qqk
KmPSx0HlH5/61FA9BwKYkfHZ94swh6ogC3j5wMzyJrfMA1k16j3ghPOFQe1XH0jl
iPfeeZIWtA6Ex78SX8HtrLbJHK6J21euswh6aXNlZl+lQpEt8MgsLFsMmW/abWtu
3g8QiXL412Gra6RSnJSc3kQmi/PutimACsan+fgVoG3LYvssX8xwxocNBH2vI6gv
Okq8UgOxAYJteunnVOE6Xzv4wZUYrFVUQJa4DTjn0rv3EiCjZMIidDc2uj2NSkvr
YXib+jQHmLigI0cxcXU0Izl6OXjY3w8/KB0S4nzs1A9h71YJgcZO4ve6b+muQsfV
6/lVBiVpXuDZ+74nV1hA2j1ob26LsAesFtQ+3aLqKdsccR8fnEPRDPNejASejPaE
oz2RJun9cY73cSoLKTD7p607azylcC8T0txnNrcAmk9/BgXEKANzCC2/k6e/D7NQ
eiMeHP7pP7lOA1z4MB81Oz9eCFsJzoqTAuUS1JYtVlGpkH4Pvt1oLhkNBoXw10cC
AosMaCrnfpsF9LrBxK2aDvIkFht1RBNG/L+LrV3vM+tyhy4EtmXgoAVUdt6bfGmE
QLkeJ8ZxRff2sXv/hZyK2cFkNZb0dLKVDVjgyuDDWUmVSO0zdtUklEzruZQpnAb+
5T0VCovYj8h20eDl4a/E4wq/qlTxLVOEaykSEr0NE+44RvoeOVihHMRLwwLFB2kX
T2mMmSD2dU7FA376N+Y16qbZpISZMmzlmoOJFM1xPzKwOlGIYutaipetya3Gl2hd
nQIr1+h81uNf6b8n7hSkouvXE6gQheQOmOxdHeHjUc6DDg0KYGCIiqn9xLl9nvaB
19Qmtc9Hbe6R26t1kUEeuVyETahEI/5xVoVo2QNE3M/drgEmzggVz168CNJX+8re
mnYaMUJ8/Zv4l2wesoT7DTKL8ajDg+dAzhP7f4mBDuAs9PwMrKi2n2Vxxu3WsyXO
KtZyhdaQ1ZRujk0YCUX/lqDhDrhKYJR3B6rmTSSMWuo67m7FUCGlU1Aa5pVpDCak
ihPYcJHTdqunvlao/QIBI+xqdneVJbb+bb0GE9RNN6boyjrY25qZWlOeJPrybXso
rTvUCK7cdhKltT/txQEWO3+VD6KlqrdhBSVR4hvOZZhg5aQohnCC5BcwDuyFZNhQ
zE1JT7TtqufKU6VmQZxqFNTUmyAMjfMC9CJTO5IPR2T25JE4ay4oTMn688O0IdaE
AFqh62O47SMWLVLe+dUittJVh2rE11JVuwTX/p4fpXPMA3w4owpgDw/eUR2bkk0i
lJlAgvv62qgMJoDJthAmy94d9kEaz7oeYNXVburo35PIXnjtg2TSwYiux8lYw8A+
3Vy/E4ruBfjohZRWFBNu4rDzqbD+gU+G6de1nI3Kc7f1n11/OmlLrdBP6oUSQWNz
/0O36/l0TVjKAZKdAfd3SMsZwfsKCZGEF6+m6HNVpOEgAY7995mouUTqQ6Jo2P6b
dK833iCzhZRuBOJwYvUa4jh+ZODrdAqqiER9S4oeoZmpANsxXpPk+SASEz3a2EY+
9P/geSOOlQlXqV5H+uKu1MA5uMgQejaWQk9e4hHmlx/naw8mu8msgqMYo3SnrLl9
Zj90COois3QYoyPKM5H7N0sly6CufELlyMmk+qRsCdh35dxYuBjp5Hg6RyS1HoWW
Kh5vhrO1t/PkMB7gkWsmO2kXfurzHQYzF49BolS387rdY5piyKiFlgSrEF7IcSad
FkqUvpD8dJcN3WcJFOt2WiOAmsuj1yWJqde5zocpl429yQyG9Rv+rjOEFjGXL0nt
r+ChBebiUJePg/3xepFYYb4GcdIbrdSfZhZM7PuR4Deu+asYF8XfATtidEvHrZls
OvBeqW7kBabHk18maSY/ryAOzyis/S9emwYkiteMyHfcTUkCsUNKXiFKuSVpr55Y
tpffp7Eiu0CoOqYkZAEWyRmeOhnrQCPuTkVF+8rKlA3XuXRXxKIPvrNYQiYyyW5O
JtrkVJQjXsDfq3VFA1esqB9WWTNVTED83zrE1ZOz4MxSBCjMD0zhpIvEbMFNq/a5
yQ9tClcBmm5cX6bqfPcRnhxH0swzy0WfifLI+8vGiTFUso8ZxxTlaIiznpmmo+z4
Shvmp4oinyjXdTOsmFrdWeL7zk9wVpWKAUrVLzgr0I+r9ugKnRCbHXOfEacmh2lb
8WmAgLQYeYmOUdD/odouMC/12IvvwsNscjyGa7yeGQBxeeTXJH4Er421jF1gz8Ky
E2N5lD9Te9bl4XYyoYllvkuPme/5aCMvC3AaGg6+2lBsGoiA8tLdTaD/G/2FczFC
oShM4OY7lo8eKWN/AeTjyJ6oIYHUY5FMv1eVTW3FHhfwxwe7oC8csnjMQDddHR7L
GQcyrIhfZptZzd02GpV3AwnfXkvYlrPQgkauWtpYRynE73TrzKu+PkpeypO+3J0M
29tAbOyy/V9EhOw9JCPa2AXzqvPkldlMdTE/EGWRHskdlieu1fQTSp9JNaFituvc
ONz8Yb4KLfDMmmGNW7clvwwRsPLuf+4R90M9wTygpZ8f1gHwb3tpdyhW09jCcePi
Jy2UkQJAX4+DCDGAmSBMzWP0ijsLb+MJTU7VVUfGUzYLRhJ1mrP4iT/ulh+YmbjN
0g7PqN9/fm3Zy0BpGR43vdUS4jboWLBqDniHkARQQtsmmxNKJCNcnfKn4XzO/Z39
IVasHojGkLJ5tqGesNDOXOCqRZOqGbzcqlMTg3ghAXYlZYE6z68T2vjwwdDLW87Y
FZ4J811HPPH2kIyaJaPG/8d5rzI+0RemhaiA+zU7UZaOXJq8IJiufucOWBU8tQ4L
GcTDWpt4QiQnr+adRa7qeo6miB/BC9btSbtCiEkbYTLyOlAPFCSvQaYiqK0fyPLJ
UZ2kSOwdKNRVg1Z+S5o2aFnVsLOHPUi3s49jFZCgo1y+UB5UKE0a8WNeQlLRpqOm
MJ6vULnYypjlMFzQUTXWEbYirERDbIl3OkC4D8J7IfEMuWjd41VyivblCIRIHDTX
5nx5PfK5V34IYiuqmS2iuPEKWczUQiCq41/lGy8SqYB8JNH83ihGRt+qsBjMOLvS
C0Tgg5IlS8yUMPLIRLwjgyHreGba+GcYVHApeIBgvimbQ0utJwWlviOY6xO//eBS
JOEA5rmGIHRTDJX3Gmu5lnISFNo6nSx8PhD38gAKFRlvF8Mtfrw6Mf62SHJf3RR2
403pxOXXgekhMiAJenvcUc8S7xDcXi9TBOe0qCObbDLyYug0hJ7oxnzH4OKpVEe2
0PcPaGwgu7hRDxpzPEWG7XMNbNKKrf11LZBtYXACXqGtLgMIogXYMhSMZ/nTB1Z+
6/kyDQ1QJZY0qDvzPMVbWtYkde1wf9gssvn37KyozmJX/dLHAi+gcUpXzo2FyGJr
1thLZCmc8H6WuPwEKhb17JE+qinikvdIu8prlqmuD4uCKX6A7xblb7tHTiB8e0m8
0PcbqE0zftx5gIo28O5/olrpo/QOI+8XKOwnm9h35/S/fa6nAGu2UP3xkC0P8DtB
8Vgl1WuDs3azsv8sd0cjRerS2n2wJzUkRqb/WuW9Za+hTwr1zpBlh4pPPbehZrx6
SgrrXdkuuks9BJLtec5dGU4FoDsaymfPeu11j7W/t8fTN1k8pgRnHeCCC8K52FWg
w8jKuan31loxTzbKCKf8Q5T2X/UkKupIQ8eNPV1INCXxXUEJJMWIBfpm8CRA4yyv
GXtIB2TaLzKMz4GXgtz2XF4h72CTjs16AY0NgINGbuHi+JfwYOcEHPNZSD77Jguh
J0BnWi7K3LZwCv933MEO1HlpwzIyn2v0nxuJKeXQxzx2JOdm7EKcPxKO3Y88Kv7F
7OX6hDU4R5LZ40b9EwgQCSxo5vAgsk/7DhAc98SPUtIZrUUdmwa1WdNTOPGK0Yfz
RdiYhOt+prUXBrV5QBbnZe4nKyHbaZnLUID1PXfDxFrD3X1hW7KylsDadV9W2e5F
RTF6Q7IZMn4s29iolts0hwLZR9aqk1mDtU3ojgYFEOGaiSlon0qJsmFx4h4IH5QJ
zmJy8NJhc1aBUGoxJ9ehdxISadzTIumlKApgmCiJR7FzW6QDJW6Z/msGauTCE4QY
QTeN+/Dgk2p7Opfpoc0pJLea0N0TtaedgP6StD+CiM62/QRbiXVZuHwPaFlDAB1Q
/crBDja1B/uo944opcv/iwAZkFMcR+8Gq/QPvK750xXqB33aSYCiLmFuSpGZ4C+X
/K7TfqTcYjsHjlinlba/ldUZBX0Ky8vhn4pRa5CExNh6JFS8Ovy7IwVkvly5MOgH
qogP4HI39l5uLaDTh02EaD8kWhUAnevjUC8/eAWGOQg0kU3EIoH098YI4QUHJJQN
KuZJP2+m6EtrKGbpTdESZsz7Jn8r6mIWd6y4XY9N/bpzmDp074akrbft7y4JhMiv
5bzBnOI/PSL4ClpzmDG1bzE9j9wXjTYpjNS7S7t/fKiUprGrJ87epz7KovzM4QsF
YqTphrlud+LYFdlK2nYZdr7vMhy42vMK39QclCj0aqxPHyi2I8QyskPMpY/v31UE
3O7+X2zZQPGI5+22sLgEr0C86jy6cBwJVuN/sSQcCkTaB1/BOYVa/kor3IKGGREn
86Ow8oTQIjFgIBuI9kVjislJnEhhd9W9jb8uc+OB89U5oH2E56YjWAjgR199r0gb
plHbVeMkI2QUeFMHONIZZvVbrRtflgWNi9QZuv7PdHl4gFnJLuNAufe8pKOit/0q
/6j6S0xjgWOOoqMJcqgyn0R4LjURzBXnLrIpQTOqlnIMvXDASgdP69fLdxqaV1Og
IbNvmuI/UPMEX/sirfmEuIv2pUexUYC+DrpbWyDSiCD+OIU3DT2WttZY6FEkVB3E
xf9xwgrqAnchHwMoiJvMjXzcyoGz7HlekOrrjWznzBGx0aSGvpdFhzV/dK6rvtQE
C4loFJYDsOGssbr0OQx8TsyA3+ulj/lzFaZGU6mGHhHVJzMc/kIm3xQS37E0xQad
yss2wmYIas11Mu5qxnl/XZxjvIhY3p3D74XWbYEWcTX371U96kGHSWTZMDqe38wX
6h33KNRX6kYN9/DiuNqKexXmO129XIuzyABMj34AeY/brQP/ITaPCEymOyD25rkE
ix+9T6mZHktoA7D7BMYqydJB7JGUvhcOQIldFsG4cyHmZrZQ/mqZFWQmF/7TKd3B
zHJB+Yr0dGuVhD+PSMRnw6DVZogS9xBTJmblLILQdDIlCVBnHbmwuMrgGa05QuJ6
CPD72/CWcv1a0mEk9Fy0Ee9RchumfmknYMTdT1WPF7hvYnfD+KJKHQZzibK6uzEd
5fBuadkyln8impZ0JTlm5Coad3beHzreSQlRGxtxcn2vcfb67nxIGb3YZPu0Yt1I
9qwrZbc7X+tVkm84pcaOu7hSlYs8On352wt/ioKtslLD9p6V3O+An11Jo+ns0cfS
iqUZxUqxYDDUbqAvRiST9w2FIKNdXC1T6rdLqzRYe3yb03VUw1mqujPW51+hliNP
jUNyTRMHMI266C1YMAnI2ckD8xNWivlDwbEKPT7eurOCi7IiDWkpopJOtZneuZof
ZdYJO5bXhd/Zf3DlPJzI30ppIXHTRe33DYwm1zL9N7S3nI289CpIlq6PYfkWXyi9
KPfhn1RHervEzDKW3CcGqdo1aCEIIxWZATBimizobOSFa9RPu+lePNUYU3wM9Y7G
ClTNidCLbVoC1Rv/T7IEeg/03ruw9xfHhBwGujveO/OLWHvDRjL106uIzZ5ShH4I
TFH4OTYrjzmHuUuw0jqDvSpd2FD1jnLfP8XQ66tHx6ba+4yFn+2bAq6A2pq1tKqx
T1M5iSjfo0H3PxWZLqhZCQWuQOXSipqG3Dma9PUbZxZLTALFYVHAmb3KS1pbvj+6
0Ouu9Dgm/Pf8bEJtpZrlSChczpJTGW7BCTXYmwbQyNCl42GSlyqoOMZAwWMT8Ubx
1/w0E5nB1xXKGpNWkZicgoZHugX4bofBMm5msVsvxeA8ckxiteDzyDHu+Xq//T7o
DwDVoCjFJwAxvs4vYwnt1NpTV0H3cVn5YDy3EyeFShNqnmG9r7g9d8RKM60IZ1li
8vA481D2hEJ3ywYwzCwbXW+mIYNjhGqU9aBgJYYAqWjXjj9LQPZcOOvaZMb9iEUQ
wKTQ4Q9yb9Zpx/yA22Z1asRBq0wSNxudWiQG0id/mzXbheHBI5uE5xrh9y+1V61h
TtHNyIYauEQDAM9BY6lFEFRRWLfL9AXjkjSxQCC4FUD0L9dTYqZb7iNKD4uoWime
uvk4Xbh9sUIhFGeaGFTqoKHPBv9LIosS+1XUmjdiVNdCToKSn2EF+ky66rIIzDWe
Kwey8vg9A/AUEXhLNeTLHjEkPzk9ND/kZYwjYX1KcSVxfhQ8V8ynaj/YomZtyoHO
+gc/v+KRU4FjdFzNCqFpO2UCk9SlzFXs1gU1r884cKbCl3zLXRKwTWWbyKHSgPsj
/f7jA2Zn392YUIILrE7kI6ly7SmmzSUAHmrOsnMxrx0ESEdYoCKzSZ9E8IkTFnks
RPgWqqhPcTArLg5H57LQb/Zri6rgxjv3rV+b+Ukh4ehgtSVBzp6/eB/hq2Wpw1Nd
NH6/YYiqb0jTBKXqHLiNrcVsLszijzVpQqxlQV2OkaxC0zShkjsuAxnX5kU0KMOU
badN+Yyy8qxmy9L/BEK2ASd+MOGgdrv4KWXPT/L2fHrhh4DTQlTGkpohA60pXkjj
CYA4lcLXfLxZl9eDkJdyXjHZCkL8/5Khh3wcBlsYwyAS0PJrBpzQq6TBobel4c3k
QEHGo47QKSoYZzLd+oqRbGYeXuk/t38CtTcbT3ULVnK3ygGS/jzxp5bJ736wY/UA
fOaI9Df5B8o8NmuwILnKBUEqy1XW+Vs4zoRtciWemgADLPbyjNyR9kkR/D8ltHqj
6Z+6fo/OlOm/QT8H1VOcqmn+QmRp7h/klbbKf+wIqCd5AkjhJNiYG8haXqbzZHda
4Auh4Rd0p7NRhl5rFCUqtCeTtDxQrn9RtFq++3naGokuhXikT0ht7VQcgOquNT9t
jC0O9BeuUC4YSUtVHIJYOWf5alrfTiH9Os/xP58NO+yvGra4cy2KEuV8pDt2J0lM
v4Y9S147MHhpnZd3fpJ05v6pe7o9Z3Q5EgZ6HyyFhP6UnpkK/P52A3O+guZm+APW
UehGd0f/LKcjeTGLH2nF+Xg7YWogz37k3TCKhMTJ/ZNrXZCr2rvM3hLlv2zT6Bsv
gu/+CMYrcg7vIrMs1rAzQ/sko1L4kmnVnIA2oIr7ha6sCAd5TG/IQ7r1+yhXtEFG
zaszIqi2l6IkXoVw55+vRxBQTEcLvAHUW+lAjs6fawk5JDvqaUD+KeHyHc7SXloG
tSyiCK/SNLoBlLkZz3QT5kJ8tCgATXurdJuxgHj+mnbveWevIray6RGJ6VQBST9T
rouaqcjj2x2EdJHFGMHBHv5Q0d52VSWUf7YKLeBUiy4gY8cSnwwc5/J4XRUP8XB6
1XloqGIRuDM6UAMY6P5EcJBmCsMtOxEFobXYCvLKs43mZcVeWWVGlZ1efBIC4R9f
Rq9ngM6nfnEVVmUmnr+QZ/s5JCnTkplTRZw5uZyulnpj99q2VQArQt8ku14dqay6
4/9OOC0czhETSbFMfrABFmdHIh/fkpWc3hD3Bymkq03q/tjy+XGXCl9G6oOQXRib
8F4/24EHlzKpeQhx4gElAlluPd4CyDzTc+mYA4AzLbl8DogyuIRAhsYzIB2stjKE
wh7Fp2oEXGqjtxJXY7xdGZyvPbN2tjfrJehIqHbuGfdw91OxqNp0eJuGz6dfCH+G
xzFF0mj+P2j0xO8Ep4P1AK/81RXy4L/T6FhihoyyQAroweeKHFgS2iR17BtlZlko
fOVIyIXo1OfxkXdcjNFnzzVZBy1DuhfBue+GvQT8OVgTwcEggfxWW4Zr5YzSDwc/
7F/9Vsf2iTHzGeiOuXvsym3glZ2HDRA9wwzWzaIZL/4Pv+8u7Oj1s/ZyYgcMIMT+
r1+ADULlNmtF4YEw8rjBDn2oM+nK81RCUSeF+ltmErl6L6D6a8ZONI3lmOlWKQrN
DmB2s0foUxOJJc+da2VcEQ6/g/y2VCPS4iW8sS3Pjxr1HmL3mvmbtC1T1aoam3gM
0XCF8USp+MOSzO+sE5K4nJep2XsCh/cRQELT/gYQ6N1NL7ufbfkP9SRoKcn4l0c+
5ay+6iqy0yz126UhWpi+ID2v9kopX1dfo4oQ4TDReEZo6FD85CVjvXUaE70FCFTz
aMSSUIXhDKWjTwKrKXXJ8/zdVzpaRJJwHG/A8SEoYvwVCfUNYhJTe+PeE1gX2Xqg
BcCLDkGy/tGyg/9GBugM1HdSzGkBsLaBj1mBT/eLFkbON0Vvh8LVGcEVBHtxiPkI
zgEusN/wY5Ly0DULdDVVZJBuw/SIgy8CXrDW7pQ3+7Ac9FuERPwPe2Y4GbVvjDLY
oyDjGzEovUjKpf3zXtPRP+6nXqCuU6Q+4PgvV7Hd0WL3+GijhCGxZ4Ze09wEMkND
+3g+/U/lJJsZphVZKRPPgkk6qwAEe5xduf+Z0VuG55UHI4wwHuxd0zWEkmPaNbSm
EYV0ujx5no5Me+LA8nYp6p2F/q+u9pBJ1g7rg8mpNrhst3Au2WnJgjbGG53BAp/F
WorlnJQ+kdH/ingRM4GNrSnxQ+t2jrUeZksfqYGOVakCMEj2EJqHJ51MKAIDSkAk
7e9pI9i0YAxKnjp0JSFKOr6esb95WUKu43Utoq5UsTXRvqY/aHFfVlvcc+cNmxIu
HdXrdx7FrAFc0/IwrcHO3nY757HR0ZcPdPxI5FHQV6pW0hhAvEybl/E1mwUEB1kA
Ac4lxex4j8++smA9NkqaA3y5g0UgBcSQ5Fr6YUgqV79PyamgbssK47vrw7CZ99Cw
3xgyxXehAJp+aKJ9VPe0JGTxzF4WXNhPQQuj5pwV1/SLby2ObB6WKiK7sP1Xtrps
BjPohzoNWRppocq3ym4iTL3TLTB58l0nH6+F8DTLIhnnEvn6KA2zmhZ8Eqf7oCN2
bYiOTdDibHzbrQaMyhlAI/b8IVapKozf2wkGF+dHEB47JTlqjxqpfN5mHZNSr0At
Eh7jY+qxHSlMt6UM0TDfE15O0dLq7t8vAsrLpyX+lYPOkkG5czJPFu+tADVi32DB
PBm5L4sGJUDlhAvq2W5mx5bmq4od8GlARycliASnXJgQ6VmxudizsBHJNn6vbfWN
OAi2epIBr71nqgZM82U5j1iZ91z22sCahQxX11Xdzt04L1vSGf4itHgf74txZdxC
03gDNTaanDeoQXfTUoS3leMxuRCV/4ktRrjl2kRVbjxq2JSiOwWp9ElLL5Cl0ZY6
qX8PylNbK7HDUDx5qovpERM8NyhabKsrrIheM7QpF031FTpMdvc2MPZ6AFe66S7z
OrUjKIYc2mEIAqYDTDff1cw9nmTyMYK2BB7H6BxWhxn2p2WK4kvuXQKqEtiDxQJC
slqwTRI/ETdCtS9Oglxf4nf3X/ywWcU/M9IiRS8rfQaaEkwKQtSK96Qh25nJHCLz
sHnJ048PLcZ5xiEFlwYxCIAGD4ngLOx68MKgTfhmeoh/T+zw1syMo6BZdo6VH240
WlkRMRPVq681IwFkc4Hielv3Y49oqLVV9qjt5r6yVJrYFFPTNmyL/y0I1gTJRiEH
/FAeM5sK6oWkh+TkQeOvpZTOGjJc3Xr8XZbQdrNsqg9TDaxfLdd5/7eykBXE7eWG
ydIdp5ylHyYQQgMgmSzhuvzdmsTqrJ9ZBgknCiqa9/osKYLESSkx8eoDRSMLEuUG
Jz/57Q+7t+IF6D6I81EJsH0XV8CDjiLtRBKjhDjZZXuPYDe/NdF0WmbgkSeUXKGI
hyLrm0BsHXe8WnQeuLu4Qen2NzKKfA7ZZWJ9Xd3+K2GBLV3zpnyDDjPXAZk/Xe8i
H8UgQKHDcPnSCkOlPrX6ej+OwjLu2MAUE6FQLiR+wEogMvTlnxL7VmXLXQQQzbZ7
vBsszSDnjSoshT0NA2lcWfj/oWdDQ5Dw/5MQpzQAKfDXlXwPSm7RGBlOQ7M6Mrho
X98k3Rie8hmsMaWhaQfrGrR2rd7nIumbA2sYAoZfNsPoIBnKVEEvludD/pmAUJc0
3pwu/aiOozb8Pmc5o2/+dlhIfH2kOFkeiep4rD2bXZWebd6PtbIS3OwnX2+gPnXO
VK6OECVuxE7dTNwn9bhRdB5BGNSR2Ni3bUM7irG/gMCNcVkXvZ61zW5a/RxY3NG9
3ApAlSytazrQyIcGAkApGWO9kXyFzgQ/K+yBZRFyO+Q8Vyo6i5oL+Jo7r4kF0Fgk
AP1baxpAZzMm27G9v3dSf8osVro821bFXcN3gIsC6uWzavZlDdNoQ/aIPHSLr0CN
bWRWvG9jxrG6sXUmi/2uOW5R+Ho2Qa6qyuTH1xGi9CZT0inRG8TDDTsYWOUII+w9
kuUCOgQ/Sp+Dx6ai3v59FIhJx7zOJNUMVQ2rz6xKFY2YCoDgLD1p+4IXxMOPj2Pk
NsAwHuk9/F5SukYNFC/rZjuRm0oly6YveTLgmQrrNPB+KBvyz/n7Mcf8ixSU7Oqw
k4XDxyq1sEyBfU3RL4WXruCuxx2OaY0rZ0p5Q5nnkQS/O0Nh8b8UoG9L3LPd0SGi
QoNAoVmiOR+RneEbDBSdoIv8vFkIQEqg2AZf/GEXrJIiWkohSegFnw8rj1VRAUtw
z8DCtaNvcQab7cCmxRTnNNQnz2mfbI0UxYEI8OUNs+9uoFs8FnRmhkfG4gA9Ff22
fBoJfIKoKfVoQly4GyZEBtnrx2fwImHVLLRhzsWYamqGoZWo88rBscEFv7eDhueP
z+fJiNs6kWUsG+mDTa/+JoY++LUQ1erhnKNmks81Rxh/bNdMeO3hEPu4ODBAJba5
K624VNhzoobOOaso4aTuyAkWMpBUTD8Km2GAzkrH0yvl6NAb3xeIoNI8Ns0qrtad
4EC4s9SEov2hnMxWWsEIu5iql8N7vHvd0It4VGC3G6NX90Fwqc+QiVTKxB8dAXlv
88lzsmBY2Hl31pANIuTyRc2yCnfz3L0TYBt3i6Gz41irVTeArh3x1GnxyWASUnd/
4++5WOYAlMzDcAYv6mHwMh1vDU7uf6TsuHETGWeNv3PxWtWczskmRHAxqTSHa/yW
j9x//FtO0HC73pTfddmrn40OVEWuXOIEYmqFkQl27zDb3Fis7Uh+4su52XrFRIcH
Hw9uI2r49kU0w+AWp6s/CXw22kD5Whpy0tROeJajMfLUvjeueX6h2dsY2NHhe7YF
Bda07NKAZJo0O6Ix2GbO5Mr3obE5vlqlKH/2wSFGPI+Si0isEAxHQLE5CbDLAuyw
VrKSZM72XImpIQFm6ZQbQpY6Zgby2e/catmia75qHkeGO1fgeq9Wu1xDSNTzFYQB
FOXQ7Whagqb4siTJVMuChMq75puFBtnwml+WYseyytuo37gJc+R2XS+I1GqVeiC6
NrMTNo9WN5D7vK3LL8oBKhQr87c9wgYjIUatLULYOfnoj8ntuwDihAklgeN7RrER
u0Ax73gavfyz2FzjRgiTeARhig01zJEQJmRzl3zvyPq2ijNPtPYUNJZDJA6Nz3rk
EEt4epUV5gwoBCzR2DsEmHzWo9QnMwF2a1kI6Y3ZdkjaaDz2I0El4WDQ0aehvJhf
fNutsq8sGTRqadntTZqcyLlpWGbB1Cf8DPQoUjj3eupU9v3l2iVM3za2zStltAs0
sgkFPaiLb2oggyaNv4AIQUQjx2eKSD+DSVTaUopiSNvgfLA7zZSbnYbCNFD2hT4V
0nJs6PF8nSsgdJeGky7tlK3hQBMgNareqLnxPGtA9bU10QY92u5rd23FuskHO5Ec
LVzd/riBGwbMJS9dD/gbDdECsc3v50nb+FkrUQiDjoEumqhRKe7t2fUi9VgzjAki
/Cd8iG1/mn3vVMTUefA7N8swTH7mnNe3tp8UCSO4Yfg05iyC4kuyEJx6wRwECQ4l
xgG4Jt3JbEzbwstZchveaMbepV2rrUvyeGHCzRXUzSFn6FwJ+NvxIek8nFxJyxIG
e4atcVaV1pPThkN0Ujuj9ysX/MNFd1VVzURzMqQyOgco8ipCOguBreuVhRsc8/Lf
aox3lFvd8WjCxQD/9rr4ZidQM+0sBU0ijXT2O5TQbQAIlUPTlZPClPCxNsoalDfL
KkxRcvONiIJ2BIqehXpL7oxFZ9nfAhRrbflZUeX9u6UZDdPJJMxFrvZtf+w36/hz
L0/JcEHhUv3qx5t5TRinfxXQVzKW6+wHJkd+4QVLUylRicJfYqOgrgUz3xpHLqws
QIuDhtCJCZr9bV8RO1Gptm6E2lyjlmVW4E+zo8QtwGwrTmW0dkQUPO/mFhuB04i3
TiiIQG44zsu9oq4He0Xuq9gbVsJRD+Ly/yS5hEUWzV0hGY2F2wSFC2hcDsVYu1JB
6/qa9oezDcN1w6nu/RNYBhjJYw8zydniAfpddU+IHsKwjqfyPi6/o6X1UtpXK7SN
oq/CX+NkgbaLYfqYC0B/nLeyX930HcewKcwfsXzOk24YCbFadhRjnoA7tzLpTY7b
a24B9NCq12VQc3U7gzbiiX31qb73rK0YTdNNY7d8th/Bio1+mv9InuUgXKIPGqjz
bGq0RPENKlP87fSndmY4MrLvW2RDpKUgt3Ha/drTcByOwHNUT0A/S/a+OlnMM850
bIM/mMRZGkZoGuJ/S3ecTgMD+lbsaPoIaAfzKak6gdW2vuEz5QlWsmoqyU+Bo1yM
Mj00f7Pxxt7YYqpGAZ7HXBkJknrKJXnAXfMFwMQzqCMzPX+XbCLiwBxB6QfrAW8q
SqPDyxCCcARTFYtrz1ZxPOpp9Z8RP9kAKWicVDbfaM7EANMj8UxSPFjzmP4HvY8U
BuiVzA68uYCE6Rec9+EzmOCQfcXKMmIXFGZ9V69zVVM6cTXh4j1bh3V0hBROgn3d
A6jX7Wvk2YCNwK5EWsFIxzVPl/YGv1Pm6ewpc6gaFsRy8GpSvH5uIATqj0y5wpKo
gQgDi3EIGATgBY5F5CfS4ets096TrdmuQNiOvVQYG7RU4MuXJ57gCw1qL2a6mrfO
CnfxbCVv9oWhDpW3di56faaG1uieHVj7Na5DAJU2mSql1Q8VsypOVwRfNzs/z84k
TIWmQVQ3aUbXa6Q2bksodh1bFpT82RupPH5ylIUM5TwU7o6h+EdkTaDu7z+xeROP
F/kWikoo7lX9yC19Jr07MttDvW3Kbye5ziaoau32HWBXTW+NhknJ1Pm3saJ1ffVq
FsuszJ+5gDH3ni+yjsKzzqF0hS8pwivW8dsivXQ8V8I6K4YbxByEqfgJCiktvJSK
vpn8VFZxsypegBgWWW8rLsZ5M0jFLTlacPtHmXWeJxeLr6TQZ/59ogdGXWL05b5n
mzr4f7AMnGBDqhJOYGBsIjoPefvggggV0YKisOev/ijBhnQAdsiCbfk2KVy8kyMo
KoUTemAi5dor3JoWZNl4OHLC4L4mHBFvGrRvbKHDc80rU7pVrfPHHfDhoYSvzJWF
MqO8tcgTGoyQnNea3sK6DijeHeUauqUTk9zE9X4KF3l6pH1CwU1dw+1uZ2kFgKyW
ZYdohM+QNc/OdXT2e7Ham7cJccLJqIwVM9TOazsamXlf7IWhiTQfj06kCc/TIUBO
ObrANI6zDGDcONV+02HfY6INKL5qp+68comxBM5vqcZ0MCB8UxX/FXalegBH5AMg
OZ8StEs8Od4ilLkMNAnm4vuWX+umsrlds5CcBFbLNCD1gbkhA4t+5rPqo44okq0O
1azWLtYZuBnAu4Umrhzew5xS99ksjU2cXaEt3d2tGhOU9BqhX7En+C3WRACpflwo
0QA3L+Ie/UE1VeOYvft43wWKts0KrG8rWNWz32l1sHM92biGMmcVN9+fEfhavXTd
cetDKT4kJcNWscsgJ7W6F/cInuSNmYMAdCwg0rU8a1UKn8f2Dsorzvy7016qAGnC
bh5qOdsdXasbM+eUmLdv6eM3Uc0BXJkGrjjawj5OO2u9o2l4/632v8XqEldy23Zj
Qx5ClkqcB7sTOiYLk8ZCdP+NJZ4DP/8ogu8QEYNFjF8p1RNREq4AtB2l6TD0aQ1/
VHmMhuoCAwBs3FUhmYUXiKK/EuRCg4AAf6CLZtOdhRm7+GmX5sc3EV4PBJbqXgZL
KW5f6SlUPLT8ShzkpoBMd8qs5AgBQW78AWME4/wGjobXD2LSIkKV8NO0jDPYC1V4
ZG2h/cwRfuwql9IQVHIkS0ODUET3VA8sniy0lEtaJk9r8tGU2igW9VVf1VrBDAMl
dtGfVUDu3IIEyKeHm21/zWCqCcjpSKODQ9pDzD+UaV3E1udgM1jZRe+q0rlcPH+/
LMB4uzU02YAmBoamnBDH/OJZqiS8vpCSusDUlXPnXnDzHKzEitIJYpwyz6nXUsDj
T4/ko3EKTVgSUNoOd/DMF/SiM7k5n1eYysBZ34aFh4l8at4hlAOB6M1xIXvypn3Y
vJFF6hoMgfrXxa7o5wBgjxI0vkxrctRF8mAAU99OK5o0SYvhp7zJEtYT6fqQ2Zh5
Qx6cNG/W9IDojUZTusFeoITblUujnG+hkY6MKxXn1nb8BEx7z8ZZEkQMa7ZZFJkV
3l5FzVGEHJMS756Z8jM3K28RPQo2zSHcBaOiRbNt4sIcW15KxhI5Wnevolqm5KAE
pXGAXcspSqsU78OIuCpZV7cNZrMCxPZs28Vt/gCOlKL2h9v/Dgvy4CKudKbTQuRK
88cN1UHSxHOEIvNdxuoHjtwNHGcrtPeq6DpaxZmfpMvzotvxqP3apWI4iYcftMQd
gy8RuAV9oiMRCQ7cz7o19sjY7c/QBJ2Fz28+cIFUqZ2uLPehVLYhAJ5HVZO1mCW2
1Lwto6j+H4YUD9YUZcWH+91gItezNlKDYzKcC6tD4lMf73NoRN8NoxZkse4S3GKG
mVuDUnq28cAa9yyxRTToYFK4FVjVpoxWG6boNK9fAIL2weQdA0Ju7V+LjJQQOlkW
7FrAJSu4dJmLBXFTCS/q4OdM4fsvlmhpWRMKxl1QJNu85emRQKjFpX0ZgYcmPppx
ZskUjnf9wGXKpnTNPlZ4fYTGf7vI3mW8fKyVAIygtiSeyonIfMDFrgH91ONAZ2rB
Fm0x83NMWWm6ZqUu77maGhFmJ+MKxZpW4RtxajEXo7RnaPf6DT7bWT8304+3ISW6
uxa990ufcudZR1BOsRlsjl9VDATciqWGT8Q9WrQ4gMmGI9b/Em0QNO9umrtdcSZI
thux/nme0BhdexJwgwxhwhqIFs7hA2eUpzMP1i62Qm7e02a2/IIkJ6b3vZncfOBJ
oyCUngCIydokGV4Bx7h6FfRoPYvaRR/Ol5XpGGUpQdXjJTz+7Gkg1d9/tZ1sBjZv
nONnQ6qa3VvlUGwPdUw6QQdDTZx4WQXrBtgYCMfv06BMO9CPun2jn0uqrbvNodVG
pwewXpUfmihPToAlWdjA5XC0BDAH/jn0qPSc5yLSgQsWRC2fkX7mt94mr4/JK9fa
ZyWIXZUFRHsI6D126M8aS1EOcAUuJGu+EUpJ60YaFMm76PyoyeIeR3ktcQPU4efF
ij4WWc6U+zSwxmgXuySNI5cxpc7q/04NFwlPYYbKPpL563hC+ZmFQibADL+09yTf
avph8rzS6LYkaZ09BW1hb9bIEGV7Udyf6nyljNFLTL1bcNItcZsT2gNBvHpL7p22
cnN4oy9nwsUqLolFxwmqfnffE58NlUjpEb/SMa8axDIQka9cihrjgKB10QMMMUsB
EwnJwjveBJFV1Ds/N15wHEXdZPxRLkF0IRqfQcdXLaSk6MuWuMzBETOmF7vigp30
ykCEYbp9QMSJ6HPx/rvst+OThte17NH9Dy0bxTT+FxrBIJ9x0LPK+Jw+ztBxcOJU
RG1v1oT1XzP4wPcKxNA02qpWs+aOgQ1Q+0vOEQZHv/8oBK6kx0Vqr6X31hBnvhth
fzNmNNYTtvh7gZbsKH+4YuvEjf5txLbKzX+BhupsINYykGC+0yI7OBFOsWsd0lcq
nbvDnOIZ6glfSXd0C5TM2Y8cex/fM7vFUEfHAWpE4kiweRfL5P13AynAqFUwEJSr
BGNq3UJ69hbDDr4OqR3MYHWhn/U1ELSf8Dwuax5wu1l/TXGYBwRO13JMSTkVYe17
l+kCuuMaZ6/oEgCoDc3MSEqJX2U9/J6qCm3oTz7m7G+GFWDyrdhaxqsydIb5KC56
t1A55LXnxRhIQlDh/tZGPD5RluNESrKR9oNsjXKTyqiKG30czLTW66Qt9uIF42jS
JJaoXTtBFfiyli0lZIstjBz+HTanqkwcHSsOZgrL6KZKDqmbv3RQSOP03YhCAPU4
QUyUD05DLG5BTxMdLlaezU/X1gUwNw7IUCQy//ONeIluInpyWNjSe4zY4W0nkLXx
/J+jr2EZUqWVoimPOZx7En4r2nNw6iW42mNQpmSkPh+/95UDuToSCbg625tfMCp/
ed2cMC0cXXKRB5sSgsrLVFjeAg8qB1SWWmrO8ZypOFrRWWTFCGaP6bLjAo2YU5QL
ssb5U8qTrtAbP5VOXWgiEQTczd4GWjVxbn8E6ASkUioBK82TB/N4WaDuC9E27Wat
48/4mF3J8is1s9aHWkZ5unjgmwX3LCldCkFejZOsb+l5ybqjCu94RWHtejAWzxaN
XRohrJKJCXaukteHIEJZr9BY8ksgza/qqVHaQefd2tIw+5fd/e+MI2Vy4DFAn3js
kx+bda1dOupchUibLps9aV4MkTUInrQGpTB3/nbZ9fk44HaZ5xcZxOaIo3XGHDC8
gisZAdzEbrJv+2v/VbSlp6uZJ1fm4dq3UZCN7pZ5fpSwlkcEpG8/ZhkSb8XUjR8g
+qgS2Sqk0Nri5zcWKPTm3LWdO85FrDVesLWhqCqLgH78pQt2QjZ39k4NfjtOON+h
0u2yWjEAXw6a1rr+LWfPMPwTkuh2gY9qjYFxZQfRbx6NyKR2Y0cbpo36UTL86T4D
puvuO3Y0mXYZgnXkYA/QmP4IuFA89yVzxj7IbmP6zk3t/0pqWOhgRae68ZGJ7AQs
sz/Uyi6BgWexgSOC0PzVP5XRjDVaxb6ptPinTlMTLPK3qkShslhgBQ0A2pdFNatK
QW6+z5QzsUutuFCq5A/9d/EYMmo2YzkcOH1FifSPRwkQ3LwO2/JYZTL1OtsgeEDj
BEWK9GSx8LPdf+O6uGv17+US0s0kODqFZnenIHfGlTJKMDkD51SDOHS2XHPkf8Mh
uRFJBua+W+iFfb45o7ybvFcZKA401uQshiXdrI33mzTvq+uyJ09cUsQrvgQgeLqe
fGV90vDOvwFKUg7CHkgs1YlorzFJGwRRPSdQIbLQEmrMchzov4gvayTtk/AeR3Pe
mORMKCkWuKdpSFiEwziwUHlTnt5Z8+WUu7OSQ70KbuKnQRSqVKqD6i/oO3MentgU
Y90pnuOzf5aQkTF4wkDOxtwkT4SvpLWrMr0WSciDRCuzU7vWNKGkD//obQmng2pL
mk2K6chbDeeEmoBV99mzJBqcyDUV1emz+LRBzxSW4kcquMjjFwCYyB74mGCCSe9f
TCBkGx5GY7PiTn8l6SkxE98A/CiYP0e79wpE4ze6oO1qzv3WE5XGLrYycBaLBVu2
NicTP1Iu2X+/p6gnkslGi+X2/Wla43UqMgWGcwbCsor0XdCApYyM/jwzKgyHR4bM
mwP8JI6a25Z1qfrFIOT5g0yUUZ4PvfB1QoEzJiT7jlXNP8Q6VbipUodET5Kv7DjX
Vz+MnZLxdlYsbpEphnUZ8LVukp1ctG66quApGii4rNibLFsAktSp7vDa7oCTjV3L
/rf8UsaCjR7Rr8nWKSK1Szp8gfsfVTDwnhYtA0MLfhC3Re/JMYFhh8nUXOjtSA6y
JgF8CHaKn0RDe9WKE8JKSAxPyWyrcYbI5GgYi408iihtGPgmZwnHl5OfVWOYdjRi
mCRhPTbF6fYGAIAaMBn1ss4/4x7uTCxTy3mYIx/A6P0jktxKMk/P29UR4ccYlZny
afubXmpgH4Bc2g7lqJJmystGtbY8f9gtCMEJTw125EOiUGPeSLv+vZjU+lt0z1V1
SmgV60MwY0Z422gdx4P98GujiO797Ld3KZC3dGn1mrj4RaCV/VMxNna1nz+RIX/b
UOyvGKwBUMRY6FGeOtsmdexFU3Ipf/oXYz/Zu2/aZtD7XYCYBUtxfdu6CLV58Qa3
wlRPFeMRq+y/yVi0WDJwZAO8S8IXwG7kF1jhxk8iQl5AGP78y0r8DhrPKbrNxDfU
//glAkjRSk1satam8xK+Wtjnvqz21bKboc7QKHUKMQY149kJ15W3Oe2UFDsobajv
T2G9bPQgVGITilYOsjZJJCgj3hs0QIeoqAAoJn5T4BUqMlngnlLPY1SjqXUNusXD
9BdYdN7kuj7y6gpoO1ePzf4AWJQs/q3Cli3B1hdrzBuErHnDArfunAL++4S0xjS2
B5u+n6GlBKhAFbdwh4Hqz7u+c+Ll5JGwYIek+mD4Den0cfxpzTD5R802SJUap3Ef
H8fHDNehLidrUxjaKdSgUTyIgFs1A9WIGNNxstpYjJoIEm2OZOH1COnA9jz738vo
fJoG83a/rYTt1NiFrGeCraqoHVGrvaZfcxnng7bDOB1Jl8vbTQlZQCOHr7wV/913
RY372dpaLUXX+CT2VZALXUEtVtEtZBx6t1h+fmvRqnY0M7F1OuUn2HP5Rm/yTMkb
IGLj7uSTTEWXt/bib7k43tTxosH9o5lMCKHJ+3ivlXuoY0pr/efOQy9bI2OWv+Wn
xtaH5Ws6/ScU6HHp7EpUVaZMpoNTg7vSk0c03X72svmHEiTiOwvJLZBdvKBXd/vJ
iQEP+gcpQ7ReQ/dTRl2baRfugruJzSlYyqRINCUVOAvOUQEY5toSbylfIXP+VT05
RGkmyuggE+2piLZ4jYrxhUW50sCoTxCo1Is9XImNVw5rtH45PHPQwcev24b6Uk9C
VmTzKPz6j7Of8trUWdMMrg0NRI50LkuyQTIkIQAMIcJML9yA3w8nQDwGGDPpFnuk
CtOsZpdp/MI6l0EvBCZjDmpEm9EY41FK/kCfbctVo4Ucz9HmZYwGeIop7B9t/HyD
QovglMnEOfsHD4aEvXWwJ5x3bhSPscpff3Drz6tJxNjQXQ9ICv/qvHhiMHJdTxrS
RRAPhUrycgY/N/HNhIJFrzCTHtReoXB7PjQtfVBo2jOtxg0gmbMXEm0roYFJ2xPe
2ODdn2GiXywoTSoZ/CHobpYljfUOruPeKNLtC3FmoRRySoMg/bwW4Bne8UI5C5BZ
QRMLA10WLCPjwtlAlkAfJgExPG7PgVE+YP7btOPIWi7OCMNZ197vO3aRlDPFWeIx
Y+FdXDy8LXOhC95a4o5LnNqUrNKeEnMNXlTY217rVXPHa8wFMHOXooB2xKKYbJ4g
Zmlk+MwiOjKg/iz+j8jUqeM37wBZv3g4PQxZ3WcfCF2UNKGUbH55n7S5q0pLhBww
F2umET1c32amDdI4R/LxR2f/bClOmEVYVePF6rp/agOfuqjkMs1/f7Zk4vV/Su45
vK5TwzVO4E2L8bq82Gv1wR5Tw/1OKXXO8jrCEvqBusvLbco5PokE9UNXcre9Mrot
G41CQaaRlQuSeV41f7us8ojOFDxyAo2e9/viPCxO33gQCYdvpYf7Cq5BUBBzF03N
gOQFR3D2ST9U7FKGliXDeozU28n5HPrel22ORDcfNbkkUGHrEUoNSDPAV3F4vTg5
DI491wsIH4Y6GG8mNs8xwjdIgjLt7GCJ1HbWmnFAbsIbUj3HcbsB10htY+Sd1+aH
s+QZg9syFl6HTrQs0j2W9V0sWpORPmwZvFLEF7lMM17NnLwQQq3iTu+ER7VUS4k9
hs8LwPmhiob8n8iqBDV9cAwr5cfNvg7TzpQ7cks8Fo5Oxtjr4vyhbZohE+ysJs6T
hrfegoryS0Y7Ig/E5Nnp9MzubIQHRU/L9dlOEAPnzcgW6I/Zojv1ReRGbmICSufg
S4/mlIK9IfqtY3qD2vC6+O5rxILrFUfjZxyvdMaKF05I1PzJ/YRWlgEWbHjotkmz
drTku0HQI3mD0W+LYH3AF3iiDkdiAZKfpH0CwvKewbI9uD+xvMRsqBbL154kqqZr
ePcItxza0cCjZjr1V+0X4NowCsL4dIJlAqrmZwphTrgATiQLJHOkVUD0bXQaov8x
mg1sFWOcwGTyl3C4J8pxj/cCLbLg52BiVo0LDTDKJU+GoO7LTsaa4YG7aQ7i3QnK
UvY+R2cXfgq1F/Jg0IDIaXuwvgc905/cdlNu0CrwlkkJaqJlaPudKD6L1lxrqDU+
S6fHqOO9eNmNBuhwLnDzdMJCkXUw8wIA8+mFPv7/0rjeuYBBkF5TjiRVftUyi7Qz
ng57DN4VT6agBVL5Pp9IWd99XCoOKA1VarIQQRpG3RUgSFX1BTJ1vkKqh5wYEXja
PBn82248xttmwZK3WG7mQTYDe9cYaGttS7JpIrl2y09UxNxAgSkhA69OM9QqybnO
sxbDeofalejhvtNz/5nKUPZLYKzS+knfWJg9C33cb5QoF6y2CKo0laSQEquPoOL7
J1tYndoYp5v1+yaCkmf/cvsfrIxzaCLsM42ZJx9CjBRVQPPLurmWF6qEsiJ9JgiE
Hy/IlWv6JBSC03/hx7XDbpzv++cj0U2OqfeaQ1QObWXfX3rdfVzhTh9D6H8exAVS
sR4J7vgPmH+LjuTtAgZeOff+R4h4J79lNQIxlEx/pwrkrEa9oactdmvkn6FDJB7V
mXZ5sW37mYjAQjjxzPrT5nJZTapxW41BwTiJB7VQVLAxliRGHrWFFYx3cyc0H6NC
9S6LSYukXVujo5atdv+kImOOi3J20Uq2KSHgwPQX35kyAlGBiFRNQb8BctyVbkmJ
tZLuX7+vkBNZfWV8DLdy/VhzmTyOJzC3ZDJQ+8t2COAbsRFY1qfr6DXW5Nv13kTV
VCHxVprqBT51Je0i7QEL9SOba8vLtagYptJon3AffaBGCDJUdjFj20hToIiPC4PH
eM8bLY8MNtKG9tceveHbJBAqVb4YScQodmShf+hRV3gP5BpVxFBtO7ac2+1/891y
8JvZJ+0biOzQYX/fXz4sfDixOEFvRfpZ6yzZ8Vva9UtNMqT5dFL6tKJJpkCRjfTM
6Up2a8mTOGER8SDtRL9iWIunLhS0NvaPxQcmhYEG5/JMdExEmlLGg40dNex3N7oi
rcflIcUBBofWS2cBtGqmiPpVExNxEMlyGYMhkOKr3Gblh/r6dgQ0kvMUKc+e0lil
AFoP4+GPhfxo4+VWWY/TT5svEgf5mEMnfCY4KBlvlusqJAlaTBWf2Ao0IIJux5SA
x/BkLmPrp+1w0MVGBhrspZSG7OymyCv0CzTiF4bu+FygtBrsaQiw4aOTe5qvtgRV
hrbAPLgypQw7iEgqMcncqArunJD7CCY8JTqns0kcZvzryIZwvmvhk096HbW1Esb8
kZ07egOSBxuNjqotTKQV33dYQd2mVVABvGh0TepRHelU3W88UpFlIlAGyt7vgo8A
wxu5V9tYbtzANmvkMYdnTsm/hKVP9nGweSLia3eL1AelvuhteGQPzd5FKue7mmuq
PVkJSHG3rnG/nZVni3kf0Ta1e8vF4K2MrwaNGbtywIZAXRVMSbqcm35LpVNbpisW
+/QLlK3JOEsO/Hc7cz3vivEKxlFEJCJ3HTy63ma4hSHLFJULTo2Sd/WO7UU58eku
Ke3U2R9eZjydkd6L++iiMyfDHPJA1LtGahKPoQzARVPYk0JjktAROo+aabqcVXhM
nONTYTdvCbJWBN+Il6d4aNc4OhQRaQ0IGBDdjOYC49SyfRi/MrNs1L5Nw+NDonEf
BP0DofN0jHDdFlOvcyRTTe2FvyuoFmfPMylzUlQqxtJWjBwvWHctiuC1ByircOTn
CD5c3+lfjNoDxu8ozL9DlXMFprq5Pn97AaI8MSLwhJya4+bCtN41GF8QqbUCLaG9
PviYp5qfRVzZDArMk+EVUY3y2njVHRGvyCsPbe4ApB78dPB/KNC6BRIQZeVGGURb
4zTqkf45YVCX8Ltsayyt0cJG4Apgv4kob4xnd5ZPHCvg7QuyvWPlDYaVx8mGKI2G
qlVcRWV3aMUcZzIQGPDmPMw/UGsmNc+eXGwCt7dJaqIQ3b8SAW/br+8qp5UOxCnD
FwB3C2vFifk7xEfCB+dw56HvwKK8C2bCzhc7eapKVSWvcMf51ebwFLaKIRRlygJX
5JFcVycrGewrPSH+k/g9ksPqo2/RuTD1ufmfHGsTEfXI6csCJ4asY1mrKnc3sekx
6hVyZTPmwDyGsOmnZL1Ca5yYqxmOVgS1HPUrkdY6auD2SjpOFE3MyLh/gdFubBH4
qLI/VYU0mVgDOv/tmyKICdPz0R6XHIkWjMDFIY8lmys7TkhdqEf/bCLcvnmybNSY
8nU4WV0rRpyUTJpxqOndQBlFLsd/wNIIULBG5uG4yLOAMf4Rnzqd6lMsbLyIjk2T
f4VS1j7vAvzW+wxT8AbvmqxaOVz7HpVJ4RuulK0IpYbWsoKjM40djgCxDdoiGkTS
9XA5rlXOCSseyqMLBMsXn0B0GJIW1fWS0qEnwTFL7dZ4WwFFCPgoN7OA/0IR2iA+
7B+sDfCLPI4nzrGohLNWd30wj5sRPXFEo3ViAXe7fy5cOMfQNbpCzUoQaPKrU+Rk
ewq0sSiVHoAfR7FDcD1C4zY3CkjFJYyMAfewHmrGhebfwje8Fg4v1oRHyXKLf3vS
WVBpxeQagKYbJsf+Cs8cwiQyyaHXV+zpTjfPY//0OyE/Ympy1YoTKTuypuBRemBb
7GkYSMNpPxT5RvEWScJb5o3xMoQYG6abCIGoxNylWuYLbr8oLnElRoSpgK1inX9Q
AKkqoshw09vu0Fka6wFoGe5LGIXRGiknqWPyj2zeysC7N6dkIuKPgOPuB5PmdkM/
To50oqDVwtYhxidCS+kCgOa97mFQ9JdOVyhHssh6rOxM6B2jnA4LCGw95cRoBwfQ
9Ge/VJgMnF94IymOf/1wLId608m1L/dL4khednj9n8+XNt9yjTHwxzJW4az0X9sw
buq84kR6nD/OyfQcgrY18hLRX2edBX7MpTzlDL5ThL/ZKah6DdSGgqw5+geOWfF4
/dPC5I7BRf9W9ZIxSbLsxwMF4UDTbTc1i4vA6iZDXMvmPLXD/bUAwuVmDAQe8Egt
dtkHi28G0iIO8TmNNIwKSPcGBTWn7aMy9lBl05IkR9NxH9HruLnUCxKgJ/5U/hkQ
l90qztDq9/DH8lQSgNa5RzjB7RriW1YLAl/pm56xiZjhVi4l2dW+THoANiZheMi2
ROFkG2zmzXK89kKdJ8cVLtNxvA8vFGNvKw9SERK0a3oOSgxZqNztiNR3bQFWRe2c
yD6UJXJOM+ZstVNLsrWIsf6441AnL6AwmeqnkTJW1ajxc2IYQ/39XOx/XObv2eAX
3k4uZwgrJwlLgvRlIeOsR/+vs3CMKJl1P0dVPofePgjV5b4PKGBtWxWzqfhY8NS8
zLECrbbH8NrPa2VoqeqoD/mz6v9Tq3XhF7n674QZMongMnSkVKt+eXUvgMPj8IiE
je9Yk3BGEroUbMjd2E8DnVT9cDZqVUfStWUbrtjaxHssJPm2y2Fr0MEqYkE9Wl5o
C3o51wsJESHkKe83Pisw5U89C7b0vBD5pQoB9IOHe/s8usJBwwTt4zKO8Yy/5Vvn
5s+cID+T275DB9Jn6nqJGpjuKiIQ1lrsnCtjDwFh9e5kU89i+bdgnrr9gY5EKrZU
txU60Vinzdr1DFuIxS86LX3g7bkg9H4gK71u2iLIaMTApxpNiF4xji/3RIyO5Hcb
3W8pezSU/wwLOGwzvxh5+ga3krlOLzavJtKsAyvCnC/myTgfDomDOrfrfUuDOmUU
DPjxHgHqnpIV5AKjdKTVI2V4YQaA6HaFqywXr+/7zydiUs45qEbEZDQl6ZBNPi2/
aoHBnK6xRcqzAGDBuVZx8gVEZzCKGtCDFmLc0dBFz6uaG3PnrpNXUhzlbbBJfno1
UO9GdVuZzQkG828nWk0h8oC8V9oHsiCv2xoVoWtdbsir2ltPcnRmKwoo2W8+NtC8
eEbRR0iS4SPKO4l3bhAalycl2xLlVUGKDYQaeBqDgbi6Ige4G0E7/M1IjN8dWYEh
Ig/2tRb+STjcCcerncx2GfYNjH67b2QCl3ZfRTkrHXZpYkmtItGIrBLgvo5woCc2
zuJl/bGb6dN63vZZvNa/CYTfKiRwrr3809rTz0O2NtAgoprl6+SEGBbObVa406x7
o0nzXYOmn+8yICfGTqC3fYqGJG0MxeCHt5rYgoqTCY1VKtkHeH9kyU8XhNQQZF49
3WfGsVIsAQ3oPfZvOMzUFpEtEUHs98SOybs7rSQQCPopXcx8NYb3pv5uDezlNyqV
acT+72EDuIgBcvTdf6zcWw6Dt7AOtuvV3Z72k6pqtAMLESzS3CgDd5+5QPYXwA+k
zJ8whJe6zIyjWTzH15JF+TdltmbTBoQg++cw/e6tbbs29sTrF/5gEcU7yzh0J7K5
rBLZqRyYNDUmhJzCETIxOcQcTAKwPl4a71ioRMlSh8YAzG2L1Eg9zfzX8d7L3FTQ
/eKtYpXRExL4jL/E7tINkpawUF3mnHKN0gvI7t/l63SMsbkYICCEolMr/gnf9vzu
NSgx+Et5uXpJstPennuliO5Y3tWCWkUiSN3X3wQHuLR7r2L7OEI4W1cn5lEujtyu
QMfOTR/h3Bwec+rhj+MCqyjDQHNNGDkMOOrtUcIP5+sVPGCf6UBTpTmXirnTY04k
OdgfdzFC6TRYkWA7wsBK4JKMIN1VIQI0sogISlge1KqdFCcjq3Q9b2tEKNCtysi5
EYmBzSrXGIdrJnmK9Ozsnkiz0iIYkideARBjtvOBXSJXVSqAK4F605aEVcLw4D3j
wSO64xVXOcxC9VfargByOptRjo07Vr6gJsY6WYigIHgPZG2xDMtLocAXfnh9LBSS
6iYchy4MXzEGAxjk5tuAPN9ygqROQJt0LuOybqdHuSbcU6iq+LNQ1mEbLMvZ6A/s
ga/kcramFMQcrBb+E59gu2ZlqeluoDPZEhRddVJI2MNjtA3fMsoTlnDbtVhmZehk
1iOX3GeQPrIJJINvvBDmlvqQyz+v6+Mi67wlcNE/YGJg5B2hXcNeWEWWB8YmdXRr
K+5FALx6VqdoogWMl+PrNSr3XDWKBWGzW3MMt0NeEsa9RD/JA2EVaVvtV51FOiTX
5FH45E3pmqslqZleyxqkj0UGTyeBU6AG87xK8LVkT+eEx54Oi95kADpX95tK8KDP
MFaxKtxJMC845KB8+/RGEjHV98R/W2r6ZlaIeexDrdi6jrxTxZQs/yXJiskmtRNw
ICeu8kKxSiMerukXUdSvv/UVc7Fen4WIejGehl6JQSvP2x4q6XaYM8jdV4YQ4Fxr
IYlKBrzNj0P0ytYxhhoLjpNMJH4ND8gka6zxrAWssz1Y3+vyJNsXx9O+7gj5CmX3
t/uNylCB9Uhos+BghjOeJYgaJmhuyNPzernXiFtd2Zjgsveo2KdZUBeaPD7GvFA2
TFBWFSnlhlACAzwjlvL3bXBmO1KnmlkuP7EjXK+qtvnMqJhZV3EP4deTj3RSY5WX
Q+zn85ZFSbC78U5QEcUzEH1hKnOsJdEAqck9TKEaNL98pr23hZjSNhI5CN9HFAbE
W3Vz7Zr0f4aD8LmgBV4OvWQpXmyFF3IgZVNnLzVEG+GcKb3x9/TyujtFGvRigwov
7FZebsLhR0HoFHXKdcpgB2k+kLcPcKDTt6+gOHasBTIa8zN/GSY5+CJNpnhUgf8K
bCcqzJX5zFjENSeVHpLXCtWkGD0QLBr6cCjJ7w2dXHB7IYS7WYWd8BeIcy3eUklQ
XqPIE189eYh/RPbt5QDXrZMKb+6JLled3TGX9MiDq4eDRbAuhZNvyXKsykfvNjSM
7QCEoQLDVIBJKy0rMWbNSAaNdOmZ2b261g6ZJ81uxpLpR0B2nq0NuWNs6etWbgUK
twqBdOMRoAG+HXJ9BQAgwudN0mZMhqNbmiDKw3OXTG1dbWRwju3FXC2auBlxA3qQ
N+6E7EwUE8WhN7ei1ZSmep27S5zYTolXKQQWlDelF3yB83BYLY1pVdQ646NEUSjp
X9MdcmuadDFhnBtDllxoMoGVBK4GIeCI33jrNBbUDTbi/lctUE9d5CRMiGlsLETv
jO2eNCo75Ay+ZYIOlSm+8cBpYPiwFXvxZIcudRTiOmKdeqKb2+I79RG+WKS/CMrm
vMGDxExdaXNvg4XbD1k7nROnUSCZEjNW1K40aCBT9Ua+TbVPtUfjq6vBp0WgIhxN
FLI2rfSdGEl/3TVz8OxmFENnnEKMsVpBw6Y5HxkANKEH9RTdlV79PBwRjCsaL9eG
4ngijm4Du6JE3EK7dPcsK6YS4WYHbTb+Qt+cZWYVxbxkMOkXgiMfcVEX2hhkAcIQ
Zk8w4LUbyfKIQyXbXDEENla9EkWRjD7EPOAbeDGePB7hG74ArPWLnv+uhZOzC7ax
FwtBloNOFWAYw1xOaO15OdRadoyao0AMboac8WTi40vHXTobPHE3okB+hQPkCm1S
nb0MIUIJwD7Z1Mxepc/yBKQo08BWyulJMF4Urh2SX9+YXuF8M+ev3jLxRWvZC5K4
n9mmGxkOjw0IImZAU1eiKgHcPetkKXU+pOKFX+wLNe5FLP5JrQGmGSlnxQP0ultq
H4vNyJEORGKOOH5+2mfkEQgyHBTorlcKhALyDufgmTG2iWQ31O9w7+0oj6IQdrms
oJJaGTToKv3cDTTIw5EwPvjWd+1/+W70t2jHYMgvmgEJzu4aXzUaiXbBSy5WrcfP
TFVy1Nwbv4G1A4P2LExss1u3x1rCkUbggUR2yjhrfj/qPw2F4tfNzs7u+lzoKb4x
z7q/nAWdeDlJ49yyEF7FTn3RmgwhChaUo6KQsz2Yb6kKliFWsYavefyyNX/YzTaZ
HfrVinjNDIlMVoov+/1JULXQvvZJ/jA4eA/IiVVBRC4NhWfUk7TOlUVeaoIWvvZ8
gglD58weFnzy3wx9nKMwR4FuZx7WxCDpkQnojcLdONbrD7bZoZZzQ0V6PhMYz6lA
cJzgwhciInvpPUxyg7zDK5fAqFicCNsRwy/2MNFDZSlQv65NBZQI0WBqncgXwOex
oGV8XZBfaDTjGd0/b+l5V0e3nacE/rcEZnSlIyOzdONOc6uRTKRWcmsCB1h4h1Sf
p2JjX219ONidHnZfAxdpsrCQ9cbzLvHhPVVF96RcZkoku59Mc0V3wDUYh+NlVa3t
J1p94m8u65Dpg81UNheoo/E3hsxmaxZDo2GOPYJ/S5rgyxEjVGFpYyIo00I9Iwwr
KqCojVqaTO7ngi5OLsQ8YzqUxIrRxGZPlRKw+mwWeNDR7NXIhpDXEfbsehAi9wM3
71F93ro282aYrLwiQMQA1aKMBJq7A2cag70PCmviKirA+wkRFszhvhhcX5gCVBne
oazAHDpLdbsR1ILeXfFPo3jHNhfajpcbAu5q0AyU3e1E5C4CIi6YACug3AApIC5s
2mY9DZYfLA3cmJHkYsjqVHarf1c8uFqRTRSfJf8DKlc3rsfjxiM/z3oKg4+M80+Q
L5IhYMS1yghgVVhAw8ibSoCTLaZxSxLrXD1uLr5Fs5kYbBC8wk85a8DBraK35WXb
V++83Bd3RmtWt74SvTt19YGHgbG+/RmKFozG53zjnwW/IQFIEtY9b8qapHGtjErb
cOT/HIFieQsN6utgRZdKfomHSf6fnJNVVVI1iz47ZFbCeA8LjQBcY0ZNiS8RnItB
IWPDrZF4/uaicO5B4cTc/9JbTkEUXrqX9w7PqY7dWWZm3T94qTdEBaeEd3YcmA4j
7ep51q+a5xFhZgiEVGCqjD8tLHawdifM4bXsBuRTjZkTwGQI2rJ3068znNPj4Yd9
tPtQstKjwwhAtO6OHw9nUdBK/lnDBSIUrDXc3hwpSnj2H55eqqz+aveU0KSX5GxM
S25Ohmu7AQqNeWrUEKMMn3Od1MSS7VLYyxc1KEMDKj+bVEZTJNayuHT+07P6Xj+B
YIFa8WZ/+hLHEBylRaBzdqwsb692GDJX1o9UtHz3NGGPnnaXarlqFfInhvk6ceZ8
qyxqy9TRAOPPeXkKJeZRtgkkc2Nr0qIvV0+EXRV6aMT+nSBZT3g57YDVFwfokfYW
azcPlnCYJnlIJ2RuHODocKXAWHfRYU/aCEmXp2TMMYgXRLJdp63fy4PS+ZtUNxZ9
TwZUZ8iB795JjDLWn511TCbfLrpSDCKQhtU/eD9XLpGJSWcX5PNEca9rBWwANRUQ
8yFRV7skWeBkq6pPVDZtEqB9dkEfnU1DdNzJnAxc0myWGlrKerjr/24Gbl0n+ZnQ
3v0kCBvTnn51roqI+8LIwJevwD/n7Df1tVLHz7OjSbkRAUFXNdHiPf52gAJloaZ/
ZTip2/OMPT56qnpxxhPBVpeMHSEfwmvprRqGnZIIxTMMkabKYAnZEC2hzI4/Twq7
zystDJifnRRrUgyymrpvnGwwUa95W1/TUM2eDoEpLEi+YjDXdBm4zz2fFdfi2AO1
Zd3qQ40DMFr3SAztsHaL3eSBRF/rmSfigZF6JgkORiq/4jE8qWX4rVU9fcYkkuqz
/PPFtUiNvsXpz46MTh9NRcn5x2Z6NUcZzVbj8C19QFrjJ8SuVeAKuiK/EbyamsGS
sC4YzxvxC9b2JpwccpLH1JfpCfVQPzhGMO27R/rK5ABnZGHntR+XaJaHPXSFg88q
SBwM0yJlpx83SEbHsrwpr/KnNPL7uAmT3qBkqE4OtVsmPyRIOQaJgoF23+wYq7p2
XKk57SmYkkNzUkao1Gf95nVQVHrvoTVQfFPrifPDswX9AHzEjpeGZWtPsgXlZ7a0
Verc4c30s1+F3Lvqo6NwxTJVazIt+KwH+N6+n8kOxKpn73CpSQmH5wjmwotjMSG1
HURmK+lXJw0yacXtnX0Fg0AtweHwv/yU6s8U3AG7D3onYl+IcH6Fkdx4lCJuF1aE
pGfMuhzbTUcdm8EOH6opwoX1ClJfQ73t/fLIBe9G8vHk3qM1RB2EXqAtnrAKhfyr
OVcMw3jz+Bf3+Je3hBVE29IWfMG4HyPpzolCjcxA1E7YUwG/H5xKG9by1QG+qtLn
MgeKix8BllwV6ViYBPekWorLCEXhD0rzRl5OQ68yHpI5AcdycZqcrkm4E76pvYV8
HAtFIlC1hgnq3hhGLPt5JF876gBxtjAcpt7jbWBESRNiAPi6RGmZIbZGZVmzN5xx
NZsj8G528BufCKSg+m8IGzZQA2utS7HQK7mEA9CHV/smZGwRlYrQPRgRoJ4Xeixy
BVaTQS1VJfqRrOoO1u0zI3Uhyb08YiOj+YmuZTPHxU0/PSNd21gkOKnHQ5duc4qp
vuoSaO/oA6v0REYVFk1DBA5D54O6uJNNuGqx7WSur5RguP0FiYsqjxS3W7QOb5PL
C4s6Mkg2CaSxpMp0PoT1PfK3x5TG/UWrSqXhpK4q8iqz6NtXTFhFPx75aatcvgIJ
B5OfAK2KoIisL3AFOrBjtvWq725BQH+e7C5E5zwuUIYwBn8SyMWnUYVWe/V30O4x
5FKJu5WxxBad0nGr+Wq9PmE5rgTyatWb11OoSILn00VY5H1jYqwqnuz9PXTIEX4i
4FNAOA4hA8PQVjeM1wqJEV1ObNmsqi+nvx3tvwIF9BoTTgP30ZTqMqgEMV3W8wgY
VMPxxxKKZyv6Eu6XVNPz+vpElM1XH7GKLV9tMqeqxnp6GENo3GH0DzUDQTK8f+VO
dIFJBu/MzNiqVQvMZU5NY2S16MaaeQarGAG/uxVR5s6797Stfoz9h2r4+gwK4C1O
FIrfl0QhRMPTgg21iAyfdLDcOJo2jugEiC6PQjCIK01x5DoJfc8RAGZr+FAUFwL3
w3qekHsdYmAu1vPPAXj8H/v0ZqNISpBijMJfsRLLqbi2fsmj9vWTqIl0pW0mfUYD
UG2A1u5gWf+HGp6U181VDW11VtNZK9YDjuHZh+7jV0tEAuV1L1dUXUTzEO/ctH5B
EoM6R1ybTEfsYRxt17+R5YXRbBXiY1WYztwKE2cGI1pYwsP/r4qP5+XMwW1F0eai
TngzwZvi+DCrKcAbm34Ogg4oxIAJcLSTqFjjJ62nxG9QAvP0pfW9Gz10+zX0PcGF
hrL8RjOwD9T5TenYZQdRilpPXKyvGv2687nct5OYw624eNaPvgdDO0XRwPAut/3U
EdjOoQU5zSZ0fSAzL7fsQRMGp+hGInbBuzwOK9JEkWG81mjswE4rp5sMlVc7k8MJ
He/T6Q0h9NKJpzJomeUGhMOj+DibuAR/dmoC8ZLLMNB7iJ7N6ik2XrulVBiGXzsh
qI/nev/+s4/nFsv6PxhkEGygWgeCd/KOwQHqtMYiQ8z8VKl+aZqhnjb6B9ISvtbM
ea2NGs5uiIKvWlz46jAAz5oYl6Vljrc7vI2V52aj5jyeGzHuRTDSC4VOSYkdifGx
kVle2TrmtKPNYCaRRQqc/hFNOdt6+UD/9hV33EtCgENGBTaZ97KTHV+f36fhjDM4
KI8QX8uXIHySBO0+mSaWU/VFiY9JjaSMpZfAwXmwHIFfHD8ppi12loIKTuSGqAcL
kCr+fgpNde8hlYeO4gBGkIsNskC0cWP9+GRYbR3qH5bRtHwPIRW+ycS1DjaH/TGx
uOpebgI+R4uSiqIN3TzIUU5tGyrlZdnVcGQwHmTwtazGzywyf5rXe/NqTechlOQk
xjhVHq7/CT8J7ikiCjvpOrI5NIz7o6aSJlRKLGXSISTPj0klcX1b+DqPUBdTLpf/
bCNty/ptjBdQOoeKyapiBoLamEI5L2RyohULElbB9z+gNPwErqgexBG4N5EEecbg
8k51q9jwLdriwb0WdB6hd0Oo/WoOOx2CVgaLNKYwnLm0aySmOTrDG3GSEyC+Y6WF
ka6DJ9RAEY8sEfnblwJl0hjVn/IVk3VrF7RUXbNg8CVtKKsBGar3ObwmLtUhdR+3
lcSlFA2gSa0slSAaShTs/XhkZEy3XPkMVadp3/78HgACIChlK+b+SQ1Bgyvthe4x
Wj8iSuX2pKMXWxdoPYMwY6UYBn3MlfMiz/fmgXpFjesojof2HgHzmMD3MRQHEDqg
nD7lLzcNKultWiLG0t0ae3vcHGng7S2TPTLuWd5RVimaoBf1xQEsW8ZuI2lnGRGd
QqK/OjCsqFgQCmkr+CIf+ovOXbf5XvUTqlRRnLBKDrJ3vyseoLRyJ0Q4ewvQiNYK
auQ/mLzrXNFjS686TaX2rldcUZNNq6QfR7bQklPCljLKRCGBkZ17yukbRQ80Ll5Y
Efg2LTaD7mtRsrbsWAaJSpy/4By7f+6CPM9ai2yuBvLM5dQH43i0uMeFYB8q0rcz
ZvVW/k75xUS5ssiIXg9joqBP7/zqJPt9fLxa5yvo5TeuTbfNIPETr2UGkCXwRceS
Xv+090AahdKlD2g8BBWfqd55tqadZKh7r8VK4lIegyPHpJXmULtndXRhEG31dUOs
D+VY4CfvoAp4BU/gLx7TE1AAp8Mw9KhYwA57a6O+/ZonDdSjEH47vWzuZavCEov6
55NKBJNqCQF4GSGy4f7b7EsTnuwlcclcuZB4a0w1JyCn2HBEmEyLyov3POcnW9zY
jYlnW9Ku92FyH09f/rtbMRtOaAvtvfwzNvCqny3dqd8ZZJaA/aEJX9+LpHTBUbyC
uxtj70TIwc5zNReA4j3n2CFJHoweG55dihHp112NW1jP9XT73cET6Jgn85a81oiQ
vpT/0uD6nF1w+HOHRG3CeugOEoqCFI1sbsdaruThCOcy1FCQJrRVqlQv4lTg+a60
Ub9DppgKvR08+GyXhdieNidKx0yA+7L0nQhbmdl0+Nzl0MlCKdoLJxaITcPBVPyO
PRaL+9AshgOiDLTruIk5D9NCr9ewhbDTLzSN4J6jVBMgs5zeeTaw4hJ240d5jD14
tIcHfZptdJ5w3vwOHI0Bn7SGmOZuPSZJR+ops7FJwy53eoHHXvVKTvDqNXKocqgt
poc5e4o1Mg82GbVXNQqdaligwCFGDYZEjug9PrlZqRHE+49c0WWGqebvI3Fto4H4
6SqgoBrqkg7Rgn/UGcudrcjfL4wlY54q8FMQc0+vCS2PWSDafuRYpnK2EFoTWH0H
FMNUETBzcv73/A5rswQGaGGAMKUSQn+/KaV6DnRVKwNOjcu+jvVXrtd/4X3nJ9YN
7f+s0KGO6IJujyO6Io/zt988ybDWEdRlZJ5dzR5PGq4uLugvWz0+3vaBuUkKboFb
VGsx1LBmXJMTd3ypYdRkHBal6+YhWG2cIlRlbkSk6kpZjf2z+LpHzLJl1svKg6it
xSj8A1XRr34hKATcx7qz4A5KYzTNIQG5kru0Uuvq8CucuCGbn4UtvKLk/CO3XUiI
4XQKjljmek+NRSMQms965n6HtnS+JvZSigbEX+/Z7h8WI+F7TYVjIcjmJTsj5s9n
S2ExYzt/T42g2rgywE9RJQHCErLlxMU8fynDQT2fzhVU6rTMI0sjeAVXhZOFPRFP
EUQXcKNip0iQzpzJxoWKiTKY7JJpmfm64eW9dImjbFDfVQ79qw0kJXL5UlwXmEk4
qjx0EBO/uvyMOeII+UWOLe0Xo/W0LnykxR7CDg0reLO/WEbIB3iDBxgvIIZdVI6k
O5G1zgX344KDhqJYB/iEWrEo2fD4sGrP0pLxVfwTLZpioZSKhE+nuOpFmofUrRbw
CxSsvD+Qcbbpu4mlelnOrtHNFcuA2VefRRGEWBkt2jezkdGz0HxADqFRw+TY7BWf
xExVdvQzsOG8xwHuNdjVlIZ0bjKslhNTHw7+ysPxA16gPmkaK37Fc9EhfpbGamha
BsQXjhm+wo983tqqKfwQYwV+wXeEdltcpQuYFlPhjkDPD/csckHQS1KuOOWGzfJY
YQM/VVbk5SRaBb7ex+zmbLN1stRAcKiBBt+T7hu4ixZIxKcgN+636PjPJuOsjAYw
g3DvT99OO0jCqRiOrtXD15d492+Cncw52sN+ZvPJR9wuxzO/du768n7lph3lY6YS
1X3KERxP4uOZxpBIQIy1MjJpEIz+X4qucEWRsvRl/95NmnbA65compKFuFzmV6fQ
1NeC5lqDLa+7OMBOpqluDkRIeObBEMlzsGA6FjMTeLwqZxi3zgam5wB7eTORdk6H
1RwaFfEmHYVs+k0nYVfZtZlHQ//D+GhwJpXHGOy9j8Ox1WfLnGR/e5ivkOUwLDu2
kI0E2cp8S1STgh6XCniip599UwxbOggQzbrSMqsINOO7prZcwPO/2e3Hli3p6vBt
D/NhFx1JYZ7R3LFUhk02OkKvSsZVP+itvpIORxr5bjCp6LAmQzK5WWlBqwxm0ElQ
4AT0zfU+t1pCBVtMDs7c13a6LKKfJQS7vwd5Cd45bg1YYTDG80j4/bQV3/WBKqJZ
4kOZMBBJTRvVQRFr74P8yMwq+ByUpiJoAotD3rbU7qmNODAu7Dg2sJqZJOKMbHLq
ye4YCK9MM161VRxa2PFvGOhVwRGM2aIiUZnfzEiRZuOa6iOe/i5p3kSzyEB+wvKI
oY56zBSV+p+1XmLlO+G+rXOduCmAULHodQiujxDfY/3RoiWRTtVXy2Sgmt1b8ZsU
HhhtCSC7p5fUtUoe3u+m2DNN4NuE/KLWsuVj6zOVfPnxUjQD7siCPExK5qENvlLi
3z+prhbWxpJ3tmKqiQ40Shb0SQznOzCdthiku2/zsyKdycojSTXVJBHuOJoqVUgr
KJ7J6pxyUuv0BjHbo8B8/AklYTDA0u6D/57yWQwx8BLZwemDiQyMBJq1A7yQykyI
jqzJ/UPepCSLAYYFoA+RPeEeruZ08Ugd9CcaL5Tg3KEAKjdy3aGAM4eZoVHgbfl6
7DuFG6OJ7Put4tCMBTSfLoSBcAFqpPL4h/lW7PJWRekpUPiLnp58pabCFf6CXG3t
PAbhxIEQAkzOP5C9dMcAF0wKeSNiRfYAXv9uLmLcJUHbII9G30dmrLCyCC+XIYYs
N5EDeoZsPaLS0ihIN+qmncDLxqqmQCFTtXclE8DyjreL6r1OILQbX6zRUcPNKotb
+8+jY7kRSe5IfVzCyRR9RWGHUDZ/CcmNHXXOWAg+75syaK0EsH+lie3XurhdNpvr
pdHuAJ1KmNW+qPSzluW5WP8S1cm+o8yf9IPU1yP4UiQCVegel/x3ulO+NR5X037i
CxhpKnKEjgrl6clOrFc0Q7PiUKjWu353qQxsgmsSzY/79n3//le8C0A2WXs47j3q
q62ohqjzKqf3T5YuEuODHb4UIzGk+FZOnNunVLCB2xtdfZwU05nb+r/1PO4JYUio
zLy0piPGjIvy6ejmXt1b8ugyO2DzDtZ14ZoWLCJyr1dDTUVYBCfZddqUkLACVlGV
vOm5p66l+vMgUl+X0Xu9yYulKzrOEyia1lGUF0EKp/LPIF4r9DD/V2D4PFqyL8f0
o3cEio1jYpaE1GWAshIRakc9VaolJNy4MmZLBC2vNQNvEoE2ZKStEgWqgQfjoFmR
3PuSU/DchOl8euKcCQtDIsWCXxjUSxjm9onmpujEnsmiz2mRuzWzzhGbl//2rdL8
TKiVdRAjzhseRLQ/JjXUoTqxZ+gsW2qYMlbO951RwBFvDKXaMiX6l2JEq2duIugg
xeoWVHHHGB8dT3JzqH+VwhRi3DN92AeiHurXx3IDe17ontRnF77oqgIBcOR5fZsZ
sr5S9oIf1Ak3UWBGZBuWRwDDfxPTKy88HeIUajEpKDNn+jc4oWVMacSfSTCyYFJM
jlHa9L9Rm+bInPhGQzdeatGHWDeOCkFt5yQv8J8qf+Ixa7mo0wj9LjiNloxD9/Ty
iFlo8VpvCPxm/2LbUAeQn5u4fu7fF9g+h+jmxKts5EdYHErlNBvJ2p9BuKGReoFV
KYLMclDKaoMnLV6fVTrJF1t8qWgf1uRhKg0tmaMEEVTg7tCbu8NvFVOE/kB5U0nS
tZ/9ehoMCsSucOnE5v1qvW0/jqexFQYMdGMhQjzZoC1yoRU0vjSnSUd5JI8YtcYI
uIUZQA92j1cuotgHiM8sna0tRnkMik5Gpd78FpMBsYss6d4Ci+9yfS46JjPT0DLJ
3mIobTPW+kjXBKiCPWn202JORic/ldoEVMG6dvoZJGRSaQK9Z23/iVP7oRux/B4L
jviajbEQZ8dkGfIWmWghxs+M0JA7gDGONT3LM0dvP3sRmQHz7yVWhcLhopIDMOjp
QWXrosH6iOgNwVmCeQ/zE1ddkFJSN5kwkJUQ8ebIxhzHCE3pXoifUsr1DnNOMCRd
7OMrrtbGw5Mzuo+ptAR6cEXF9vcY3eqYQaXcef5IIlXR6KcZkrJY+nc/1aTdNraf
vQXr4eytVidwXr2h6Oec9yE4FWNCCgOLYKjTyZFQ1VysDx1fKCTYdZ2igP54xh1K
YSKxTOrGK2jmE4pwHKiY0ufStrnUYzqdpRQWjnfSIIqdhjEH6XCisIN+uDhG1mFP
Glul8HPFct2n5PZ6cvo1U4yI841tOKVZFQXuJDaVc9mmgwhdnfXtES7yp0I7UZ6i
Y3TYye7ngsLeyNklFGMyzCxQlOk90he6HV5huYv3DHRcaqZQbLrOYZU2mg0Ginl5
At/92BzqbqjS/QH3HTfaYOpTTentZYMRLH7T1qc9fth56s3/uoLwsScv5c0YdgxV
qC7OWSqHhgOhabkbwYs4VPXYNlAlU6ka0AbE+es2mCDxnqbrJZmaiAKF1yffSV03
H6jVsAb+iMYLA12LL5LYj1q4PTtqXx4Ps0/WaBNh57N4snEqtulgvsu396IthA/w
QvfFVB4vAJvZPVYSRd7gh9PEv6pmKIxij1DBU1Lsgdj4RQT4c55m5CwQolln7b07
U6+H8euTxMXsZ1GfTZzeEbwpdUxPHs7W34bm1vFzz7bIrQyigMG9BhF/oLhe75cB
3RwPeKN/dCRLbRO7tqP9DhqnSgaeNxcz4RgV6n4X1cnko69swXmoCUQeW4vRSPJK
BzeNEVMKxnQ/Pg54bf7k54Snxqn6c6IVoyQhl2+g+hvzV1Hu2rlKW1nz+tq4KInC
99CjrBHr6QvJf9oTrVTNYbDum4xAn5SjOp7MSFpKeKicj/w8ffCfPRxS4ibVfbSp
kjtY6NlVhy3DAg8rtgvsD/V1nAfOB02YsVVSbC8t6MmLrBlYJA5IseWohTvm5X/e
BRy2yI4J6HgS8cecXo7LP4x2RrUe12XIvnRcyAQ98vvYWbva8ToGSRkPi2hi1xS/
uN0RnnAjknYnWARHY/RlIXqx1ooUJqOu0dwWc+uSN+sOLfwMwCfr/2PJSQMDCOvD
/RQuhO/To/XANedoTm9UPEkVfRkluKUEPa0D26i99skWpglS7RH/suhKiMP44rVU
FeFCQTT8Oo5vpoddG/0ju7TKbra73byHxe1zK6cZhYSsz3T7MOIOZvK73lLVGm3f
e9Cuka1uPW8a8SN/fJlSwbaU8kGXD47MygmLoaiARi2b4hAQ3D0vFT+S4VHX1i8M
QT3ameWIJUPtOLe/dkmHtzO/yzxlddkL6Iy6m6wuJl/1KOyf+kzuaCCqJmH18gIQ
qovIw1vnLdw91O/k91BApDv3S+NR/BXy/DVSoS0sgT+PIHUc0rvPI5/urfD3vl3A
3wAeNyNTEdMd5BNRm/t2ffxz4Hy72JMqQgS3IjT9AL/vI0tno29DI0zBPhS3V6hG
iQeEXzcZHXXpfI62LZoAH8m7KbJqQI/mDFWXtbFgldPrS3wv1huHhDueQIbcNRx9
4FeJnp5TgoU+BbNtxv7PlJtIgg+j4eVpif0+IXAg1dwQuD7ZaYbHeRew0JTHwWuN
SUi1kBPfwa3B/Yh5Cfm/Y0/g6eMVn/SUTXU/tW3VM6o0oGEjL3+K6UPKrpnzEST9
ldF4vtLrBWn2rvbrCazB1SxUP5h8tOuPiFE93PcWMPr144J3UuU/bKsja4Sic8xt
mPPRClrVKBRGuhV53/6bdcdQ+QJOXPEErI1ZA/wVbIvS3lqi9YifGjWZWsOtcs1L
+607r4cUN3mncvhsoqeA0+SUY7hc/Wt3GxcwiaBiH94hj649PiFiSvt6z+vVz0XI
kQJDe4yTbV4/71tHMNwsu8WWeUCiwVxt+N2lollTXLjHvTxgqQDxTlp1X8lHl9jr
5j5BcN4fVWkQU719+330f0vejVxuLuH2eyRdrTTQMcyRSHX3uHC1EKKnkPmWTpWx
i07grqqgPef0YXC+cS7SkiL1L64KvQ5K4lw0q51lA/BMwmqn5ZwUVzsQ0DxPFdYe
l6J3WCjR5TKn7nnI6zMK8wzaBII1i6ROM1vZNXMbr8tr0Ozry7oT8edgvh9YnR5c
o2ayosOr0F3w5SM8pSlSVs7VdebItkbtgL/Fd3YPoDNNPL6JBMWmRHN5CB06vTgR
RL21QrYo+Tuyde+dLoOIona9Cqp8dev9zOYH+rsjXyMmZnHPWli8/JaERVkAfn1U
QtM32ThTlSDBEOTTpPiiOZmDVA/ZrakbSYHFY0m9FfEBomgUmnUwdD97ECSmWbgk
cvabGnaoomXQyCvt0nanAk7ffWQCXyZfnmQ6dCYBSFApyJrPmqzHWX6uzPGgZegJ
W/FU5HrBmJhxBa23g6KXiR6tphesmHHat/BhxxN4oJOJCvi6YJlmoQQy2p6h5q7Z
ul6sR++ef0z+F6h4dTFMBiSSPmg9vSKocZq4KeWPIwdDmjGxeGrYEMivA6Bgphsh
nZNZQbiOGwYPyTvUzfHpkmJIOljyr+9p2vvmR484FGpi/jdiCNRzjreq2qA4vSGP
b/OLbi+3kUMpfpfCcV6voA==
`pragma protect end_protected
