// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:40:21 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aLDz9bvvjaTU7BKAx015+8JXCzx3J97vHiHO4gqmdpWD7vwjDbZnq10m5e90zCx0
CgLdYZwc6n3Tt61o4qAIcC5kxvdP6Pl7kXjMEmo7Nt4ZV78OdmkTC3RC5+27+ypa
Rhlv5/xgJBqLBUChsnvgpVc43VGm6M9/Y4feioAMaTw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21920)
VKui042KHE4WQYfwSPyLr1XDhT5VMVx4Wgfydu6PZCl62gw3ruxhw8wsLBc6IVHI
3ep4HsaiHzLgiB0JpeAx/S2C/ZTVrtmP5cjwf/iI2SW2eZfWS1ZiEjouhqBxlXuD
4xUuAR+HYQ7pGk7oPoeHldSiayx0tWw54XIg+Mjvt5StlrbzNhT+cCGOoqwj5Aud
peK1R5LWsRWNUfRTBAktpJQtx9z9s30UlCIQqR0dWJztbRxJ+7a1qs+z/Ix5SmLn
2EwCOAec5/mUgqXRSsG3Z/YKKbP6nHeXUFB56eViVKNmHk7Hu0mVv4l9xuzNTWbU
QID9YnSQVTtwKLiat6EEvZT7MsFZ7YCsyrp+GvGO2salTgzJiOC+emAJTmVdqf9q
AuJb3VD6+kqGkAZFa84txK2kYpS5WvAGd1hgWNDh3PJJtTxnlwsBYCkQdPnfLsGU
nMFSkKSSlhExW3M31uyJucST5PeMucROitzvY+UC/KZaHpZEC0vYTjJNgdk73/T8
7GL4+qceAWef+LwdrhAb6SiDtMYy3+BcgwqixqTjfrYrq3OH/Lpm3OxEjsZ78Zms
3l4yFAymdrltHdGhY6/L3FoQK993M6Gr5OJTbRnYejzKwqt1QOiheIiDkCPWPil5
sY8/k1tKl/PKzdvVPEvgWhHrCM8KhClXTQemuxty57QTTZ/+mSWl8Vd8ldQRKI6z
HeymIiLrNtpSoZQEvuCWGnjk8DCTe4NYoSsv4eNfztiWLYbWqULbSoKBeUvwyp5y
ISyd0dSsIWHyuldDnkzKWnGdy/Pc9uvcPj2NXQOwtr1AVreHqylDQsr9GxFcj2jk
Z8uJAYivJRwZSsvvkv/eoPWDzz2yQy5KzOisU7IWpQvjyKWzODuPxnHF0EL8eN39
E9wis52IEsBIlAEdY8LBoy9vxDmQM03OgdPaujRk9GyGCh3fRgDjfR9MUsAsWocW
O8QPXVGXv6VCoJZR1NazFbsUEXNzsZmca34GEUXpgV9zdOMmQ+JgVKx4OkJhRBgK
R15+cD19mcdAO28vT7LqOq7TxJ4lCDI7tr6eufhDUJ1OSZqjiYx9ppQdc4fy3rue
r8sPkUe2ce9t7ynzIk2HJi3naXDfX9wYHO09iHA114DyLo/5CtEBRw7PicNW62o+
kX8yPM9A+vWVfBRP3lkbZvwkPqGA872ovCbA+r0JsoWa8mOn38Q7vStB/E154FvA
NL2wPfz+DGeE8YQn8o1k9nGx1Qp5KEnR6n22GbuOB2zVS3EYaEFsSeXAZ6GvPHi3
/REYYeABlrLTsIjL0OG8dunjSVB7SNT/W6RCYnuYC/4Vi5ufzcelxxkV7vv1dadU
7E/7u4JVNcygJPlZvhP1i+SM7foFJuXnf99yJEFGT0C7iWBdF8MBAkQGUvEB8aZz
stTI7WxmUU2ERmZoAuYzXNDKzu9Jxi3a0TCmHm8OrcPCB+zXV+ur5Haj1ZTuYctl
EBo35n73bC3EGQdc7SUwyuOFZEFnN9Jy2bb0RY+WzZUN/fNnK6J2/22Raka0ufl/
iT52BLjXN/Ru36u14t+VMGes5rC+yKKK+TWl+s9hIvTS+haY04n9Pz4NXrScnP3q
nu8LBMFe77nYqur3JeySOiTxLTk97PbH1YeO4adeDfP5Aai4bOyqF9LP3MozRrGS
3HgJY1XJatN3odAQ7WUd2HG6C+/MTTMEN+eb0JT5dlrlJ+Hx0vkR+R7WVaED1zvY
IqhF1To2TnDFaiBLcOjEEUtluQjP3aXAqLYf91fgMkTvNJxlS5jNGWy+dGZt/qmT
OZpy/kppbpssDrOkU4Q6YAFygpGOGvWF28ba/4YKArxCMfRVvRQsw9SSUFVu3Qw0
n4e7yBVAyQL+9eBs6aWqW9HoLDRA2IrQe+iNxE9OxtHsOBS9Krewsdxa+UwlWtp5
ZEcI1ROQEKGXwYezTkf9Zg2wVRvC+bqNpipxFHlrR+E9Es+P2Q4CvX9eOxrPBIbF
NkSjAMfowuW3hR/xNn8uPQBCuf38jO5L0vGIsq6plx4Ippu8vFSiIyP2P7oRxILg
RmtAcWjYOmuJgDGnq7tu3D+3IqgROe+vllT0g/C1M1s0Q9CiOlpeUSSU805xaTYx
QjobctIqTXnmkGWzNaUvrH930fE5T7aJ27/Jc2BuxyeMo9pChbGuKtHHTiuJizGQ
+sNPsgar/cIzdDx7ZW9HiF3Q12TG9uSztQyxc1nrMnhQx/6BRBPLbzJlwSc5QxZx
SIu5K91r4OcFGFNhD8p8CcoY1f5sGaC5lFYbS3TcLtAhXqLmLxCzJc5eMVglyjqC
NO64peITlGdTRPCSSmfY1m36hzpQKG1Jj8ZJ3F1yt3vG71q9cs6pxsD2O9E5vA8G
PAyUbuRKhz84WSY6Oy2zrexf9n4wwqyAlx5aSbWl40zgWpGn04QhiqfyPrg/CYkS
Ft7fqZ+3/PL5YCv7FXh9ii+hkW8EJcGxX2RgiCslbxXtr861ZdVUmF6GXhthfk6q
J7AqO84+9tkQCPoANwmxLYUTvmcM2KWeQfTXfq5/q7c6o6QTbsGvpzzXy/90TZVp
maL/Y1dfHDTTADizBOp7fVKa6ApV+pZnA97h1NxHkV53oNoyjgZGR9+W7TebLdGJ
aivhTDTkXg41oVCCx6CTV1KREA60GYhMou7NmrRgNxMGbN1uNOa+QX/m3EaqkjVf
iI4TpD80c4/igfNKreXXc/7V1/wy5C8Q1PMKOQ704ZzWEjucZSl70LLSJmo0laGp
o8W22+bu3IoGIf+hKnbSy1y+pP2Pm2AH+qlIAiEe8Cr/by01/smbbPMYgBz4Akca
nFwod/3UIs9v09YOB5X2RjiAwMiGglnyR6YHM8m8tNpdyb00099jMMmNKT3EfwHr
aewHkGIKMWmZCuCM+oyfJEAANUflEk7JnE1HMH1a547Hynl3PT/TDlfRc8RvxA9a
BqZVyGQoAUngN0S9gaJN8uokup7od4SNXw/408/sOVsbud1gH4GEPEnkR279PLsu
trvl+kXVy1nPn6q+7uq6eRjHe2rjMJeQXTx3wcfvPCPpsasewbDqpXWRvUeJ2X/2
QPnxWnK1Vf904VmJwgaY6yxdq4mdUpujqGPB/RcjSWvQSZLQYNtHS/3mXT9L9f3E
O7cJ3RCfSQAlwggKEt/f8SxGGGi62YEIw5EkrSGz2plxaGdyGlc7QrtE7H82G5Ko
9lqhJb87+qhClvZRaXnN4sEQWHIrdvMh4Wd9hgoOXI/34B1e55sLX3Sac3NlNFYg
olErg79QoylasqzxryAUwb6y7tGuuM6S1Wd2HxDtzVisMh9C7SKBkEn3PUdc4Ftt
M7NwMJ5G7xZ4vylyqh7MkubgejUfPHVhDut3X09tU2lf+p08ZGmoNT0FyWbBkyFP
B+cSefsne8j1ExN1RVtddAH9SJyJGokPuvG3C8vyympqrQKUYAmptU6YRYKC8oaK
kESwDT47okjYmxa9csAT2LZ70R5RotGtmyeCgt7g9tTDLNO55re6tyhUSH0IeLkI
Hv6ijRbrCJQogXcijzoR9lCxUZ2msaDgJ60eqduT9DOXllLm5jQBIlZKhXniuOhf
rHQ4j65HYlUErpzd6uur+KIRr2ulq6iZ0C5EFSEfMr0dlSK6LQ96Yv4Oo+lu6jbE
nxO2GZNeUG8sypRXOU42p108bG/yXsWBPkn+uwq4DcAmk0+FsDJPtRM13RXogwPw
DuVjOTHafAGw2ncRs981iNShD5KYWjfSuz4MJ1cUIrNbO/wW5pqVNxQURsiMJWGw
Q2D7LzZtsX9wVEtkehCL76A+UNT6/D0W7632GLiV6+MuHRk0hm+9wTIrfSQreTWK
P3z4FauAyka1iPfScQYYRTWAQz3Jynmb5QMuFmfB5V1ndegATljtwmljCS19JM67
F7F3eDyljDb301mLPIFSNw4bMsWLJNMiPMPbALNBB133Rel55I6APRcXmXvBlvCy
0a57/WJ9KTy4Auyb5OIwR0qzBwG2QCGUNT/uL763wTuDM7bF+XH0YZDp8M+ZF46n
NGuY0I9UUDHIbiwd0KHa3juKt86Rf67mipdrOXKU/AuRlHHEiNcyfjzLuqMWdz6y
5qB4y87+wbA+eLp6O/5GxsNz6XxYM9JenXzDjKc8F9fyziSubLG6gSPWi0bpekd5
z5JG5sX0PgfoZ6y5abz+Cu6TbqoH/lic7TrypsT4JbyC5cRDLGfE18Lj4AWif7+U
oQxNf0C0GHwznQGXY8Cgqz81E2vC0B8XDLUkncbL3uV32XIL1Ebs9o6FQ1+e2dDC
CqIxC2ZEcwSlR0SWXKvacgUSpTlZHploY1oHx7OzHwndc4WITf+Fjd6zCy9XehBW
lfeIYtV8xmAWT9duA2/963L2Sq78cZALBeGXeiUFAcZd+TtRNVXrkg0V0dQBZqVP
l8vDd4dhj0M5lch5q4i+OZwN+45J7A4RluwBFT2wDzlCDfBRBM5YyCYqBelXgNVB
oQD/w80fEdgVYM7DeDLgx/Mk1K2f2qXXvsUDFcTMt/S59ndwFvW1TXjx+LsK3s3R
T6nAwHR+zC769JwYmCMdB7gt+1fe9AkxaM1pSehSpr3beTIN0BtXDE6r/BIfZAsr
ewReD2y9fGO1nntOXkxtsCa6xrDywCiIL6GM9Oyw/XieMkR3nxXeIfAcHu5wKAHx
+VjJF/V7OtTpHq1a4NedSulUbz+xOXLDEWzdmLdJq5XD50moqxRfSNEAr302RsAI
Dnr/KO/fwH1s3odm9madkFUxG/oS84Eff2Rh2ZkkajMfn0bNN9/bxKsGhoyyugj8
7l+zTzEAT6ksonVa6L2bzd/2Tw87eRnCzfN9bnKJXg+dpCn+yL6EPnR5+kgPGsIT
rwS3Mc0Uv8Gwjb4WtAxyhYOxiVVxl0yPsEkguY2UOJlFS+05hDUplXA4aHn9Wl2V
ulztQPSF1csfM1UIm413jAcRZBmUyMDU7OeyzulRqwWOYQ/XxKZ8UE88hJHry/yv
sxHTRYfF29ieLFYUc9krAKVYIghY9ct0RSs/AiF6/A1ZeAsoq/UIkDPlVcblZX/e
6noT6cwTPEGGYDRqwzw6YZqMV+g26p2YIt1ZRb6CKPjv/1QBnBu2FLuWghmtD5H3
8mVTFA2fwGBMjS0EpR9BWhH5mY1V3rGKfVxFBCfpG+4ibogEb9G0OmabxgljrkpN
OBnxmjh90X5VikIProERKtI4NSiyyd3Kl6ILWtPsggxBHGyh37QSgI5PzSRk/1y2
VuZlC42elzOwSZfyap0XSLDAYCmke1yyBsL7tMTr4eCNkUg3GTbHsdYVGnoURDGK
iQiNUCIaTUD4NubuNR/Fr4fg2Vhvrl2r640BtR82PXVwlzSokX7O5/bbpOCT79U2
MlHhr1AKeHS2ahGlggEv4CVgucN3mmPHZLxQ5ukeSKDlBdO0HJiu0E1Hc+Ua+2Sy
40sKWJ4HiQ8jfFf0G4ea7TTw9TIJrW/nJ8HTjpHSMQCbUWnLuomO2BmX5JyNIYQ8
VIDRzGIvFu6Krx7WOiUQ8KFNMIH5gazzj7X0Ot3FXzUpGCQsg4vxmCVGhhN8ecHl
U9XnVIGMefqqYB/79I8mfCuWwPFwCjFhMlAGeyXsPi9+C8JPiU72f/efjYnuSNGh
UsPG1cTz4rQA+sLajl2jm6hlUT1aSih+HD+jutgs59Pkk0tQut9EROrd1E+kEkaH
tW9UJyDGzDcmOxNXzcmd34WeA45FVgSbVJRKAnLj76V5rDh+d7/sp3nPbLWc+Miq
9oJuvzz8zv8vr6d7MKBRccNssLzZD+lcC8o7YdEM51tTgjNsbSavGyUqMsbtf47F
buUZNVXTO/wbLHInsm623cdUzuZfQ3D2gi6ArcFm6EP9xsoAJ4V8n7F74Nti4KKN
+xCfn35QMJ7bfDoCLvpWuW/Wr26WOigxtUX2LCda3uKdVHKRc3cWWHMxKj96GkWX
MiTv/ZVCmU4j4R5CjFOBxZMyBY6De5LIjTe1blZ2zJUNN94xjvclj7lfM/OlvFKy
UdIOHVRizntqHj5JpKssfdfsPT0lZyp5TS5R2rASZ44pJXhihSB0fuaFvvDrRNQz
OHvV54SIq+wHSlLuR0Y4vQVfjHZ/ygOKXTo7myT8UvrbrL208EFj2JPVppvya2cP
NM4oW1aL14sbY21J499K183RvBEbZH81GBf3JumGkwMXg2ThRwueJ6ozCvgn7S3N
uBd8K89wWJw3dFxbTallFFAnxhqEERUwbQyrpQWAcDwrwqv43d5S3CrXFRGee6NU
pPlCL72glGShzIhYnlyEfID+QJs0uhkA4GF5NUV5DRiiR+NJ30RUW40BcPl8tSK7
0SOjzhTxKlIXLfV2FPNcrY5mVRfQduICkjsA941s6ppPXF8cEAiKCe2eUzFpHn3+
WeG5AWwoUrpWOOrhPBZw58ooh46VllYYhjZX7/zgZytobj4y7rt+v3POxejbkqcr
1U5WNkcjQ1I1eHU+eUYLGO5boEK9LN5rSOttyfG2d7kv6JedpfULwNe9BNmp29NW
Ra6RegbGqORYG1zu43Sy4rLKGHe99Eu/3b0WxefVEFm27zMnOeClVWcqEjYr4uAV
oUbK7o+2lE9juelD3IBxWJfoHUNSeYWqeIOrVG4hFaXcmK3k073t7ZANcp3a6UVJ
+mTsuTVYpnM8LPAzJ72+ZVXejGh83nO+z4VF46awaoDvKkaPP+XVEO8nUsS1VwC5
wLbSdCdaaeRg8GTAEcjZIVQiCadV7OsKrVcvkZU/W8eFjpRSkDXwXXlCa/EuCgev
CP8hRR+VCrtjmDM2keBKLsxSZYMW8xiZTGLgEPjNdVEjCSmjYQ3LhlyJktGJAqmY
5kzyyxg+qrHClTsOzIgkAMDRi/25ehJdClbhE0l/9Sg13+u6dSKG0jOgqTo+NEeF
d/slBsndh6HRAknLdhovYXpPBFS0VpDNAp8AecrzfEYA72gZ96U8eNH5+nY1x/rX
8xhq3YfqRWiU8O6WEStMzRVST5StQRaWmhrF3w9ACIBtIayEtLxqMPLBjUouiuTj
EfnqAcv2SgFGyInjRpy/fe+Rcu1JbYNZbFV4Y5KhOgMYyd100gbOe8sdWFIeG3er
5iFto28NpSRAjKiPbxO9+V1UVUKHEvwG8fnqb6dKACK9b0zz+7jAioxQAE9ynObw
zcxejnpHeKVbPCiTV6bH/4SQG58eAYWNHpzz5TGRwt5xWTUJCRdUPxecJXHvd7RO
eVCnvG0mZQvxeH5zTh4vEC2ja5KQzG7AeU+Lsfeg2sVjr+15D8yq+d8jsGVIBRm2
2h9aXueEmEr62sYENqgx86QUKFeh2mNTv7Q/ftd3uHY1x25UAqmOZB3A2bbprflG
2Vv6xDDW+EqwwZb7c/OeXpRrcNa5LJeozFwDRY2DhgAYj3YvH7VIfnwTQ/hvZIwn
IT8H6xcY1skc97rJ5mnM1oFkOeW0S+Km73eTpTV5dTaeXqWm1ikFwTpvt3g/5FSe
9xB13G2ThsTHrrolSlAnEDHK+SZTUsDSAFZGiA/qDEXV/0kQM876bDaFo49O5KTq
VMBXBnVNp3jJVVanIs2tPCWjST9QarXD8pcQ/55TSiv4lMaqXgs82mFc/gZQ3WBK
8ohHVQDug8n7r/rS/jPsD/epuAeu151l+wFiI3bu+AmOS5nye2uIhrtpd5Gq8kxo
VtM3N4QHllxNg8xqNPELVLVu/Rntaay1ZQTQqauO7vSGPz84pgEOGSfkJAn6s86P
LmU1/EQvA5N15ZEFPbqvnWzy/ptZbgSRepNG1QtsCkYARMQrF1Pofos8a9Y+fube
fro116Mzzx4QLAoQ4xkrz0UeExbd+ZnChnzTX9/PlslImpeeGI+TlpJPcuHr5yWg
DnOH47w0TVtRrTDrBFrvlXJDjeoqALcWyA7fNaTXSi5q9HBBZJmXs6MkCIS+avg1
oSskMG5+EtmOjE3q3GHVFgenb+moayZeWSWh8XoAUbmCT0augW+wLNndrtLEvEsQ
W97kyYeEyVsuvVVlJ0bIn/eqTegn+hkDeyEjuDERaXRxoGUEWsKoKFiqC78T+D74
3DC/P0M7P9MN4tJO7d/lN1NpM8LZyOTIFfL7SWTgpcGyXt1gHhMJZ36ijGJoLa3v
QuaYIrVPKevGmITVqn6HMSReapRNLfq0zE6dukm1c/Jtvsg3pjI9renfC6YW9ggb
Hw6Ghp2RUBsHkJpxQDRqDPlLLw5WR0pngOHnKGfoFzLiNeJW2oLjgZtte7yXxwoI
gHKoINcWXIujLB85pxhsXfQWZMuOeMxyNAoblCFk7Y1YRMlKDpYaKlArQWhyr8lu
8Puo5eXmKepQ6qX93FDDMKDhNii8wdd6EDTXYWjknBDwXEVWIfm+YCbFupiTw7Q8
hLzdRatQiA54uwcahLG9/0wIdtxfVFD8gqH0JLN2OHU49mKaOBxAxERQzth54Zfb
pcQaMvaabt+pRXCyNy95/BgbidUOyXma6xDWsBidiMzJG4Zvv/iGMZEo5Z9gRLLu
K13WZVla/P8KpAFrCwqBmKyx65e+l8/LhOUEMMnsYvY2/2lLLf/ZYkHcGLQTls0V
FPXxYtGHTEVIEzgRI0tby9gifIzYQeZt6OKff7Su8n3Q9NOXx6hphPYmmPWpvMCu
60/KEpaKjjSEh3DiQB4sO12yDegd0w6UzwpmfXFj5zasayOHr9O4Dx+S3uKPe6Oo
9uj60ZLUjhj0ln0B+zdUbSsYERPM/GJ6zjLp08qj3ChpkuDcuDcrbN+M0zjP/27k
58T7j8xQHXHe3uPl6XBJap7XH/yyr2o4RVvJoqskdg5NufmZfwPQi4bd4ncsQveR
qHHmJh+Ffcz+fC9bOH5F8YEwqdQ/xkTqJk1Df7dHzlA9dM62CZbQikTycmqj7vkz
ee/pS6RYuCGlgoxa2r+jPVepiUMSyixGT5wrtCZYiQcP35Y0fA+nL6aDpK4JhijV
4dCAG0oX1cDFTzUL5rFq18gp9NF7WMxGVnTgEFL+ZkkwON1aXFMItRp2gK7304QF
wYFl+dLgh3bGXl4oChG8jX4AKl8vknsTDjw7V+JDNxeGWbeXgB2SBgYVje0Kct16
LG1FfoVw2/6QmNductCGN9KX+5yE4XIQY1XVym0iR1qmRcr1acwSH9SCP4IexKLa
ac44/EpuBbVUisF+AR8Rl4tkakphE5zqub1XfS4lDqSDc1uGB4NrrYN/Ebp/isDh
J98PRSxIb6UW5nObqR7QAO0Q7YvzlRZiWul7tECx4FQBHsjGUn1rW+s452qvKrID
ZiaGdREY9GMGK+ZRafvHmzrSPfVVsixl4ZXqI8w4CosXhgcYz8UKe/Qcrn/lvZ3K
lSvoOY3Z4y5iATNOPx8hE8lc1NZmg0FRG2kNQa7w+fTJvSehok7nvERfYs0jD30F
djmfGF/86x4rik1E6qq6midOodvRkqb8vXgKk0LgNgE21IPaX+BQqb4SKLROf2+Q
CHVS2rXCilz8JwcOVTipu6S+OkKDD1V/c5y3UvvYaAFK7vkUrrclRNkkx38+4CZB
X95dfd4SmEPN04QCMarZpQflf6/v6o6JkskJsGPo5ebg2O4Oq/4bfjPLmfEZZLgN
xS22piTdmD99i2GXgFgDrSTAXNGitfCAhnYvewbO3psj3H04dVJl2eyTqYwnmg6h
cdVy51neHAYSgptTWh1DdDb/DXnUPxPAo/HvAr7w0erdKSHZbc8dY0pixQh+PArD
MQ7KiURLzlX1sLqW5AzpSuO+4iCFtr75tWWjbvUDguXSZqYXIekzLzy95fzXvfjv
I1fhG+aiks2wJImrHB36Qu655hnyIRKi879LTp2xzER+V3kXoI77DpBE9m+reDIU
JXzMVdLblqkMG8aZD+VUjkUwRzasoIv0BWwF6R8OAZnur/g+vviybVNOpo/n/vl9
E4OGFDOJUTh/eZoWlxcG5ZS8iGSjnei/xiwI0yvmaaQweT3J0tDFL3Mn7P1RgEvA
gQ07W/2PufeGub07Q0Oe0Wq4R7vAU9nt8DgJolS3A27F35GpIlpNU0kIYs3qxyG3
mU7lU/n3XMEkmRSqD6yXSUCC4oNMtUOmETo8ANWgWRh+v6cQgpE0QyYeMNXqNaWE
r7npSsgiMeCcmjx9bOaLungnu2dqQZsnu73riPcvOlowWAzb1oE9A1tJtJTYlPjf
vAN0iqTq29NuAdFg7Efa7beqGhf5oFhHKJdIOx7tUso8KVj1uFQ7h5peYqEHFKhp
78bQo0htis8CexijFDmxrGIZD1nEnbNbusZXYH7cI/XFfp68r8U+Nw47ka27G/3+
m9RTLB8WX+pEpgjsS9nhL5cTIntuOLafQ3VHgy1jUPxEvVJ1tHsAAxNYketa6TOI
I/G7lQKa3TjyR/r2qXPC8wPw9RKy1pJKNdXq8wKFQbb9xT6UeBETYySOv9SOQfa6
tEbiE50W7qBdSvEpO+bLyRXjln1WIyQowRYzkMRHDRWldv8z7vz5q98npUwa4BuT
GZAAvG7aSOI5S4ftk96OAYTpOfZPQEPzPsHVe8k+hA5mSfNCCehhoE/anlAzJfn3
y9F1/+cIILPPQ9/fYnnUX55hTdlzbmZmDPRtyaxAG9UPFnn//gQO/+ljtR458cRd
hR2F7Ys17BuG7JHYGuPAYnqbSMxh/+MW2K5RusXQ2j2pVwWCoAxD4DYWx6o/mSCG
HG9J4b4PkDSShOFC2FAvs3TaOXDnUMyvCyEsqYRlVNjN+DIWEjxwZsLLDQkohtMy
ExOM0Aw7I/v4SHw3PAJpx/Fqm602DuVYIDuBky9l12qkD85/RGVkKccIeiZxMGw1
IFUt/cFwkms2CuUpISI2I3TTZZI6wS6fgtyHid3GVhFM3LjHkADrHqz2dj8abtBE
r0KyJeF++FnJJTQnXQMEfcogToGXslHUnFiVMbcbo/rtsuChVGDrKVL4n7Wfk7Fk
GAe0gwsKX4yIrQe56DiTv7/7yq33xvhOX6id6gdo3xaGs/6wM3bYBApOOgSU/TY+
+BFW3hWGI5UBSJAt0BmuC2fGy3HzB5Mvvi5Am3g+bDVee/aeOa1/iYK8utJ3BKn7
jhm5yjabA//0a/oryniLp7k29WQeWjAy75UNVNXkH4OVM0Wq0nACtK6o9xy25P2n
mc2zKavrGODs5GHbYgcl7D3CRpaj5O8vCIK15aS5nTGmkr4/6yCM69cnUfSoS8/K
Yc8mskbkUaQWDRrBVSlluGyzOGWNx45v8kfCM1h73PDd/a4wvYcukPQdnpHGrocS
IziICJPh4KcdUNVlnf6vz0ke5JJJWmaCguRy+3rkD3hYl9q3ecsdpkmiXpw2gdY2
fPX4TUtQDPLjqNohUgV5xXiOYj8gfMP/0yfGK09v5mtB2gw2ClhLm+BETADW5XZV
tnaYdfujaMpF4OFFrN9I2M2Kb/cruGXgDado75mgB1ct1JJMopghyd8P+REUQN55
MRzQTuVkvQxgx8FSfTnJXZaT1N1lTur9oBl5XqCFiFSyFIAFPwRyOd5xrB8YJRTu
wSs45ptB+4XkhiEYQvqThtXPGmEviM7lCFkAaUBhiVf0jP7CVurPao5Mrwg8rq/8
5/14ut+PRzezRhnE4OJWQZ9touwGztyXfMCiumwEMYpWb1Jl9DZNHxqpm9nCbKNV
IkeQnkc21c4PNtqlCRQ2O9MWnNsCw/zAUOdCHttEJcP730Yjav+zgnx18AePbOxY
A8zS/xMNRlPWqvku0MmqiAT8Gxf3mMt8euQ74Wah/YoIMvRMB7C67xlavRg/pdGH
eJyeUVmcDeS+G0pX5YQPRxcWeIWdc5WH4iqD97ULEK2klSFqvYsZ1sZlayJRNW0i
aNCmHLdedw1l7JuyCanBKtPbzt6BG2832Vw8f4ankeOc7aljdOczTclrOjJPVJxc
VnL1loX57PIFoa/7qPkv2dXTDoYrq2S/Og4leiOHZUfYhtKQaRQ5w9anJ68/KDtu
AtA5ap5jQNyXz+4RXo3daNRytnpptyD8vNKOxeBZdc55kcvdu8O2Iy5Y3Hfmp2pV
zHYbkPJBAEUhtHpWw18cw8tuAFXy+oUIK/4GrAzZaMXPGrnjveAJrdv8D7x4zmdj
JPEg9T+QtxIu1tOx4ju+Qh5hCRz+xuIuUOmjoGeLhNATEXkVNhJwJjwRZ5uyk4cZ
ptDnnYn+EjtkTnpXnSzsImep6Uf6YRD0pEcUM0VaEeFmbtA/+bBHz9eu6wQ5kD7d
GosXJubGRUzDNLcAD0tiQuxfHTNxjmgEQ/yW2hOrxqR30HXYm9kbUAQouvi4jdUA
aGy7IhVxfTDykYwqK98Zn0XGPTKDplwRPnEuBLN426reJG0FrLpU+DynIUsosS5/
yXl+ezFxMr7j86DmgazB/1Ki310vLuh5eOJp98OMyi7LG7qR0hIsHIds9siTpL4C
PqLaJ43+ir/kATOLBLyH+7laGs4dsna/Vg2O1aftCRUeGXcehGojNDkCkQwzV+hf
zmwt6eHlkKsSj/MS0wjMnj7nu/Sepul1qIb07fvtGBQHw47W7HN3XwJfBEaJl7qe
OWPacBlqr0uqrqOTyNGMmYvuxSeZld8BlY+S8odGzc0s8N5dPQDpAu9GOwrMLA/6
49YSYetGBsFeZ2eu2Bife1mKj6Ubtfc3LziReK1bxR1fTBzhn6gDu93/weCwmX7o
2EXpmafsPbZtgaoygib0Yug8vKHbO2oNK+jW0rthXbIG9hiYST1YVI6ejB3zjAly
jXOCwwMI5z8AOCK/ela9XkXCThdWKNHLl+eu9H3QYjrgHPMR6TuT/lWMJ4zyMO+C
CmiPREa84+ygO/diXlvEeurSVnLDgshRQBfeGrqGYB5m+pQeylmJnPFWENZg7fwL
d2Hfd14+AvnXm/sFR+fO2j6vc/hwHTjsFHpsylGbcXnwGlcmiPj4T0TLRTlDLttm
9lrBefmFQ9FJxN2ZifSmKqQ/Y6NQTJzhbuYOVcs6//doZioNZ9DecII3x7vkX2aO
oXr2kdUCRgW1l2vzeNnJcIU2TWk/G9bfL6uR23KPxEpv9w08DI1L55vMn7ex52YZ
szsVF3C8CPTaZrUgBNXVNjfLD30sdN/mYmI1ueN8hrqt9jtFOl07+aNHfIf2pkZq
DorPAbOfeTosWMAV9tCwQKjOIe6OrqXaZw5SOLfE06g2QelRD1Oj1IuOc7xE87JG
GFOBqxoR5sknAceACfBJrypHAfRjtSvb5rQr5XVbwpxqnVHTvIoYui0gxXHdzVX0
0jsuhuKhr8SYTKU0z/QoC0NAGPTXK8amJAFncdYHnHGp/vhwlORNz+ziQdJao+UJ
a6QLC5dIBH2PyP/zMPCtKVwkVMwiScwuecU/O7fVOZExBNq+M7khUP30XIMNsUPB
5rLK3bSV6QOByIQVWxn2/aYcycQNPl3CWhyggObl17582ZNzHbes6qEbE+/M8STB
BnZy6ioRhHXgleeetlxHTkGMvvzCJ1gpZQ9zan/PH4+eeva7tZh5kQrjirJpms02
ByqeQQon8wkucIDik8qBayK2YPv6LunSLU9AcCVwXOtl6Nkm28b3GVuLjuFPHTw+
U0Di9yZOrODxAKYUv+Vsl7Tw9SZes44gRhW+biARh/dEP0hRuF4Fp4yi8izV0SRn
bZuGJDYlbfDkS4vXSoYdLfjOPSj+hAM7G7ZsqhhtMTNGBGq6erauDCIqAV7GZOa3
f/1sdG2Jq4CPf0HYFLk3U0XhBgfMOVRsZsA0Fxlo6ZpA+xL44X0K8rDCUiNXujn8
CIVJEYyZyVNz47dtErZNgoj86U9yXNmqIL7AmiWqBCzpGMADf6aZRNhWB0ww1Dcj
5EQfUCOYJtqm5+rGoceAVQTxXT0HKKsDWqihyUupb3rXMBRnC45OGLL4fjXjFOzK
yYScrTYUcITMluBMg6+aFcU3xHa9ARrLYiAWl9AnWwcx5TfR0owMpA5V5KH4JrEd
fkhK6HVF1kdOoLFCtXmHE13CwABZFgbzLvF82xsg+uE9M5agWkBpton9r/IYDZO1
pw0QSJO1WgcfO3zgpPf3bh1zrFM0gkaFtOPsmX6TxvN3lic7/w/xvz5F3GeUvZ61
9MlP9JffNQ4CNGgAarmBsCxbtrJM7h4hmyYc8LbEejMI6gcmVi2a4SKx/c42KcMn
fU7HXPOSacqC8syxOJlFrxX7NVLy8nMv5Hb7ikwIamxGLJOxPdqCtmywOhu2vscL
LhqwGH85z+OmgUeckaPGLUR65/4r0KMgYpVck51mYt/0WIOQ5rGYFsQlqE4cPDKX
n3M07ZbC8nYcF2YQHaWtxhmDK+6UIIMgKQe1SBqk/3XP6utliB5LGxG0ANMXuo99
2dYXkagBKO2fRqxZmhW0io11v5a/nt6ZR5JLSVseE5yv24KGcepkTdmL8LVv25nb
MQZFqWVf1LF8DmZD2NuHu+7h2pGnstp/yXnXXd2XFw1utGz60qE8yukBISQrjuIX
EkcBFJ7x1NLh7rWhV23K+7sySFDv/AhDFQ78jjD/e0IjM5Ya/jjuTYtcY8HAbRib
KFhF46yHRBK+m4CVEKCmD5cZPpY04iDGhVJ8Ab8XumsVor0YqhdX6BNjl2rGW8+T
qc5wgOZGyMWbquj1BfJKiiS+o/Zd1wU0shBjH74sQj66Lm/nwdIlQkFv94rxS8Fp
0P1/cP0P+V81iC0oJFqzkm6uVYNt6fGiulPkBbKeeS43iyOb8mv6A5YqjFMoLaes
MgMABmGHD+iJx3QjHqMuLw0x9OgSOQ6bxvri3oToj463Tj9VJ78o3+oCQ1vXRaO6
1Smeugvy3+01Q7lK+bBCNFulz/CG0QnUQ9VYKGy1rpiE6ttWGz6mVppXaP36BcZM
kTztrdKWEU2WFQk2ipZ8/X4AbRbZAnqQR/599snCDero1l9WKqU1bX9dNzh73MUI
I9x88KX7oMTbu0oFaf/EhOcH6RcRuXoDqG8cdgO66Hw/mBXwjvsZLQ4C6uINeWJB
ceAn4uOPu1GXOHdrLpdFsgboWpQVr/cdWD3gMpcj4BNOXkBnyiv0prjkA1Zsle67
GDMGFMF8WwM3NCNe/MqvwUMYBgIFfYgx0TbY0eALG9jXCAql7rN/2aVJ1Y12/wUz
/rGDt9WOvU8PLLLKHy1tinpqIe/NcvHhVeGgQBHdvusydU+7X9HfZ8GdexDC9UFp
saCwe58j+jyTg/SueokLkjDRz63uiTkU7UKNINPy/tRiEzH37tDJ5vN9obNjMWNh
/+m+Fm6Ej0ydaM0v42Ta22S1IyiK5kG8GJ27oQhXCx3BIIkXVTBGfCFo1CRycrnC
LvtPHHVivvivKRRdCMF9kAH3NEdPyH42w9w976Qsl1RXP5mRGO3ECQRE/pXSvvFI
0c7scjB85B4uYiAYokcsFRQuwytV5/aP2Onc2pZumERNezPrC4jVcriyK/vHHmXm
Ln4ndkQwjVkSUJq1ZgjeNjCDgbclyde2aOrHRumT8y/HWzwPWwBJ1uGzo3RXhOMy
5iwxNbaWGSZpubk5D41A29Rc3NzUB02RwuXA9A4Wm9K3rK54A3Es/oOl/ic6Yzzr
/FxjJ+ZNyCnYmDQQBSG9a28DOvhUbNizyh0fDw1qYx/fzT+AkJbRIprkTcZUjOqN
ncZLTCovDfy4k8UAdQEYZ43eHprzWk6otI1NSW17TeCxcIm07uLBaBPXaGAQP4Kz
FhxawuQfbRkcQqoQVPHAVpONuqoBoFE35KFBb3KjpmuvwPO5q908LEGssMqgrjfK
CV4J7kFagHJymdeeG7ojLGOhO1XFlA0x4N2k/Oav63zoHrZnqDGvmrx10r4tXm7z
bNFenAAa3mKzEdZn5TRUCe8GyTtmb0UsYL9++g/zbWo1+7tVl1yXb24Oh1S2g0fZ
djlaCvqxOAGSx8aN3h4nLEBjKEkG3ptCif+8uqpa/M1s/EOvmB1KJa7n7zT/HToq
XEF+z1hko4oE5Zm9uB3heqBUvJvamE4WrfeLiVV+DpvhGQ2V7Lq73w4GL8ZQW3ie
8Sw9zQSa+27LV+iVKhcytTy55PuZbqQf3YCtHEdj0a7+oIaszr5UcuzcZNFxCLCF
/gRWWUrtjkH2IQQ71RC73okncDik/HOjmnGpUQiefsxBlCNSAvdFqVMZUVDjBf6Z
sjDKyIIBRNkCXubShTh8ymOF0iK5UTZeXT82sux2ZJEaEsSwM7HtNyThvHW9fspf
S6gjeLzcZl5FI6+Kne+auJk7b6fuRpVbzvpIxad5y4neoK3y/2/sRmQiQFRV8nhe
GCCO42hGMZn1cb4Ss9SbPfenYGBGqV6PYc/mfQjWRWUWbAgMmoyvjnfQD7MW7lOl
OXI3Lbm48Qgo59kINyGICQHp03XRW/zm8dUtOC2VOjkS5xSIfgpapvQ2XgXC+hgG
q6YIQ7+0L/67Q65TraBDOgXBYnXwhzcTr08+hkuN7b2ggLGPyr5pqW/mEMuEHwNG
e4qLhJ7IGSJNxkWizEr78dFw3oms7D8Bz64P9NICMjgGF9XYvWUCwWSxvb60Swby
D5ggHMYx/EMHOYMGsyCR2q8qKEpsB0O9okauREjmcP5KKQMbP36oCr3dxF7Sc4jE
f0zEzEOohyYAnBkCbvrhhUiRjcr/l/z0qDQGt8U3wd4ESJVEQRa0yLwm8GdiT/AF
ZQFPDwzgqDJgEYCLO6WaaN7srZV2wMsUIGawlfYKmovj5Zw+EmfsAz214JrHhH/1
WtJa9AtWHB7A9CRZ8JX8qDrWyNce2UTgR6IPUyG35WUJiG95IAYYETAxBhZfSUid
iW3F3UIer+80ljLUSUPfi2ErQ9OlGxkt5XziX6Q/y+QlaTff5x1h3CdyTGsUDOlh
iJYAoOT5YO/9Xufn75S+80/HQKWidLZELGEnmDeSCkSyfNQEaEVIkG0Seg3jnqZJ
nCYu7hL62TW7PFpMCVpI++DtkL7p0R3+/cejsgYGdhx3zuIUHzxHtACBEGD5egBZ
NWuAqi9ipbXDbNVD3h6ZZ7KS+FaIW4YVVcroafHnlXGJQNiDcPXDFCDU663kcxPZ
pqKkUuIRyQL4hlmKWCpNO61B+qOh/iIQ6XNYh3goLv9l4P/xmvQTIDQXCBCbAebL
vxvC/aloSJoXzgMoiRO4eTORfHCIRrPC6f9tZa1CjGTSZZwM5Elsb/Lgj01C/Foy
TEsJ+87A1kfvqQZphCqjmER/4iZDxKGA9C8cNCNSLAVVsbo3Aoq7wxL1H+J1SNq3
Gg9vvf3dAyY16nOnSP94bEN8w/I6nubhy/11mal9+kp9zbPE1/6h1P7w8OfSs+bj
4Pqxs/e696i/1dKo+mK4Iq5bf7+C5QC0UYSjJIbWiOrjCixZ/aORbCAz7u2YcAlu
Icb4fLTrLccmBH74Snd6e96Bd7/NvY0rGhZFOrOQVcBkk5p24gtUtz5STMl6M+5s
miLsmEw3d5ycwOOo/dSywJQ0DnId+52gw7fz1a/6Zy3yfRX96qzdUxqknZP/3SH/
POwQmvPKn/GT1tmPBA2ruSOel1Q76W0CeMaVrITe0JxJiaXVA4RX43DOWjavMNTS
8fHQrPFkwk/JpYEOpsbF7GLwD9HJH15W+hAROh/VDR9TAB/WUmbErWuMVuRuD4P0
Dvrc4A9U33bDlFsI4KTnkENLGsnfbG4L5d1PhVuSkyu8DSGEDUPo0gSw2M65a0aX
L3xsTHg4BoKad83WUbS0Ga3a04TCXRsQ4ukTbMnh46M2GrSZLS8CtlKP0z6itUNX
i/ztlFT57UZs+eKpMWTe/nNZT6LW2WVoiQNLhpVbFOiocwdcd2ezJy3qWn0oIhCm
iru+hVQpmIniwqgSTrvCFPxAb/YmmkAqoe+fY7IFIvcy8O5jmDRKa4S9jc/V6/ul
znHN+OILVITCl7qnUQGPbo9uB3b5ga0f0qx5MTQB4hgN5/adM+Ep0p8XGnyLlZtl
+2KT2KvORvA67KbXjMYc9mNwMI5rzFcAqIkU3d4E2cd+JynrtEFrzWB4Q9mkOd38
s2dE3Z5bu2cVeC+dAgreq+bMKElLzN8Vr+SaRjNdyTyB6MhqpNAJN0MCkI3FK8Qn
yPYu9+lBSQzWEuhU05gIfawB0xX6Ml2c6lRlOptcUYkeYjYjZfN6M/6auvgg9r8X
6QQfiOu6eSZBzkWFXUXDBQ8kCh6sig+1tdVThDZIToOWJcFEHJxkZgsAb8y/ybSz
c7RcmOHPaMqGllVbGCE00KxmEPmyd8qz+EVIyXLqvq2KWEjPbPtx7zlINzs61XAC
ndIklWOrX/GzETG5Tut5jQvHhnwOYM+EugK3TaCz9VNcM3IGMfdqGysJHTZajXt/
Guc2WVHIQ+SexhhEJVUWCXipu0trfhDpkZLV7xPej0u6uWkH3kcy2xuu0vghMxTc
SkGVWv4TSGOHJtzS7aln/HNDA4XnTh6WgkQNhNFSgARkR9FOARXvc7/3Wkm8+Kvl
AfJ0Wz46f4g8gwpcDN6NCFzxDFYYqB9wPnl+7y+2uLiF4eL+2h0v3KsmEZY40/Dd
Fq5+mDr5Fn6fEKbHbgY+PFATRuMhoq6qCLoV3O6gYghHMMI2Bpi087tV9iR0QSnY
BXRgZ/wdVw8Ay5Ter8bUpJeb74ASlGZWA6/pAdAZhF6fCLqtDXRnxek28iJraaPs
VF55eMm9wdlPgSlKlphIViHoKF2DgWalalTm9fBtaNiAp7mXgy2aKvDwl4TSIzZM
wKs+cCVKO/4/M4heWI9/cbXnG42Os9qfKi0KrZwLgmybEq9SY9R3JRmwhs2BWKYQ
yUP5DRePBLU3rpPhYAqYL7kPz4V0dVY+wSHHdrOaCCzRUaDLVMHHDJn44R+oGe3w
dD4NLNCqfvfPnkxjqe8S7w0c7K0/NujJAF0QxA18LepMRuTEztFSrPbPE7+cz04r
uSyKIKEDBvrplxdIjwhrpyWED+gKthbrST2xU5M8eJ7vEHNHXijarjM+OC4kFSxV
BDsk/rlcz5WFv+qDFxOxF88ZmV5s5Xph7a9LDSfcqPZ6KE2YFk1G4kuATYkxADRj
yJ/J3wSY/sw0tWKkeiOl2jl0vHZu1tKpOnbhyMVz/SG+uyJwCeYh7eHv2mKa8i3j
+vWVu4YcVv5dkcIZmF2iNWP7UsDO9NUjEwR5pB5kETUO4iHAhcbwunTjcmf9OZhh
tK89p18WE4o49mG/96ZetqmMwZl6o/jTK+QwLFDKUWAHeXQv1PnxIA7EKvC7LHPy
CZRUr/UqJbzvgoBLBirQwl/y1CpOOjVr4Y01ynZn7U0uy4HPbNaxndZnpZsduDVE
PWwrUlMFl+Jes44Urd+y6k8C90GusAyQRuGmR8pCc+dTO+YrS3jJkT+xY2nnbbss
VYuCCFtcpqFUHGCjo664HuRqP2G9D6utPGPAc2ojPXbcvUX0OzmcT+0ht6vsKS6j
YsOpUweXhVN2DqQy89c6GG1/b5lfu9OAXwEuMMuGoUxMRQ+n8hX6o1f2ujBM8wIK
Hj4mndzJ8LSPNkpaORcDd+PIlxIR3a/F8mj5Wjk7HweJD3RAuz2jDrVmmh6uKQdY
pqLxO7tKMuaR0Qc/m6qSto17WZLXxx30lWlpuikJ+W8saAB1wXi7afeu1ar+egGJ
DhEq7d2cLL5HHkF9bJVy3e4qLwHtgUW/1w67jKWCePdhsQ/gsMBBFif4qTtWuYk4
I11DfDp4fFpujIziBQoFmVoSt6yb9Be3pvqqgesFWgisdgEXuu7OjjQpYWkcFtiy
kdQhoi9aD4JfeXJcuzQ2hZLHLdMVeBncqFfMIoASRzWh3S2ck0h42pJPzXQI3BAn
A9iaPyvbYRqxh+5Pk9E40BvKpocwy8pXyrxKBv/oa2E/kljJrKP9USVBVrw4Egvi
2L/y3A8BEoDRiueZzQ/yHLY3gnfvCJgGcLl0gl8cVEmrj0EIgcb0JLJCjwI6nb+O
JzVPmU7SRefTB8TlMnwznKIXdlnH1X/EsUULp5Jda851Xk+WVrf8rlUAPX6ZucpM
94arm2hDosen43UWGeKkd3PayrwCekIGOvZYGhvPCp5nLTXRFUo4b+ueOJovh2qd
sRoA0pMjRZggFcjLe9cJbQkwBOSi/7CKGT+5xpdRUySDjmyvuG2g6A4tMfQNbwWS
DqUQ8fE6VjmFEGKjNNGgsl16IVP+uTZMoc6ItUFJeaj2Im9RUGhvXVvaULfEV7MF
pNYMeQ8DByeWR8iMBy1fxrwtVRLixfma7kvzGttRFiHInJXWBVIm+ctFXmCGdL4y
uh2EsSsghyuY1YWBv7pFMfCFCiwWMOOvTRAbfLgztK+v3SI035eEqND+nCzYjr3g
QH7ed4tHYhVgWZVv2RIN2fmIDW7voD8fBiWbOQZVgiDsFBp+ioh+5nHzRqDOTL07
hKyepSVHH22QnKLn0GgYBDVvOi/sgQP7S/DkuvVbjTzn5WQtKNbF9qGI5K54Clj8
es+sY2aBlp4gUg/HGkVRv25X0EbajwU/S1qYUFwAxaZRzWO/IqcbeInE2E5NOXhq
/29r+85JsRAEXUMwVrUFOIU1JAah3AiUDrqjso9HkYUYp49JSE3AQJuYEnIq0E8B
svINdB3cqGv0vWhE1z0gDIWjMm34VKZSvfh58USracwWoNKRw7uZx6xrgfFElbZH
rnGrAGhTEJnSw8okErvqtjUCpjwc30VgBzO/i0yIJ8CpJVId6dUNScz0+AxCuB6Z
srBlqgTiWkgc1MmknKnk5o7qkP4R4Bd7vjETr12UK3yIiq5/u3dUJ96bBk+knu1m
hjyMzIgXy71mvR6wAfpUpBsK5Si6V4uYTrjg6emIYRTo4Q2W9NmpvIg9OgtFcWzS
tMNwTmzRRil/qoTV/qP65G4CzTAiCeYV8Ph9caQM354c6YAI7p1o+RSv84JnCHw7
9bYEWz6z8hGgF8weybwW5ik4tRE2oiDuJlY0xLrEcbkZ1LKqRwo1rpjDLou6uwIT
MojsKMtYYhrzEPXCQvlCev6FQkpTc0fbxugGDqR05J9K7A61ZtX/W6RIquCMSS8Y
kfrD7/P6V1dWyKbltsomMMed7GMIBsjzBoTF3CrDave5Jm6XWoIOmj6WbP9SdZ1V
cJvL2lKhoK6ZjEjAz4OBK/QdnD824JUPNQiiW+m9tf+8d1hjdDGQGqgKdlg2tdAd
VuqWrzvIXvbrgJGk5RN0jpOqONtxm1yMHVQgXaky4A+uq7q5HoSz4ONXDLi3XGLz
WkD5eJreITZ50EV7CSHlwR6O81vP9R14EE5PVQD9KUK6aPJzqhAQEr/wMexid0yt
A5NrBeVy/zbnmXfDKsnCRgM1EUPK8q4fWelCK5F8TPNaa6/CcitnPoRcolpsr0mx
vlKw7hEWTqBoV44cU4N087RKKOkPZJ87nL6LaFFa4Sysu5C5YXjCMc0B3PYBp5OF
zoOMikLRc5ZzVP3TiF9T6QIvsBOlmrLVQHgjGTqCFO13q2fRCKjLcbZkXfPBSdBu
T6QQe7Ek384+ybrAXeCF1tAYiEKUI8DQ3c3yHw44x7WyeJlB1Ev/EsYjKg7vPJSQ
cu2sebya1uUN1SKTvWJnPWtV8h87krhYeB0c9mSf7rYuXRiVOITsMdjW3PoaFVkb
m6293oXTAds4WzX0JTDlFTw4AqJz6bi5FOWwZ6zqR1XTOOf/OILjxxrSlLEDVqmh
WKxb4ddSPWLv10wZw9adiJ2ciNIK5rdyIOXGGxLOMJ2zOnRfGkkWEL4johzEvUXU
c8wMI18M8TMJ73sUOMWnqNYHdvDMA0AkOThzbl+zVFYgSh8+otbtOH8SFa5VgtER
QDOkEETc/WfjqfvtQro1yWkgNHkvnYgDI4FtX3W6Hrln5S/KOE9GZIQ519Doglh7
69n57twVSgkYyeFjDmZ3+8gn7FjWDbEjRcxXYIyXYhrsccqMmXMrGZK1aVHQGxSB
+R0Eh4ESer1K/IRibwKjeUpu4CCeuZBsbj2cM3YYhMCy+Z/OEO+AYH9+F5j58esk
yBRjTPG+CbjmDaTlHFecFM9WYYpsYTFEdfYgJxEX0TT1nnLFfsgOhlPpgXwXxp+1
P3qMBLiV/jww7cy6AKGFgyuq4VU021p3jR8Lk/kpi0gnNHGIDwEFmIIBKrozMGKV
oBYgMZeq08YGvCT1Aq5bdO2X+BERS0/uNasbdG7dEIgzg6tU6zXzU61b82CYn9X4
veM4+jSl8CpoexeOJPrxq6jt9FFbEpQ0IbMpXgHZ8NukTFGABPZWi80e0PqXcyPt
t09D8a03eED3JuI562KZ3wUymJRPL38+ooR8HkLEYdfqYyPRBZkYUXyqSX0Gr1yq
luuKqM6J2Qx+ajXAVrYbxsTitSIMokgiSHBPfy3PmtLKkzLQ3MtpuJiu8cKivF+s
MU3UG1eaXM0RURmwdD7uF2vPU2OcQsSh6OL4ZZl7F6KDSsXapXQUvL71T2duDVJq
YsrEr9EPeSjbg/8e1T1FQtjIoy+j9H77gUKLvTYAhZ37X4iddggxrCrNf/cNcRwW
hT1oUrsCyRb4DzQtf8QcwplJ8G+5RUyazSaMVzdtFK6LgrESYj2x6siE7Ao2RFv1
NuYh8r6S7douTp+yc1/2cgV4rYR4I2T0IEhTalYXhOKlVMj0mCuEoKnT/kVPMjRd
MwcE64e5QfS2xCqyAZyLHo9naKMxU1cwmeKF/vPb1aTsskaEDiMUGhcm1kkpM8Zm
OTOnKwfgK3mR+NA8bHjlL+5xVn8k4CWo3XsuoT+KuQrO1p78Cd7/XZtRo6pE9u5n
ANspekI9T6SiPh078QARzvzUBziljO7WDkpVlSMXb4TQrp6wKW8COX78/j59NXcn
8OnikR6s99qqvhwzROUuNxbAafzSMF6YrMu3aAMlzeCp8Rsfx5BLB2E62YCD7iXG
8KlExQMXeMuu/TvfSPrVUHAKeCY8pgTsi6l4cUYJ/h1YyJZOfO3AedwMeasv5LIm
j4IE5Y92dOCMp8YBRyK5xHcsyjF1w1ZPNh7+FoeyZjLPXDOM5R4EqM0IImEWSKtI
kzR6EDmW5m7wQ9MHr3Lxm5/lZY5v78yy1yBfG52e4wlGN+Dz3E75Up68nxO1Eycx
wySRFsgRU+yXXzFGPKcLQnKM8Px5jLaIT1WekOAcZK4R+8E3cbGVN7iM9C4ynFNq
AvW2xULJvvW0pOu3MVb30lc8+b+kdUxaPvnvreOvzD/h/aIN3E1Ldh1amI6PquhK
IZ+bFv1vtfPXTEW6LJTGcICqnXMo5Oni2dQ7XKdpb8qN4bDne+0m0ZJasdAHVkYD
R2f2XWBq0RrdYp6TNW+gmldG8I7ePPrx/ZMYeWmpr57Z7qICof6/Zq2FOSrBcQwW
RafLVsJROg8qB0NBYReBTLqnD/7ekrv+D5IG2AYNXn67Y5BZO2cKlzCUHb0br+GH
lhW0ME9+YxiXN/K8GYcaEwDlaOfGeGZ3uiOrb3NmOQYe3XQDXxjtNK8pJPVAcxjF
1C5t955X9mhNrVQJj+EolSEqkpJGF1wJCoBAS57Ax+5jpCKo9pSpIJ6CRnQw7cq1
NZkWMJ9rL8Jy/zkuCnPtMnHQs0EHmwxDIwb3rVqOVngP0UrHoLcBK0rI7oDOOYiN
DvU1Wq0WTR9ArZciQNEXS8AZE5nFfd0yz/IwzIt3WMvMjEPY1zUpfAQQaGJtC7Ff
K/niCJgEHp9Z1Ca5t9eeOTiNaNN51Akc8QBL2+BGQkWPjmFk5wuNVDCcMFCZUp9b
G19BLUe6hXDKRXXx1ZnDg2bLXZLMcVL3chQEAKrnPw1dC03SrhX/Zi7w5ITuWsR1
0wLVj3UoGbrEb4JvGqyIAhoIpEGa/qSzrl9DNMO/GOePSfjHER7xMOgYgzfR+GGG
tj7p8Du/FB22/ZmgWwMlf3G0F9QyBfSE0XqTPI3pZrb8bMkWNhjuG7I6bzctlfyU
RX7iQXP87e35pkI9vW52Xii2AcVONpgMZUzPEvfjvYLSHoUQj2pXuwVEUn8MsauX
YwpsQ9cHtnk1/ulx9eScMPgjD4AXIAuMu5+ZRLWSQGG8nFvq5RGmVN2+3R8++qal
BTFZ8fuwF2wtXPfjN7m4cx9A8nIP3fN0l9TTKTFzKw1WKxPmp/Yol1qZJFefz9Kg
MLIrQ1jeeHl+FljNvXVh+B+qiX1iiZ7NLyggo603GWIMKOs6zXEAvClycwlNlafD
ragH34NtJoZ3Q/6oZR9kku+pw3ukXcdtf96IxDrb59Q/XuToFM7adAVRU4ZatrEb
eFp0cVRIuGHKN6Mu9jdEsniw1DxUPHtoZ3LGj+LeaefpT/3Kqt1Boj/WK1RsG32n
qwpA0ZJ5oc9xK+luM5Kwj5B36YNdrEBzdKNDisTp8QSIh7bGpSFlduP1qGGTT0oL
N9PwgZVKhGyYMAbCfqxiuYdGiIByufg2c0thvZ6ePv+jky2qffPZvOFqU/gSZFTS
Vagv8v73DEO0X7iR3nn53bUkDUpkYk76gT6YE+rN/F/QjtoKOjadi+PjMQLgt5XE
hSWIZ0INm+7HwpJFvi5ftP/N57Y406eS07qL7WpD/lAsJ5Ea+reOfcR/Gc/ZVCFx
mCvkF2ndlkQhSgTNvtJGGLePwvjucp595b7mijUfpSufInMXi0+50I+vp696uUel
XHZDpNR8+iq7RVCdhimzs5NN7Yzkq3hZ8uW9ZRcsMia8hzx8lFbP0awos8Mpr5se
J8kbS6ifi302UmvbzlUiqSD6nRCJFc9XNCw7hi5mUqD1cPWaYHkwLE0HVDF6O6sE
oLxisFP7JER+4VgcR7xOpvUPa7TPNV0hN9dBU4OYwIF22WMbrGRp8u8W3PnkCNdr
bn6i3azT1v2Qsi6q/IoyVuzs2HhG2pkcR1ISWUsv3VMNJw0TR5McN+XPVCuU9mFF
ghfHNbS8Qf1Za4mZYKONmmLuMJpZJkOucXiXx0z63F3sk3xXKjWub1q4ywUWNhUA
EeqSFj5zgjwme0dzp9xnwi03j40e3/QeCm6aDCLFcHo0Bj5IlBBtwr/Sb27QlQhF
cQibLKS+3OveQecGD5BBdKCGWLtqmmYRoQtx6Zg/l328HzumSAe58v+vI67wjac5
5eKsrjrWAWsvf+xk3d2hPnA1e3dyGW+pu1Scnf4s97Be1W7T/H2VOW3K1IivkUBw
UyyBVf33jOR4aDWFSwGnkAuhs7qZoZOuJx3GVq6tHdvl4pm5Qb3NRBv8yG2tATYB
YwLfFR7FgcyW893Tpjm1LLA9ccoJWNrTQNSHOekb1BHAE0iWVRQWj5PhVoVrv/G4
miEb8x7hkxQR6vFCu8EsfRV+/ErZY616RPaN38lDDQ7atybqw5aCktUDxn5td9TH
9vf2cU1qUxKteX4HaUAw68UEFRW+xhpekPFTk2iSogRplVDdSg1fSRekqXZ5cQ/c
InZyM9rtvsEJ/1qYp3zVKSy5VIA6eXfkdDmOvTe02oli9wIzZpTEYeDn3pU2ZT/S
U51xhgBGHqRrmZTabxEeK8N6sBa7fb/H427hZY3loAWmle4B6GxoHBcvecZ97Rxm
CWCigWTW6TSbXHF3p5MEhJ1h/rdgPOEQSL5Ip2ojGs80vwiELDw+lB2QLveZoE6f
4SUjpYCaY3ROpqnUBc/Kqnij0P4B1rs7178YFxSwY+FL/Bxfyn6edjRBbfk+Brep
SnQIRQOI2wbBWyhixI0sHyQJAKSU5T1PU2Y51SE1Q9ZlM04XuuRLICZr4yGyEov+
Bq0WoIhBqXIFeeusnQYLUpX+l9V/gn42nH4chWEcmcntMu1mnYgKnUOEFuaGELIw
fN2TxBR/4xvUneYzCAAQAUBgHFOUxYdYEGXKaDa/qLnI6znFuX8U6MxxKuah6p7L
3LOnBYtZ7/xPJkBv3fbapgV1r5lIOQ93dvbrDj34mOyE9bfSa9tHOPalmipJkK6G
XTpB1u+8THygil5fucsTvzEsikQ/8gCne1x67v3l2d0OuQ4KnwbI1CQLT4w9DcsP
LGMqQQMZfgKQynccUgvWuqcWQnjISKNj3enc+GaZfxmt0aMqFphz2YpFdpQQAihZ
pZvi+cmeIFyLJTB3cebNGBd3VBCdvbZXwPzrszheVGkzAOsUzfApImcUaQDV+yDC
SsCuiaE0TCXdcnrTjjcvxt7SY+HCS7SV1C2CiGuv47Pf5NdGUxweq0OnDjR6vHSW
KE+wQDi9GA4jWTZxAAsAdavbWbvkamV02bVsAj9E2mNHuc/YHejZtUi/feQRxZlu
4UilvSW8NkYGBQsO0gDDR+xmfZNFJrHTHFCSg84LwHhPqB3pZE62XjILxZQRL7fc
GHUFAThcnJcgSzqrUiehNCvEX1NhjFcN/1gG4oPoiB45u9Udqi5d5IBCaeAUJt8L
si5IZOrXS3WIDqi3SQM1qSlA9rmPmpeviJHdIV+RxoMA1vj7qdwgNORVOtGV6OZS
csihzrVNmLwGxVt8nZOyfGLqdiHij95PXpxrlMFT0PFbSUkYQxw+s5V083bhhjjM
AfLIILB4fAZk3jXq89BbBYBdfMbx971byJ1J0fAxkSrCWV6GvKVj7qxLkic3XxSu
YnlQJiVjd41MCg5YMyYc4F+gN0iKsqXkZapgmgaUcbAbeQw36KfpTUhtIP+UQKzA
rm5q0rDo6p5R2wn4yWN62PnXKvCi8akt3mMbPqOy8HUiIksWlU+wCvdGdpQxjv58
Z+UN9s4d1nz83LTzV94QpmTcNIXls8MkweEuNjG8Ionn8HLxSfcdS3EiRWEK/I2V
vxSBXnNBCbPs81R0UxPdcQyKsflDp2Jbn0gLuyxxQN9Bz0e7Mx74mZOFOa3mmCMd
SREXTB3TowHzvKBnkcEEjXPMT5mqq5sTRX53uOnqqRUtZ/54OrBgyIluDnR0B/bT
S8tlWeRsrMwM9jZ0b2voPhHKxrp+4RYc1arXWxhnk5sJ3Sad7E18Gw7RNc186Rvb
3v/Pbe23NGfXe9NLW/fkjoIIFihY5DEss3AeTmXl0nsXqLB2yGDzZsP99edP+00O
mCKBOLD0O/Yl0SkTPaFrfdPFKAhC09erqHSe/VtFHKVTilNXFyxMBSYIXyOoeSRZ
HUY+cEujkDfFngH2D/79dMVkK/GM0zsnGwNc4ywVqqu0GNaFSCJOmJ9TBiIsPwYM
L938tXO53cF/x+SqcKe+S+lNza6QkdKUsqEQUwfP+6NT0+6zNfw0CYVUKNfLx/x4
HcKz2WpBmr8s7GwttUuFL9Mws9t8nZ0/bsG3IDEL2uSSCpDtzGny51LNELvdykRK
tai7dWfK7POnHRHQijBdC6OTQPSKDzmzyTmglANJgv4wsv3lnPPE6Qx0xZg3Yn8c
wjUnzZtqa4BW1FjmVX2ubU4YPoV17OVnbza59Yj0w1At/QoQaDbxx72wA+PHjQ5N
t8OD2l1OEZft5BFK/Qxy8wdm6ybPprq/Czi9eF0sIoDEhiM+zh0d9uOdGtGtO0hM
EHN9AM1XSDAnqUFMniS2Qa+wtJCLhH6MSeEPUSajv14QM6EfIAt61psBG7KE20rD
JQkTUyQa4oodD9Mzh20An7+8t4zhlE9KUVWKGtB5VaSt2buBVMW6ogJbx2i4kJKy
YG5QKXtonE1yIVizZ/IKv+hhKUlwpTMLETKOE0Q+lWWzD3nANG0fiRr9zrgcDdb1
cut8s/aQ3cu10zG4HwR7z6r41o+RL1ays9lB1NZqbxpFTOSIUhoqLNszeA1Cg1uL
lvFp2n3KW+KeW3VQJrX0CyS4FzD8irOpfJIIriiybsThyTh9tlyLeyfcDsw+xyGV
d3di6CgH4vYqi2oBwyY1PAxoylEstQf40v1eP+4w3txSEuX3xWWfeARRQY4S61mb
134fyNVAS1/9brPTGaKyls7DE7Qq5hLnHwfL45+nZXYN+jxjysJSOhAleCq38CBT
Lsng6K5OMJFFa3+vaCkW50X3LVJsVq+qTT0nkvY127u6mvOm0xV6hV7nHaLayYH3
djbtWDRy9EB1LPFd7WXAIffHEBUpAz8Q17TxAVq+997E+szJZ7fY8AgutwoYHadT
vqlClUqISNVE0UcmAlACupkXhurugkYxNV2GNSjNgJK1Wh2dmwnTpfoD7S/DnwDx
Iqlk9LEIrXeQDVJ/DcAYGHHDYI8uZjMeBuj/Iq0K53KYXQ/Ddm/MMZOn246A1lfz
gQ3cDPu/j1Kr2xrYHbYavLcclx0MeRvHWs9XmNY6h/AQnXXbf2OtPwrE2GQZNYMu
bClvmgHrOO7wqmV5E/4bhDRP2w8WDeW06v5OMUQiUti5rZquvOJ5DInsEU91XbZT
6KfeUitxtLTlTsSWPTNm1dvZAOEtJz+Y/75AYVXxUFxuKpJPc+cxOkJAqV0DGJuC
zS+F51KlqD3h5/gf5dstImmEnE/SW+0qNHWxNaqHnGX+nzdDeqIdEQ3syrv1SBPD
jfQIkSdXDlPBpf8TQYni8C7ZcNmk5O0O0+zkRW5YoksLtIWD7wQZGBtn7NM4eqXv
cdw6i2pBQ3OVF42fWuA0n54N/QXAAebwvliIZNnilHprhItIJuD78osrcDM/M5vj
tm/cCmaGuFNxiCMjHGfBdHRSZApCI/JfSSZ+ZoCWKFuIdeDKNSi8XenoJe0/YPy+
tqtPsa/vTxhUrYzG5X/bI76mdthaDOOBPh/Aw2awG0sDuUjmCLLMUlvymnlUxVi4
SVvO8zqRgD1stu85WxiaTBuEs7PS0bTNipSEYFBQVTklzicrBVXma388H/sobOYP
2zR4u8HFAvhlvUkjbKmXWhh+eHDRPOgKe3ZpahkmirWUWDtQKVRG8BSW374QztX9
60ivBsF9eVbiRWj3wXuA9PRcHQD2X1wPwBLlhg8nBCnACrJr5ITuGrjwxLAWhBWc
Ngh/b8Sr+JfqJNczG0E3x//UQCKHHxn1OKNFnYUJIgVApVocE0geid2LAviCinqp
1roAzjLlXJxQcgmeiHFN2wjDEbLXqsCptiQcWrt77Nwjixzh+eyEjlUxbJuKhc+b
B9lXn6sJ7mPJTHwNxe5gcOm4Qhn9HQO70qPyPeifqyhQD73dO9Icyasjy2MhvrZT
75pjBu+pKxMXZOwrV/GEQIkyw3mWGolfkAgrI8TGbDcJXL7EhV5weyiVt2hL4w6J
6LNEY0cnH02TBTPBuL5+43ByURHELXn9aqg17QYbc5WcRKSv3N/pHEwtXnA4D5fh
h8FxDrsbbrz5i+mWQoUCw8dJjxuuYuFlEydFnTg9e0eWDg4esiDLQ3QLoPVwa/lu
nZDRfw0RINHQE+GKLPKMI7SKH78d1SS+BGrwR1BTzsE=
`pragma protect end_protected
