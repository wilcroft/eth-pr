// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:13 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lS3qgHezPCm2k7J7TRpoH+3CEXEI5m+xMHBDVLTNvfRPdZw+77JJXzgvG+UB6SFG
HAS2v4CQzSeQEZj7DFNYmE4uoWV2CsY7ysMpx66UHHUgvszRu93XGeyo/4g783y7
b+awS0jtR4IzWrtAbnyb7Bmyee3fsqyzKoohHiR6eVY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 46656)
r7n2uWKIYPgyLQdQfhkro074ZRWxtf+0Rx0D8C25LWA3N6MQD9mMATfeOisc4Spn
Rw/fYo0nR4yE3T8m22wFuNCURz0CDjKmDxdJ72iyfalxXIbMPxo+VK6+xWgXNsgh
kBQ6VoHRUFlFsiENx7Piu6M9Q93EMmyL9QRXK/MW/sQw+OzlnSUE5/SRFoJHAmSO
bK7or/agrNwGM6rbTmknZOyvgW48ZZiOr6kQh2m8jXx2w+CtAilT0BEZJmt9DWUi
tfAF4iGlDZj7MU+12I3p0zq2md7tsOaIFpa5Fl998zN7Ryz8txxYjR0CyaAHaofE
8OSxYlcXdC11bxVssEx8aAMOLLbkRq5DlbrV8ehAWp8YRBA5NmtNONgHUqn+iBO3
PcOcVtTBED3VuqFKj+X23N+tbAp4uz7zMLlEVc9hIzxLW8WASYFa1j7ryb3Vm1Xc
Cbniw35ONlXwNFrMdtW6lO1wXB97CrZgBkDXmCoSrZqPaOvWuHC+g2yp11UOMpgr
i5lMpX8/MYGL+AaM2uUNQ/RAUFy2GoxuzPUIqzA50n3KhmzzwsGvREYygX2qfan6
d0e5E3dF/T6vD0KbvmuGl8xY4M1441BG07Op4vyqJ0fWEOTbvmuetmH6wiiwOcsT
Jckyus38xsOku1Gf4Ugu1MKqHGXJmPUf2IgQ7WTuHcgx8dkrskRg5qkw6mlZMjtL
qlR5PQd4Xxda9CKT+gKuoPB9ixBmPoY/8lzzHpoc5zT3TQu/hMyeHODTvbgd4Tdv
ooB79avj9MU6XyuGLmJnrzDZWuQ3Uak2p6xgUj6w2AkCGEjIMWKv7+ZiU+D51Kni
9+euzcFwCnMROebC5jQW9q3pseK1Qomf7qCNE98xWD3WtgBShJe+Zmq4Sf4TOqDU
CVj6WI03T7uFtPP/fvxuhE4DWWdB5+CzxYUfYf879D6+gkeDQenQLuw5AYDN2aS6
BaburEuZhtxFS99PaJQrmm+8LKF3YRdzjfjG5Si7ObfHUyqCExFw0y12IVZ67Cez
sO4vrJGajfmDBqPu19s3kw+7IL0Q1YXSXFqeqnLeNIoOLIrxp0kMLbAPlAEUVm1R
Pa3f89ExIEDQ1U/itZK7O/FlvPNNYX4hy/wK2zrGQ7MuWmdV8I0jJHUURafRAj32
UNTKgjHIl0byRAtXRic/uW/1F7vCn9E7XA3XvqEnJ2F6MkzgsHaWveGUTaQJbWKc
sDlMU6ZzYj+jbig6GOfekBhTIJ6UJTbM6PLOANkMXEM40+FOP+Emlh4NxIG4LjLG
NI1uYh02nOOFVJpOblgUT9ocHVPwmJaeEs2LSnAGVs4QpnmLi9goAHFRfmt00AZg
IByqLdMPrgnSpAj4r5Aaxcgx/6mt+X59/uD8Qao+EjzCEPChONCuAdHIWPzVfUck
eT3XdziDAk09ZuQPeWu705BsCTQqhOjbvLzDYij607ORoB2E1DmKkTb9p98wRJet
1XkJJP3VrBzB+Jpupc1HoNmKMitMDOfabTXs822zM97eOILCH5DBhSZuOahSu+jL
jWCXWKvOP/ZcJzcRbUaPELZshbNB5zdwp0gbo/lChPZ5Fd34/Vh5EFNMe2Cxxrev
zZe3RTDqhEN4+2+h9YI3+k6zKRDLdDBJBvWSWwrgJJvNNQZX5mQXe7qHnO+aZYxo
S3FiMV3vlO/hPgSBRqcmsGa7JgZ2q4oHbdQDisgTHGybk8IXeBk6rpXVTh6wL5rN
tucRXw/AW4ytqY38dMg/hDaiI8kW/trTpOQg8+z+aftOGheCLrNU9G0hAatVIw2g
mV8URl9Yq+M2tkmQBCyGoDyeZj3nD9zQcAbmUQEoaHtCBS1JADeG9dm3Q1d4NwAh
AxyXuWCUF337jKHVEOZWc8wvix9LD3vLi5se5ZD0RZYb9nqPpb+lBh0/sTVmyfbP
xnTPPJRyKZZlycVKD75cT16J1iy7FkqYxqQMdewGUCL32EXcP2eccY6X/jy8c7gF
+ObKICU0KjOrXGtI8xQLKrKSFVfCs2iXKyvVDcwEbch3Ba6FKCjtdQdgq7JgHad6
rD0qVeXnMg1Lue5w8cS2GmJ8HnV3aMJwfCx4dlNEQ9NTD0iXTQ8rUjGhBnIJn/EV
UM3dd55VHjNo0+qN1+8CKXUZU7VixXRoIk9uNaV5JgFI72aCUCBBDNESrx56cLeI
oJgWsrI9nqAJKRSwVLaev4GVcQ/LPDOx270Vl2fLWYzvVrgp00L6zSLUQOBFq/Ss
vQa7f7IgJ9e17oJm4/jwOU88xZ8pGlqBlZ7x45MKDyvDfoY2wkmMWnkhs2W+7mV2
sWSoNICFHHYwK/wD5Lg8PiuDJymD24S8SKipPIKe3BL1aj2V1/rCz2beeDR/cWK7
seUzXRmsztERWW9Zycgl9TTdTuV7BQ6Epoc4zyfQkyPE62wdUqhd7Y9GvbUa1RbB
kk12Hgrpr9DeHqkwit+npIOxQo3aI73U4LnPikb2kMO3sXjTeztu5ia63hgWRS/q
H4qPXmfnOXN77GSBoVAsoFtyIkcvJiN3Yjveu2VSUnn/VZfWfoCz5XE3yxwPNPO+
6JNcpwl6UbW/mKQZB4iMkU4ALV6YLvCLEYIz36e7Tj7b2cYIwc7q0vlsbKTZVizK
mzdDCLyTOl1iwJnXzFsGxCvb22CHXGPgMkl8tP/b6O3+leG8JO+xALM96nfxPwEP
d71lXpuqyN4xSx+CN+WbqK856Unv/bd944pQEGi+JWfJeuodKF+2zT8u4XYihSMV
+ovyGuAbq57zP1pfWFjbZHsHKN0EuSF4duqCZ6zzB5bD792IadaZJ/61EayVlggS
jUbi802Z0vvArbpyOghbE0YbPKWKa7zOZ6my9vx0Yam1ILAwcTgNK3QtZc4YhFEE
oNBXffPZsbnCiuYk8qK/5cLkWfMq/Rvlnau2iSQob1GUe93kcNqSrIom/30g16+2
ouUC4oTzX1BbYVj4HnPxbyvOK/MVCN1OkFMTsu1chNt7UhErutoTzd7nir2Jflzy
onSNcxU1ZfadWjc4u84ElhBnCwPBpa3uOkGj/Fnn6LjXx1VUP8Lt4Q98HRDfF13o
wrU3q+XOlR7+25AG9inWHUxa8evrlR1AaXVKDrLP9yt0Ic4rnY2k3a35dRuQW4Bv
j/pPJJix5DKZ18+lsr/TRBKz31x3nC3KocZVKjNIgR9Gq3VaWvoGD//sNMblhzhW
CTyqIbF/aW75xDdENeYc0xUFkOW63X05TYgl7Xws6iczBYVB+vaTtV5lrq71KLE4
ceOwmpE3zHGvn6bJYSPkl0o8vVOhMblBPh0fI6QWewNsfZlsHMi9UUWKtm8/FHKr
OXfmoYpeip3nDUAaQcVd6xgz496ydNW7011MLX+03vY+1BXuCkTZQBe59ue84XN8
5UMCNuVtVs08SviPGuUj5Cz7cojUwCiSATY+lsmB64jNbghuUWCs+dYQxAEMTIT3
oSEiB4OTAOCd3uAyBQVLyitpf51lduQMOmn2u14uTnYoweskQeP8G6CwAdDW/sqt
YRenXPVf8CK4Tel46XHKF2+cXBu5JuJdz7vbTDFMPuZl0ljdX26w2akN1bJytrXY
tIVpc9+RbC9BOzIhYiAF6tWlEUir04aT/TiGQ9jvkYjudL71swbDVNjncgogrHty
DhqqB9Fb6w2tPZFDM3OKH/Pi4VJ3hcQ4rQRvKom1L3jSDeLrcGbQqdCTqvckOyqM
TUlWx8mVykcr9LTslpJyDDZQcomOclsMbcW1Z4r5ZnnF5wbEmkv2s1YkVR2LoF8A
p/Gpi738Hq9m45UYfje/GZ5M2Lftbcz5XT2Xakvl7FF1LOtjV16IuLAAOr/U/Vlc
1YBxWA+gdSR7dJzlO2IF57GQPEpaE0n8IExfQPxnJ2qUv5/BUHaFn/40/pWcu/jL
oeSTY8S/Gk+8bqNhtx8uZKfXynBvcXd0dCTwQLtPUxQB/dgZsit/f0Sj+EoLEvP1
RAoInHEFazxufqIYRu+S0MNnDo+jwFMRj1ciYXOuZeBuVUJYNqhetpPOviHz27+E
scTDDgxPdALjh8Py2TmKC59S9rpRnCPyNQhTDcEN46d+bjwzRXUAFUPm+Czs8QpC
tZT+Bl9KTHvzOZzTL+tDgYwAvXCtATaRKuxOvrdSjKuZh8mwBx4Y3OdWQS9QrccC
OYASTU38MtCPfl0F2m9eZ16uECKCer+20tWMAq4gmkxcJIwQuZB3e82KgavLkdcV
2EvqZE+OLpaxNx9H5j//HTnHuUtS2tTwkN7B+LNtnXkyszzXt1euqZ4s6LrU+4ib
cP+USuwqwYNGx5Ylew7F4SmXmXncn8sXjLU46HhXfZ3Cn37u3qoLS8dYbuVaR5Oe
VFruX/Gm++/vgGxPUNaliE4Dgm/vcKYEVKHcx1Uv5AkrhEaEnfEiYbJTPy8Wcymw
+4iF7fk0SXImrJSeRgX2MVW137wkpQqdZpVh/jzTlBDYIvoLdeXdwvcvse952G8a
mlJbkRjsAs0seQ9HtK9KzMJnimeFnixaPexxjwCJ0ddDOCN7kSYZoCmuiI+8d3gB
ole8IvhFkBVzmhZigUoeiac8ZsTd88zMN2Lp2iWljtI3JIi75OphxeDTmoZbJiok
CwyPWbqJXBVcMn82pmhZc+9wYeQnEZwfR7WCnudhSXCmn4p484fFQwzvePhmjEK5
KGXHSR170wdZ6A97KOERikYG4qLk3Fw1pgKqwUXq51p4KsmGLDsA6ibIjhMq+8m+
7mQJKzZJk29u56QS2BCQsyGXvd0cwUQufEjnvOsjeF2Elh0BWRQPEic1Zq7BrVAu
Xi2MstVA1rmtN/li9231iRLEWZ6BTZNU8u6a1gez42KaIk3XCGGhs0/tI6m1mg2U
WpqQuw3rQxIEdm3AwM7SrMxRoK6+fN3BhaqATQ/H9YHXi3SC2Ruv8Pb2cIQxGWBX
jrybS94UFnXVEDugv7zJDpracktb9nsoGNzmOMeT+tW9EeD8f8ioPw0lr8MasTV6
kYDVjmHAX9ya4br8/qNQfoJW5tPt0R+qj5Fz4KkaFZzexZGLuBDjjwxGZsfPTlGB
Dwjelw3+0/zaEV227Djez6UpMI2sr4hITHeCw8yhYWemjht7oNVMWZVvIGhaSvgD
XsGWP2AH01vfQ+Eas3Q5wdsUZUGkDbxR4tulKcqySnU7RDh+dRmMeMHuWFASKfnk
Jyf8+Fm7E2TSY08mqdud6RVYApxGfhFBLUMoMeCDwJXzftCfjjEIpeAwO3CKTlAb
dGRtdrPhBblfBrDkNzKxkbhdn4zddw463ZMUPJUQcO9N62Zijb3fI+Mot52bUkny
+Yu+MItuK5kmUr3dk0ceZt+HhUoR7KiJ1MpaCsr/WvqmkTM7s7xVonBcoA2KpwBw
jF/BsNwWISsHsp0wyMoM9GC3PKlkmDpIKaTWzVCbQphmHojqgOsK9ach1MsOGx57
7ujojUiXHLxaHV70J2oaHzolNs9frubf/0LWW0LfiSFiuESLJwNsqOiNaWxjnznj
NHNnDyGm4+zrp+ZLSYaFTeqHhY0AEj1luM78aquPhJjaC4ZAyhsrsHYz3anXyjZJ
JZygzx9qG5HBHPce9WnlL7oJH/R0jwHYBmUWbLj6dH/+RBKS+y8EKygb3qIBf77g
/kgmhjboh5Od8ux0pBo+0N7K7FfBgEBH2TNfscAANFrslNjxc2pjklYYBmnTK5kK
t12NkLZ4Et8HM/oHbfvEWM2gh/dSG3MTEMfLmhd72qeWEXVrHD7lKvFofhpZ7+nm
XELk2huohnVQUesGOCc/x3yDAjW3ubGbBFmjnu3IaIR0C1h0vJXi3GvbU5j3iods
db9NT36VEDnFMncHTZVXmr4iE89d2w2Xew/idb8Po/tBTFdede45Gcg9gm7paHCW
2Jftl5NBCFj2jdJ0Hie3roR4v0+4Zc+7daSkN1nJoc0ggIYrw0qJkFbEC8Rh7SXj
GeRHA0dUu8cNMNvqojehtTe8kZm7Osi5nfTzARzplr1/vo4KM/LYIEz61veH/uRK
4hODVuoDJX3hNRoYSuMLsl0N97ZHZko+AO9FPFzX9jNsBEV4OfqC7Q6uV+oifxts
bBGzVA1WBuZwKcwuJmGnWpegsab06EZNZ+M0K7/YGT75amlWtp9RC1bA9d6xb3Uc
tF3BJYwcOHMzYH5Eb4V6nlJtK3m7pKTQRbH15ZXVhvL2SpyFsHHCKc0chauoGqJ8
x6FBAfgV11RTH9+AYw2XEhVy3kf6MK6Hb+CBFY02NW89udVhTMOgh2p9SOFEEl2a
3WheXR/LOUphq6IPRL5OvOBiClPtE5fc1iQ0ANtt5w/2V2cOqu5+RJjU1I5cmALU
HBSeSFdyWafpr7WG2i0g64nobrZXX5GgsPonxWObY7FeJxPe/pRfRR3/YlNd+rbC
sGCEHccuPeio43X1caZS5/3eVGpmxLq4dj8XMl4LbkclCsHxvszemkSrZZtrAvJJ
BDjoyP0s+hTN/LENNerGrg1xP6Nt/0QbwyaHczYO3D78lWGcfr6B28OWwYR+inQA
aC/KGNiLW7WfFXYbExRURYJSwI9k30E1KP75GON2eRC7IAVazAroencZqf+QY04l
p6VLaMjD61ymP4h50MMpapJoVyj5fS5JfP9hkNWttcveELt28rLcjGMOtAYinA/B
IsV7k7bDJsVlBAt0dZH18EG0QtzEr8tRd5pXOVWUCzepP7P60MdvS8nsPMRvwROB
VZcpC1achOqhUJi+vb7czw3oE2XRHYlZk0jLUruLwXBoeRd8z3lWrEj8Pd73Ho3s
JRwXPf1nctA9siL+lrOZ3D3aWKWdcEPHLBgXxMTken1fft4pyBMsV9ue/RVAL8th
SWSM319F1kC3MWHowdxypTbDsx2NbRlYGu1jK0tSELK6QhP0tRXdj0ZR5xJjBsYw
F4jQCX6MwszFWjD20PvP3IDZc/MbDiy71mDfFAqYOdtK1j2Kq5UDpYQ7iZECwDvO
WbUtRFkOIa7sghE2+4R1w7AQh9WmEVRxKolP228QvxHJZlAH889uOQj+T3wyFVMV
D8aye4QKI5j2ju2fMAZQHNODcZWq0BKEKI5gNZsyQarUezkMmRPjSHrgOiPVu66B
mkGYAj5v5kYGbHwu/VeRJBDcZTVUq1nq18UZ8X6xru4OFlMRtkfGD9y2jI7i9TV4
4fTIjwCR9CprPy3lBoSOw8XWNiQkCfPSrztuD4+46NH7+JSgyM3OTbFBK9QFlfiJ
qv09m6gH61t8FOevn6cEpQsunOPe7J8aXY9QpudQUn7MTZ1Hw/odvDmpG+WHd0tt
N3LWslCNX5KL1YpTqiZQf0L3C11KjFn9rF6DjbJ8kJTEQgVQ+buSRJmTZe+iqSlX
6rs7insy8PJFkMJr6Ssy8ixbCl4MwxqFqG8BAChsBNwDKx3qi0BGvernGFBix+MS
6B3rQYoCc2JV+GwmaU6Qt8pbh+LsZOPCXVU3JFZLu3mfGrbjeebzogfyjwxwv32E
lgWgbB3Yuk7deH2cq6MuW3rjgqGqNgObRVRcg/hv8wgwx7FJiQyHjnlVPrszyb2r
IgO8WP4zoxhtmrT5MTVzq03s0KuFJBmJTxD7X6+0vvADrlR39j270DAMF221gKnO
ufi23SvRhpeKUi1tHT0jnWT1Z8WhccF4dx6HU7M6Fo5oRiRNUT3lpqDjLxTljl4q
5/5/CYKfLqmisfXpIgupmtwRQRju+aAzrrcM0MUcvX0WDXKg681+i+B85m/Z/dXL
inN9MDD3evR77DCGgC5RRTsUgvL0cMJG99RV5mr4Pm+wF3Bf9oKChSjQ5DNDFHNQ
9UEFdZ2KpOYEwZla37gYAVZbKZ+QHhBh3Ofil55hkSDtR5aUVPE3tAFztQP9ZNeT
qI740hswqIzsxCzDVdEWLMHjgyJOA0JcvzQQCeOVmkO7hGm5J51o3XjUp/RxXN0s
hD2Bdi78dHSKtUDtf7Vr3wGP5e4jarZIlePYhIj+wbkKEXDAXEMXhG68un1w9crs
2FX4ruwxCsWKPF0c9JYr++91Y44pK3oToBCEBFuka8KZlPqN4/RFoVWgBqKYRBnr
Q/8We1m9ej2255YsCmF6xIX/wuOhUbfDaVymVe9ij5fUJ5ZMMVk8kEem0KVZyWFt
IG+GwU4WQM96wUpMiiMmJJD5Hu7Maykj12WKw7CRscwgkRAO/EVt8MolHi2EkOza
GLngIKEoKtmLd41u8XkmCkuxVGZDmp6xZv77+86/Rsw2oGYfkT2ISgSEG4x8Z29t
bxqmPzDlpst6ZdcsO9jOqQVtVEJ3LyR6fQt8PQ1FEdAFTSDc8DYwxK020yHdC6f4
+isKg8X+z2mnJG58A1k8OuqXYwX1yXQ5/YvadWQCNtgB5s/QikEYK1utqoV6hqYS
7eOCf/5laqDlhDjSKQOmdG6nZPNCOaG2o9EaCGSc5LilTpdHYFT6Y8I6c/a8J7sw
5CrE0YgNQT8uzxU4c4zmquZP7yx1TPcDdNEZUgLp001cC6E8FY9LvSAvUZAmk463
PNCehPXv1TrFPXuCwVxDUycBQIUZM0hkQbjaJVwy3jW+bM/w+2qwC0vOGLVoxAby
ciWw2jqLP6R+XdYeRFgcPBR+AQuaZejekFFFlKWnctDzJPMvwMZF0jynR73TM7No
2XZX+vJzJ8gA+lSGUNnFqDFYU3ne1NWS30beg6vA6/fimscQy5BfC07lnR0mfFaZ
JocdOj5XA92rhUsDSj34YpN9OYLOs18bUlXvX/R/x1JrGOoakSOKlsZMZ23SgPJ2
be1zzwLd0H+XJLbO5ISy5QETJTh9aq10Vpp7faRBixkfm/GSiQI0G/T6/X4UG6Gl
Ud5I6bWMZWBz5pW+7l+l5dqj+y2GunavMVrd9rdDzYaelou7bv39+MdrrcM+nrGN
mqFr2UFT14mwC9ZrhZTgJla8iNDGM0J4U/WruXH++IcEPxtSg800EZ0prlbOF7+z
JNUXYn2HVqlBONlAmslqJPmsREONH6QlAZG0bgNQmFVlYzPOwzhN5KybIEnwufsd
mIl8zHpgsOd9j1gUx2OChEnIX/m8umGVC8m8k5xtQBt/G3ZqBGiQOcFNATFZvJss
Mbi4lVYr6TWQyqfLMUy3cfRrmEnA8i9aedla1YzyvMHvOOmHCsb0cAdBUtUUNG9b
2vj+Yo12F/WCj6handJFl4tCs8HjnYt8YStHUDnxOT+Ss2X+0uwGGaPdYcBzzGNf
92kAHEp/cS+B61XbgtZ4jg+9oHVTzZlGlTG3eNRulrGQtVpKfjGzJryMs3Sbn1ip
R4ejAkXopAmWPo0xUBSpwmhkOYSnbkTnaiPjGWBKqFpzAuoS2x+IWNr5mrUyNniB
IwmRLEoqyy1cpSF7xc+Ih9MN6DygpEcpWKbzTVvOA4RrZjd/flqcTOK9+DicDOOW
qBS+NcgS3AdpHqXne5dH2+7O8VFEA2UHUBrR3KOmJXsK9o19eK/pGf/8Ht+hdvp5
T+SYieg3TMYiyZZ8XAr/Y2jdQF+uDiAHhWHMXDbJ1HwGk5NdR0Fl0ZpuyoQ5zFw+
9JxjlHGF2WLsbaxqv9WhpI0d3/G0cS28qK793rwYPlle8ErD7CO52cpXbJ2VQoSZ
zNeocNNdcaEOIAjvTTGK/fhY/Kg0z1kCoOcCaFKVYFCU+yuSDcNjMZQnPsPUVcV8
5Sl8d/myoj6Yk6AQIk2BBDoBKWR3ua78hHc3gnamA+BfprcajUecHP2409erKN8g
0nh4Ji6S0ginFvxp2ueLOhqp0gnLAFKIl/Ptt6mZNmIZHU0Ofuf+oe28GquwNLa5
bcK6ULIuCXi3SKIeabdr9+ipY6fGfrMxWN4APJjlyE5U2INbaESkP8jXdyu0yojk
ePAtXYhqIU4PigPCnUFaT5Gtrt7iTFrN75xHCHE+bkY07r6a+PJVcdib+coaPSUr
ZyRrr3HM2WA/UZlVnbWcnHlTzP+yCau2+YYvBmsyUHl6gKqA+COzSP8gkpN3pK/T
2dhRpPUVps/XB8VCpYHxq6750M+JO2eg57cS3mqM/JSmxmE44xDXHWTMSpXLkuPV
1BPeD4ATxktAc2tiGvkE6Sgk+iD6RRfPrJlxeK4QdIl1/jThiJEi6PRoMvVlhuaW
N+Lq1DFvlXp2xpve2vW70pKhvKN5pBLt2WzoT+rAEV2Lyft/MnNT4dSfxuzlfNHO
ZcP2CWZDEQat6lFNVgML4HnFphU1cqQk6+KiiG7xs/JM3dENLhUMOvjpkONSYnlI
QiNuSfRkKzt8Gnsv9tmaNz5K2y7ASu+xAp3YAtUVjXig/wit0xqysRJQ9/OEi755
VHDoTcQEmOM8+an0T+qzkJf02+Er4mWm1kD4LPsZp+pLFuiru05J6+/bdG/p40MG
kG+El3sNz4GcppKgayRsWQyO2WCOucMlJ+NJtM2auVGJ2dDPahPYI7igZIyWwBHt
YnR+tYhsI5GY+IDw78wbtJ8EpaWisfycJWfj0IeWk4dJmp/fmlqutDVgW/daQSy9
bPUZ1xwK9etmw/SYBSMaRTlYEKYOWmU9WVsQ+clfRDTRnhpn+CeX02AVy6PCTlxd
KXtQ5hmxLqC0ic7moPsNVzJwU2eU26EVIOzScuqPjtTKl6iOKoIt2YYihPwSF8Wv
Sz6mqdD2hXnSy7FoaV9Wk9j8UgvDi/drL3DYdCOpyT7o1xhhIEuZ3p4nYBaB+Dnw
o1+I3PI8j4ai3T6kxsCJKRYC6CI6HRUq7WLYp8EbxeGcEPrUzfqs9XzWN/wVWvtH
emFaWfMJRtatwytSA5Bm4BNXUiokskpPFDTyoVG7DukXKAyuWVFvU9oA5ucz7i/6
bLwVS4Bau0hzPe8qniPS2qA8irdcfT3Z2A2cC5AguDpireSToPacUis2enIA8e5/
aSrn/HfulWtRbYI/MOhnoSJZUT8fxb2OqlEPSf+AB/R/Leuueyp5LOtQVpSV9ROs
ZvKDNxV1Mlso+TvdrLa49H8tiPZUVcd47RMTOKFcRMRU1mhebBKj/a9qoV/taPty
eSfsdpVb197lF+okz3aBWeXuu7MC0+nSi2+hg8QYFI8McZ/r0w4Df8ydv+XG8nfK
Vfjh/XDDPOu8QTR+tPKqnzjO/bOwsfJcuN8RXO+p7ozPlIRGmd0G0PtZZ6M87FnH
XOL2hYQp+IVrsgaJPmRrmY8YcjN/TQ+rAknaDJwYOKh5R5SMF53j1NU6S3ahwFIy
v3qo65gWqM5EOtJ/i/O8BrL1QTULSmKoTOZRi0CeJ+wHtDPVJQ0gW5PxEy7kF9fC
qZwDtj7k0f60Gz4N0wtzYiZAcPUVANCyrArxn4gOIOBoNOTEYKzmtvgwobn1JWD2
3xkavm19Nq0DZ8eXKXJoi13j18iNwcVahGk4eO7+FfNkZT+vLKIuwzEyixOMMrYb
6yBVY4Q6UAosZtFDmvI+AnuZiOBNmdpSt1ysxysdTU0ujlBABdQw2UrHESJWHeiX
ICBONrosh8WOLZ4pifmm30pll2WpvvFWVCUQadKAn+47AOHo9wmqQVhUEJfuVSVO
tiew6zEGcUXwxYhEG7KSCnDzwQBnoD1Q/Qh6YLWEjHGKCoa/a0D2XuP2RoIyiPle
FQeBOx4BB0caJJWj4ywA5WRmluGkT2gH0aQDYrQvRf/DAboRJlS+alSq9CQ1r2jY
2Qfwc5Vg41uzOiymhr8pJZWQlDzr77RodBtvxR9csYBIeYazERkhBak068CZEhkN
D2mdzObKz+xQfHGIeyjpwxsisLqGFrmiqK9DedMdHep5W41Iu8/vT5d9aPYHdLFi
Dv12+6TrpUibPRBtGgBLwdpHW6Unx2PsXva1AxR1bgvZsXkdlcxUHL2SKUbKQpv8
WOwlxqwfMHHOQRmTz4Yfg7f4LMVA4m38u3XBcYX5phfowIXwDTeWLlE4sqUSdKtQ
sw//rZtV0RKrK2sqG8s2T5KSXV4XoIF/uFePeLIla13Px8IJHT283oR5vuPKJqll
jieS+aot/rnqScIglVq+Z9Woh/h2Ujx70KJmvxRf41BE66cynupU/WmdeJLea0Ig
PE2z+UmtflTP4a3qlPZy04iqsYBSI5M4H53CFWtCTlS6XSE6hzhqlYMHnz5S7oe4
C4ZN3vfoknI/yliNjdnFZT8wECbFlXQEhfCmvmDqEJFKWhCgZV+qd/0XUcpwGsZe
RNi/d/0CQu9izeFXbbtwBj3+RfJe5c1vEHXtK7h8iMvSdJJtSFVRTJYwEKMoIfwH
2pFhclyWQhD3lRQ4ka3BNqPKbfvT5sV5JHm0O3yoSd6KhD8d8NZZhb5S8IlQSU8q
E2vc3PEnNdSwVSXsClSSZdCXXz0j05ktM157JXp7ORE5gZ77kNOafB+TdKqhR1fU
PB5ascwFDqUfMFln+Ji/4JQQHBgZkB/fq44hU4D7Kkb36fohn33Xvamd8s3/E5gT
fUCj3b0w78nsdA3zoCdU670nh5X8hV7NgWWdlkrg659ofdbxQMPbBfdwijpTfzEg
YCPybE5TOs9PlL6vh67HPxxn0ssyEp4DoMGkI4D5EYxcxtPUJTiVQjz57uHlj7kz
hdcT420h70comldHeEg0MNR7s2cji298xnoWxvSAQsup9hjLUZxCx9SMu+GdHaYV
02zjX9d97DvtRpzZ//WkOrb5FXsfSSCl50HSqXTtSPZNFLcGKVjquyWEYMiHqsxw
LMXHiHMd41fyovMF7ljYgS/9FzrxItFnXTR1Ypc/wVzN/cydD6s8pZ1NgCmQ+y06
pQWWR46jSZBlWeuPkv5pbInUB0K9/xwFVNyyW++/l+ZE7zm0BgtAHAoimzJetNiQ
tApb79it2QdCiDXichh8jVH/pRCM4vYv/WDxOr3sGtH92IZ/g0IfrLNGRUFfRyE7
Hka0LpGlplNR1vaAhlRAmSyqIlUrZcELqLc0HRWhepgoo9hmFMgjE9M+GKbFZerP
c1xdb/ws5atbnJjNBrXIkPMt3lvFn0R7Fs7gvPlrQDMXmuRbXl2DMElfAEuhsdyk
z4kVqyQOJHR0zHHJhhUj42kCO2EgsWj5OwW8pauHbOrLhrXDYU+zd2RUZoI6TrGV
XeDr65qPMCpPMJ/GnYuCarRX3xWOI35cNfL/bXVzN1mbbQWPnTQD1VFVt7VSfjgQ
rQj9C6oMIstbLJDdXDZIF+fr2mfcLw7qun4ZPfYHQSp5vLRuowMl5JMuwYbwf2OT
2gRpbEWScO0EKScTSVaSC3ceCAPAS4XnCauH4T3neOYqV7ewoFZ2w5+QW+u4IoLE
s93oIth6XsOLQgK2x1U2bEyWin/synU23VoaQy1zMlaHzn1wZoplrqiO0LUaWV5O
mb2vbwk1m4MW3qp/gOwjuSuYZ/202hwxmITtkz+tiLJH89oHUhSxpgB5RptPLPeZ
xWmjM4k7WGzaUnLyhoSNbQYfPnX8f+eEKgjJ49+AUpydLHuk0t8NUBt+dLa0OHkw
EzssIN1Ri60V7SyBtVoKlRG195bNIjkM/4DVrgc/zzW81rYNPR75v6yeHgvTVf8+
NgBmbIv+Gl+2JxHKdTOtsH0IEMCE7byn8hALJDevoM+D75vMlxngQ7aXLnlGnqwu
9EQhh1Xe42+8UeBzFL6M4885dsknOGdAfdRedzvu48/5hrVLjbQql2tselJTAUeZ
wjyNwTFLJm502tskQ7ir9U69N+QFQJ5scKdgSm7JZF56s8F/lq2p+nDCiWWWnR+t
WTKka7V+b9N8xtegW/Ve7PO3/B9GGMegmNENZ7qHWTvAclEC0XHN4W8ZSXMH2ssJ
FH43SfzKbPBXN+iMzVdU+BqWvlZ3udqC4nwOHayDwiog9ohq7/GKpcIHONoMcidh
5rsXW40y/Fw0gFSj53tuKpUSLkSHVBZj2f66vpMxwbLvnzXBTPRmo8op1HnDWlGl
fRW7gLwBY98WbAr0ZyyN8tOLS49V+KnCb+gYevrzDmmorVEFU0Z6Mmnr3D97k74Z
Ssre4pdvtVXwlvlQBTNyQnfipDbDcNske1jjXDqNAlV6jblrkfbHdqkq55cjcnMO
O4oGBhUoUHUI96UtDjUPqiI51zmksMjdyo3JiJ8CKgtczSdPRjdL+J/pSXKpBt2t
bizhu9s2qnA9uDnBqXZOGv5JIBSDXuhMPL5uqigfAHYf+4LEslGetodo6vReHakM
4+JSxNnGh2+ZU1aMlXjrqsCdWpidmKYIC+Vg6XkGm4jERH2LHC98J3Y1+bqtSgvp
mby3qJqTbF8FzMMa33zPTZlT6XrEw7s9SD3yrmCYAnEUXai9jD67Y3EReTfM6hqB
diKreaGlDys/gJCzCRWH7TsPrUipB6D34/SBVsz+W6Chfl8U5Z+Rb97uhdsB/ml6
xfnrL1HwUuXkK1IsYfm6+KBOrvnHEsmZoSuNNQLEgXYZng/GXlPxO1IxVXaSXvy6
h9bsIZ+9Ccm8j1Q1blCoTWkK4BtqL6PGLfjkAl5BGqYD42zZKpZ9QCXhSy5Hd70n
du+bMiTi/Eqww1cgwj+iyfZsKeEQ3pgVxb0Bf2A45V5t4Y93+CBT8bH5ztXG/xJw
kNVdZOW+/d0GU1kmLGlmO42b0gqNn19xyXGhSfeWzrBgL/c7ITM8o6WsbAYIZT9Y
WrAb7LkbYuJT27q5n9OO3etNlsm4yus1opXDQw5ig0Vggx0H0LKBdJ04TD7JXuz4
hx6r9p0RliV3ScnzYr3C1K5cnBdlU/sYbR5LpnALPtqJ1BUze1gZD7E9gn228aTh
sTEX/Enu2Q0Y77OQx9bUU/w0BRDwxxaIoE+qlWw6todXsG5tIpwTN8Vm5NJG+Uq5
Y8pA6JJAI3UQWcPNez2xS8drr3kbvWasRTitCl8VZPZeaCSDpL7+0aTEwBeiMOnA
kQpyWGa1XfS5QTR3UEhcwRLF8lVAzUX9N3DvUq2tP8ai5W6Ym+CU2OCGuWgA3gjh
mFrNZSu396uHIMY1o2rVwvlDWR/GAxqkahi7fVXEVjQiWx7D4/zu7cPJYfMO8nAb
CReDp9f1quiBrjD1Pw69pSNbV/DyoODqJb7XSSC/Da+fHucHC2J4y1cBwXUQrcwk
zC23eJJiGhfipAgslLm7hp/Atg2XWx7jUxxBqJOjhpw/1CqQL0FoQqyRmoIwSp/P
cTzFYwXGRQHs2yV46wPIFgbh2KoD5V3p6t1ETLUtQxKatQyfqN2e4V99BidKmdkH
jjm7NwHN+mfosBvS4CGAJ9d7tSPdHT4PRo57RqrM7Hlt4fWwioDrBUxwpljSpjFf
5Dwdl1uM6MRTSxbgGEcGOmvL3qbgqpt1ii1meBEkdIXEHLKQvwTVqWG90HAr1Hrz
7qR78rNikL02vzdW+/GYsy5Qy7qec+bA44MfJVs0u1ecZyDLcnss9UmlQJQmnmJu
U0ycd+u6+LvLmA7iiBBT1/PWW8h2ruhiuclfuyRwmyXWsqMPPjjssrpP+R/rQZzx
SdfSDGvkXX7Yd9GG55sA1F/W5HVgTqqWgK1e4bYpVjJ67REV7A9i8S0FFv02FSle
5y2auhgRiuGgOLxvAc81bSrTmIpiipsWSJAKD+KsQjQTWfZgbZ+SQKnege5BHFLC
Srqp55zDNXJH/wZElhtPxvArlwGLAJZQVQAXE9DcDAt5casFUrC6B0lm4CPzHfyN
bAzUBpxQg4hQME8mZVN/kXV8c3RrZBSu/c+ySiiPI2Zl1TBq2WEFiCKr85oWueU3
IxtX/o1kTL0PSvhW+KgolsNgb1mHfJ3aHeAI8MH24csi8IkYow9blUI41DBI1eBx
jIUm6EL13WWlNThsg3G/+KD8eHyTyn2kIblC9tB3fnNrcYYrga5gdvQE8m3SlKG8
OKY+CQtNlGFefmywlpXNOGPsD1ChRqiVy8sc3PN5g0oC06ewbBepdoLOF7up50Yj
9QBcRiJqAkoFzoLDY3E6IMU22RFMad4S4641maQaHFXvYRNSMwwUi7/QB+0Ud8G/
1zJmGneUV/E0dE8MuO2GCtEGuOou8/2O651aQcQIsRwyRpDhshI+Y3dfvzmTp+2j
rM2aqiGukOn6t/t93z4TDCLDHzcUtt+65NJR35oqhcm6h9y+n9Jab5YzmTMAu9gU
xtRpuO33HvyD3Ln+SU7eOR3dYpjMU3nOUcp4X4+Dyjwn3m7Pus7+XHqN2guBJ98z
btY3tZsL9rbe0ebC01rtRg/TIdc8wMHL/npAMygmU6Jg6pkXY7dMxBs8VuqR+bqh
QmvuJdyEM62ysmV5AAZJXZzBL3Wzx0a/qqbWaLQURTA0TZ+2oYEN1aO+e38BwROO
/jMKl4cF1gMWmJWJBnXNLnqvGiaLl1e+3ha4WM3H1baNqFMgyO2Gty+wIEk2n42/
6SVGjl52KxDvkg1YyLAs+0c/rVARHhLz3miCtlDOnaVtG2PgZ7oqhWxI0ZNZp4l5
12bw6tcQxFcBD6dKF8r4ZdpNHZneYkGtjMHqlnqiOS7TDV+1HweFnjSAy5VZv+od
kleR0o4T2JUXuTjvRkDosOwSvVpuOUOdoHKeLG7JNDqGHmT2SQAqwYbY0SAuo1qU
IIz/CVNSaGLZxAMdsFbCnwIrk0py/rZBtUkm1AU+fn8CixcFHFEMn55xquC38Lqe
yEqtUQesINrvJmpus4vGPt5Jbzwfg1xDafGtcnrVH4YAaFIDMzd3sYH7+fapLwIx
BQlSutllztGlZJJQKKxR9o83BiUfBi9rE6f4Io3JcQtQYFnlHhQXkrKecAnUAweS
FOsEHiimRrARzFBXQvIGe1NJcZ6s5tRVdcP25OmrwY+GP+1FHNEDZwgHWZzsM26+
6HSY0zN1xs9hKJwhYiKKJ+h90v7FsGuT/xAq9oLSe8MXb76BGHv6sJ4GbnH5Joqi
CvjdWX5UDSyx1J6ns+BaaSFx0BSoxQl8BTtR5Qs3XemZG5JcfGo8G8wmFMkGskvS
rWOyQogOv1STpM1L0gUAKPQuzUJ39BCIUueto9xgyvNujjrcTEBObv1qsyKK6Jme
cgrM5ZXCQGkFIKVbXysuK8z0mJfhEF1gmDc1VXih77NAq4BXG9z8hlSPhug21FIL
wPaznDHhec3OwYdTU7FVyLSurKuT95cQGjQV0yl5RTfwJXxO0l4AYBtbsfyMrDK6
AcNsPKrtAV9R/S2tUV1sC8zf5oPHeDcBxciekHaX0Ajy3uZ/blYX7Ks+i1eWk60K
QzZztVKhUN/m1OvdqixAO+mxLOZ4xYVyqbFElFrcia7qGiiOnDakOA28xyBG/CPe
Ic4Xkyo1rCH4SzNzDniRiMz561EB0Vk4ThcsZ0OJmA0DP3Renjf1kSnlFCkOLwy/
iEMCvk5WZFzyawqKYS6TSqRWy6kigMwvnhGKrXCCs+do5tasTsdIqlKVo6wza8UT
lfYdyKZN/LWQKjz3Xsn21TJHwjOmist0oOqshB4zottMetv7QnqMSijUUNElCLp7
uq6f799AQprot+rldVVLMhXvTKW/zqO/50QTJHt9L81avHGC8mNZIDaQ9y10irN7
B9z0B/oIMUwqTRum5qLtLBDrByUio+MxKuZfChdXOfYW3S+cO0EsXK3J95Yvgzna
Dx8rbhgNqMTQjpMbFc4K4iafQmeaMGWMOAem0s+3hmbwxKtg16oqhflhl/1njIZH
4/fuI46xsef+nVt+5fBn1CwkPpKgwksysPIn+BQpQZP8L2niZ32lCQYmnV/bPuTs
MN17E7H1xKrk/0zyBJXCYa5gRv7nzlXiFZmO8i5+EXPIFusTcyCb5rNyudlYVLou
km/s4rJVwewJO2T7uo6YUusqfDV1RlzRXrexBDOoBITHzsC1FAA8glCzf1T5uZWo
/Eog893kfoegud9Bl7mTfXGIkW6vb1oTmsjDjkhYtcGHB5DAui099joL5xWErU87
kjV0D8IVdHtp/Y1GhjVnuD+pC9+TuG7LtsM9CKfiTFHvVEPIevZZfOkzVZzrFQF5
wYgWyN1Fd4MGRJoDQZYghtBUpPyxAYtaSl9WPD2vDsJ0Lut9EjEMWem5xS1bjAmc
fFfGdkJd8FqaPvrdcUk9Uj6bi7hqf3cgb6lPWG/2A74nItbfplO+j5Zeco3LnsUm
9/hoYkzMZfkMeufxQfn9fOL2hgXRyzlnnVLS80RQHVLWXQgkg1qxYVrvvxFc5YXz
MfA3QpKZ7E4sZvH46+yTuvKWCdTKwidHcgMmW3/ADYtNzBc1PQzj8P28reqgAtj9
88HyFNwIfmDdaagtDRXSmWo0jjNdsdtkeOd2fT7p+eLYGNOekgJv5Jj9oBMiv7Dn
Mt0QTnTHMpYEiX42HSMz+PZAbBqEzvUiQlexxyxEtxVQTS+T7TBhKpNHAcoHwDRA
dUMTNwC8qt+w2Z1Kicd2MA6leMJeySXI7Uzk7ufwK3lKLD0MeDLT616F7FU9jU3Y
BJxHV4Y0DI8psFEclUbbhMjW2kaHDX66v/FQFaBdGtzQD0h+0ssqxdLcTF4IKMHp
dP8cbY3RU/ZOxrE2Wd4+cJiGi2LplkRisC1yG4cGmJhDqD7vifiBhbaDbNw9Ocnw
fl99RMvuHRJExHJB8raJZibII2PZh9rVT1YIv/PokZY9V3TjfKile/+nRh6kZ9lh
rjFUUSqfpFV/oJU+xadEKB5ZIKcsgB0OzHlScvdoHHJej+P0akoRvHO0dA5jLpK4
6/1L5LOPk0uosTfHjLKYzzpetDqkXNROX3koffQ2Vk6PPgln7PdOVcto06eXaXLX
5bJ/GNauJDIS5Kj9TfJIZzjhovDaOgqdM7xte9AOX04vg1kFIJWNhv2fM79hgAaT
9iAxGX8BgFfcDoF5lEh7LQSixObPxHWHdonKYzOuuS8HKapEvKajDTTYWwZr5DPT
N+VFPhkx6M1UN6w7gibKfEs4EW3DPWJLa8Qf36oGNerwVajv7l9AaOkRtqGZxVjU
t9/ylc2MLrhxruaNRLlJVeXuevbI9p7eFdns4cB3NvFY6hJlw4D/df31aFXTBPFM
vyx6Ct08kxR5zpHON/IjJux6EEaUhgrWoV3rl6xPcq2JBJ5wZ3oC2wfGAjIDsPhX
9V5phbeda9dS4U65otYyQyTPyQ/Yufhld6u58DysulEL2Qr68PjQi1BCBL76olBL
8xeR+0TPHI6kbS+797jxvYeYvw4geTKFW9F2cRLfuyb1ce+GC9V0vmd4+9+5vQzA
Mfm5JkhZYPFWyxIb6TYIAhhRY3Vig3+GQHYpKdGYYWpeVwC5camWH/unlrjdqQab
uuZcFWfZ4XNrfsCtvxbEiylF2ZGJtcGpS+S7ugcwAG8kgvnt+6D4hW8efbavOSRT
OhU2V8Kkcgw2u2WoidDPJLU6IYy2kQwC/HaFbCrBpqahS8mvy9O2JS1frSltnCHw
T81qtDI/ngAkQN6G6NTK6jy7OCYCUtusQzvEkuSuR+DVxF309v7fWPbSAljdfRO3
iR+sp9qBuhSLpyP5XaNsFJ3m+yBNjGU8Rks4J5mkmhl4OKnQJiV4Un/U0vuRCmhi
Gy4UIRNVWrL4+eqv75NAJdEZVsugfvALfUlQUIUrtI18ISuKqHxEwvKSSJTPblD7
lpVR1Nvh4/4J5eiZZ4hT6SJuNQ4698M4ueZrRXIGY20CzXeb1ps6DLODohdgpDmv
oHTtvLu5jm+LyLMpgdio81SwKQOCYF5aX9bY20GtKH+5zTd65k+tIKCphxYhA8Or
jpv16cKMVfXdziAma6FI6m2GhwGA4Ix2aGyM0RWdy3Aob+jvBSJWqruW+q0cEebR
kRKbJUYVRp+HIqYSzVCqGfC0wJzdHnJhP4tT5X0mKmn8W0Ccsef5SrQT+AuayvMS
PRLvf6d/buj4hOOPmnColfJIpdkiLCdURuiG68E5VlF8nIk9PrDBIyKAUjeTikaG
fSpkji7Mv2WzHschMO3GDOIoNTQCyRZ9fk2z8FHv7jfretA18HlvHJ8MXYxnS21t
27oazUB9i29JasflBN29624Z/MFZh8nmLvnZa3sHL83z3tSuahDbMWUHRHvxRNpU
D1eSOhnX60n3ucbkhAMxQWCdfykgS8I6I2hobzg+uA4f92qxf0tOWlFYfsf2+s4y
7wXrr0dR34EdKkoTWOReqScHyn9SJ8Rt3fMFcxcUkKJ3Rz/FLGoNvltUnk216i48
b3Pcmddj+HKPIn5ge6WU2a26dYwW+OSMOdyh4QTU0RC60lVGnDe07XneeTIfp5gi
4rDi7CqE3xfgt8zKvxTsAOMc9CZkFTafd/CA0nQ42fzMa29/vz4EK5ivvEc1TCah
QOqPCi7Zbu4OnLFUIB3u46/airQ1qFK12PV+9/xMHXUzLkcVSme7Kklu+A4ADUds
Kj8YdldHZ2tv+ZtOxBQfJseL7AK+yotAEvpyfRttaH2+Imw8k/JoxoJJvcMuPJwo
hBVmAbrnJHfA+rQujIscKlOfEMh/ExL0oNsVfdDljM2xtTcxXYZ2ToMciyzuKDEa
cgewD6MG0oDcWGyPyHbAhaRKoZ1gGC6LTqdDH8Sg/sa5VfZE++abUyjov17DUKLG
yz8tZj0EvMUglGKZssKb62Jnl8ely53GHO99BVs0oZKAhUpq9zdJYnqaxbEAtf94
SjKujvzX/Uhpbr+nGDM70MB/wBReDbyWkdarGuWUC9VD0CTkVX+aDABysTsGPIoK
VORIp2oI6UZqF7hXsltlHdBHyCHfY6iNWR4X74owcd+4PI+F5kO0mDMMEGfYz0c+
WjGbr1TRS9S8JGRvJZOqzgGjFJzBebMtulv8uzK8w1GXjZ8pEmM6h0FGwJPoqlbP
xVkTx7PvxrhukGUwPVAYF/Ts4m6WWK/izZp2GWBV7BTAS3jLt3nlZErIk3Cf01Eb
aDQ4umreSIV4uTDp1LaeXu3REgSzGLQyRuWM9bbxqoGVgXGWdAxAGq/WACnrAGEU
PkChLinhJQYzlcfHufi5PCiuHzmb/0HGu/SNpJNJGD5+0QVVdKKnoAOyYul+AQCN
wYyyXCNelr0H51I7cC0IJroHTdnTN0kTkrGo+nl8sBveSvTabO5TBACLU5H87Y3A
copKb0h2fzn+sq7CLfdily+gsWtbriNRf8mWezQ3rvWokUODi/DNaS2h4NUzpAkM
CrR6+AEbHdgQl4JD/rxPirxJpmTVI5nl2dZ17DgpLtXgjpDpCNAJG9lch+PyUVSK
5nJQdQCrSwTvHLyJ6/EMuth7GqNW4IZU4GMM1bOqHZseXWrJEF3iOngeG7zLrz8W
LJQ7og/H4LBHEFWnHyG/YK0GhTVjmR4hBO05lfhbsuRZFM8zIXmHYNVh5DyZSD1E
o31+4uQj72Qk8Cs5oQmrqZCoY6vtic3qRSQMt3hRDsbE0YtPIY2uTN02sjnPczOE
u3yO91Mvt1LM19JnAQ5q1ucAhPR3cxzsHEKj/++/uz9VNdoXh6rzTtXjIDR89QIM
/aEpwQc+rlnRp3mwtD4SYPey1BLPEpvOQXfg+0BmkIH4s/kSK8zAFaSpWHyEhPrs
FNKS5jieLf5uBOuP6TxT+SaEogA9iqBJYucimZCcyNB9snFIKwtPHtTEq2rVpiJo
D85gDbT13xkBcasZxw49lVrXshRUHU0VZWWSC1A4A0YYpF/1YFsWGoi88cqz/w9y
zRAnrzIq64mB1tTUg2/ADiQJM28pbthLVWD9+OnBTtI+U6viY2SR/3I/mgOiYEUc
4vfKzfHpYn1XJzc3YYjdsBT6Ai101iHXfcU0HYhK0K9SOnOfkQ2OqOPP3bIspB5N
WyWAHx8Km1PYzxxS+bQrEBszpV1TpCGIpyT2p/3jYagVmokf8mqhf4a22Zk13clJ
j+7dRvBB8PWetVYwjUNYj1SE6rY6v7O1aJASscnssmw/LTkh+PDX8kDfi6Z7vqQT
lRVaX58ue2NtV061iOH5PhpvEJ21icYQ/FfwU6rudYb3BgpXCAXb9/hHu50RVcYf
VRXwyI0e57hADSM04dxemCW4fSi8uT8yciA9tFL6HaN6Hh5l/p1H1cM3xg47IiPM
CaVLi3rAf3HMUvXU367sz82meXxgV+SwhSfp9gJ9RcqZ7qCgjTojYNPYDcP4nk2S
kTOqTq8IuASFXNTQ8UjHPw1tAw5EGW/20F6JuFO6wHJPjhEm+F8HcddWkXH+Mlh2
eDuxmWs+Qn1xJrHECkk1IqXsL2H1kDKniOu2V65oAkNv1ovVLyw/JONJPZteAbMg
ZvvT4AWS4PqD1g6i4gNxCbRMKHbIids3UF7+VmWWU+nDBDG3h8jDTTIdXO8IDCon
vkzRvYhMdqBm/HKbJPQA2AMu1fY9EzYPRIuIn7xBGUbngDpzfnGjPzD0H+2uLiaZ
BApuDNRt7ouWprcNzZUviOQpZPe88C2G3/vqcfjIv0jQNSiUbSXgA0xM/EL8W6ML
y6z8Fxq31dwpfDx7QraDp+MCf0mVuo87khy+5bQRQBL/FtLXrylcoyWSCHEUsRSA
1H694JLaw2yh0MRwI94TC/poDaV4lDuh7bwstLZvAbJtvREiNJYlIks6K+525Jm9
EWAg8ES1w/mG8GcQzWrXHVmTFlKTz/0+X74OFBO5pua7xLt9AbokNqSx0DIDHf8U
kYbdVVflyif81bBp7bmftayFXJrPq1GuP3E3ex/ts8TwiUvFH7CTRSOT8/y4Nc4w
2y55cykm0tlnqzR8U8db1DkzUHV5HIZWIUPZjpZv8IqDt5mAQYww5yU5MUsCHsj/
NRUsQpSN3VLkgA8lVd9abhEfUFM9OtYDMyDV8lYKgiwxZJcZmMPrI2PVZy8bzfTS
7uAQiuK3YXYgLQW9kDnitUfad2maEG/U6PBg3pfhVDQF5Qq/+pANOzLkNeQC7XcA
4FyzD5BNtCSwW2xA1CK5arruqcOVXzQeGODssSyyMVLHoDWm97DsOaLfrVG+cvdK
nPk+D8uxnDcKwrwt4Na2nyiIcFJyHziFG7quDidAqsZyMaev4qXncUT8FUqKjEnO
k8BfsNwASVzRzhpwvk2zlyvME6tBJsgjsuGXHHaijI7e/o0vuw8j48KxVRt5ZJLa
yIHEyx0Jk7UCXPWCJR1v7cykRUUEdAS8W4u1lrS4i6lOcZJ70s7SZLdM+Tifi/CU
yHxaBBMaDJHCCYNqZRtBx2NLgKFGUtJ+UFhbZPddavSQ7zVt7oVrp4wOPZZuopYj
++C8WQT+OPfGwXch1U/4RVblZZvadgflatn9S7xN+V2iLt+mo10YNi3mal8SzPJM
bT6FmK6k9+NYDFEdr+FBLNiAfEifEI/9VZb7CAxUyc1nRYBn/Y0W7xqdDulWA30L
MTIhTGYawvODNopdyYEjA+jocZiHcWJ7HBCLPpFnirTS4HEoli0xAEwv6gbMZV/W
0svEr8zSEubBWAd7i0VFGAxF9jx8rXovwSTsXSO0HdFx7jv1yyUHZ5aTFgA5gaEG
CVivXdT2Cym3D3G/fhxJwiG3SpXTyxvJHz0oemzO8R8zocM0m1uIjZfV3MOPT/T8
gTjBDLwGt5frqt6TS2beL6UZPkYxslWMZYbJN9edi2Z/fZPA0MF8UrNew9R5bvFA
0hjyyX6WgT5l3+mvbxFQkUc7EXSLFFiG7A4kq06EDvtacTnBYav/MISTlSUICVux
FN7Qtn58ibpsTFoS8OaReuR8/kVi6x2GdzbDcjDrCAQFjhUC7K6ocqK7a27RTHzz
+L1huD3jlHgsooAJV0pb/Sn864sC5nsWMQAc8AWRgBH8puDM7PnY2xJVFndagA8k
wN0P0PEf+zliOjppwiq96/XFrDQrb1RVRZ83bNsCQ3AoLFuofJ21PfiDP+men+vy
4l/BmPF8thDe7YMcfeQW1QdVGRpdZjo/jCd1CI4IV6Xr35WW/sC5xadVg0Lar4G9
QmR7m8dKSjr016UrlO7R4T8YkCrnGImgogYT3on6ihVCQhTP4PHtNMfRsPexhIBp
SxEqJMAVvPch8wmG/BSTZnktHQHH+q2wE1dl6ius3VfCATLssqs5PcC+LCi3duDl
EbEHwuYDEoj8NOuuoVctQ2ISLz322t+7qOumWPH7F0JDz83Vz1Bgi/QS0STt+0YO
Yiq4RW55ySjAFbgTgz+JXnjVxwiJoLWMSv2rwFS8M6IP4lmVqDp9WrOMDBDMHQDv
NAA6EokGDIzwbLLo4ADKI7WUTuQCwNF9vFtIG4e81XCI6BSyWy4SK8tWJqsKY+QN
039dtHG/m9wiIfuNl7L2gLVdiKftRiHSjVueYC9zwGaYmmcj44MGTmCGKu/F18Ky
wQKP3ERym7UzxeYXP4B4kcltnUZ2tqkbTiKyHXsGKWFU+F1eP6lW1tstF0abRGBF
dNbUIUP4kJRHeSh1HnGJyQVEFTvdbr0SfQsDFRJ0VQ9X9Ae5t3bYoZgnlNNJwk5h
ZmSD9Wv+0Y4uplh5H18Chm3Bakr9iya9ogsr/OW5JHQjSLVP1PeeEyWa23C0ubTB
LbspdhXDdR6xgL984OiTwac5nGBI5IB869W4gsxcFNa3uRdRyl/OU6CCJ3XNVYXB
M9guVeQZMw6hmSwEtEufGFalY5GTN7Im9CU9J5NnzuGHcd/LW83Vx6N7/rtgIgoa
Lis4YPh7BWXDqa9+r1+Uw0pEepds56e9DxHKfuYQ+4Z4hfvxnjIZPd5yteqf8x4e
1yLO5xM1MilRJNTQ3PNJW8A3r/dQ785rMglL5E5kEZkqHOyaU1Df/Fu01awYVYkv
MFntyubZLRBRfI3JEsdRMQWUp6KgFS8hDFL4WweIKxRn5toumuCM18VKuq2D0ty6
Jc3z9O4QkpiPrN0wclvgmEZNvFYodyBxFbIHp6a9PA1/dMp1zstq91s57fSgJCnU
CuONgWPPhn5wsBNSpTEB3MHRjxpEYJFkHe0JXVRfRWpXp5h+flRrQO9sfKlqd+Qu
mS9Sn3G9cr9+MmuB3Db8FIEyvRajPBr1ZXnTD7Tz81G3+kCSqxQqGSfyd8tmwGoe
ygKSEwrXESu1eqUpqzsZRdz2wQsDRZO04I/aGUMHYGWIQGwMIXXOSj6HURpmNavO
v1dRKgodeS7cPqAGb0LCGls+vB09hQm7akNhxCnUvPdOTnMwyAlef+aG8VUFSiTe
qYMuoYAnimDcna42nc0GOwwOVS2keNkRJF7Lha7q+M3NoTBXVVNZdl2YzWSCq0Q7
esvDS4kDXybnjGDcDH3lCccq6s8HmkVemk0OzfavNli8WMpPlhHST4xTd4N/sM4N
bSebhPX36oRCCH4M7+W8aO8oRePj1C+xiU+MkdC820VrTYGHN05Xc5/e1j9v10Pc
xOpKWyLztecdJ10Gz/k9UKyambEYHu4HYxdbDEXVFYfTwkoLiDdXWScAfP7rmkvv
zl5yqzGRO6j44NFFJfQ8NqIESxnS6HXLNx+JelIzzkoeopiEM7BeI0dA1scCJDWH
5E3Hb9R/w0XhL8L3YdVI/AXFFUUQt3atNv2ItIcTjftRzbJHHAHWN3THkTlGogUo
U4894OjdjIbQxNt1/6R7D8MgRDlHSQjSuGr27vWgS+W3GVoEky/iV+aEmPR/yhIe
KQrTF4NDE4/2xlAnHpQSFKdVzy2Arsqzc6xFnR7Wmbc3Y4lSHAeF2HowvEA97pSv
yldXyXcjfLjL+tx6jHeLsyXlLcZcsjaObOGspePRjOgyd6p7H5O2dXmcZtBNVa6I
RpXqDqs3amR21f4BlcUpKPasZ/uXQOOqE0ZtWhYpXajYCyL+QTugqBV9m2QkZLdf
Otwaat8yDYIZ3W7x8UJ3l/k5JRSq/4+XqEm1LYDCdmaFmVeS6eXJoXx6SeHPf6JU
Aojm0xJoRRGj+CXZkynGRVcrLxHPzCjroU/70VXW4bsARbO1K/bkQlcAodB22TaM
Rce8mh8Kmfhy7kwn9ADIDn7buxv6RyJpdP/Jb4jiVNO6ouh5OzuOBNe20H+mYZ7c
PqPIPOFy10kTc2HToJVIb0bPTJ8kDTy6Fl2Be1ShBpTopsg80BEoV2ih7ULdIsnz
TgJxV0rnot8iR4INEW6woj8Pan50U56Q9MBQmbjIAa94y/ayMwdMjmwQPnswY+rU
/lPtELJ1TeaQjWLv4A3LGF63Z0Pqqv9eT6lE769futityU/l4Bbb1W3WZ+0A2lVW
18Xw0lXoys7burkBQw+PbnCFA7Lx6fwsXSel+cscTwL3o0iL/uFqTRWwzyzQJkjf
waiwefWBuILQp5rqRgJJHBZXpXf2dFMlLVW5xQy+KhIYG/7RZgnpkhCiSPEz07P2
myzv+lIix+MZ4zQ3G7d9Y616r3ik5YkWMFdT+F1skHvN3FiPHsoorrat3jVirxJz
1jk6dg3sCb3+Nkl6E5RwoBggB+wRhDi0Cwyy3nB09vnGc5QBMYSE1OnIY14dUk9f
yxAB4Xd3T/CQKsEKNMyY7NH1zNvi3ZwOE4FQ8tWrzs4GeIEe45XnwqIIx3gR81gz
EvaE1U16W4uIBmjX/J3niINT8jw4XFYDhe5KmnqqspISm8qS57P/5BV/3mYgp+7m
PZclB1LmDQnZFxwtMtZ43mw+ikprI0iQ9z9netizZdBId5ZhaR+/m+6euvH53MH2
Mj0kXBlXprhq4YP6M5mDbuAiTO873C9rzRDW6SgeP+/EqhVNDO8n/jA0JLbtq8fi
CxnwNZ40kCDBHx1m83RY7zC2g/9ezzFCTqi+zjpwYQ1344Q0ho0zSDn2E87iIos2
da2zRmtA1pgusVmwEwhujaT/SngOktmjupm5GdCwZ1afXiRstC9dTme0XaraUStC
K1ZPqx2tQBa8oqDBz8ku6U6kW7xjumJqxfSd6SnQige+1p3dm/ZmTW8kp4PGTRyX
drbwIPBQLyOHfyVwherG31M3xq2rvS73urcBm4scqGoAIPdxQyRasqKF2DltQnfb
f3gegfUuqacRI35o4jNdNVorXXwHdUSZTjOAthRpolIkmbq5hzQDBgO3aJMiGVQ8
2mc5QXO8r3yKk54LkkBPVNvzmIuNYZOGt8Iey15uFkBNhl340Ms0aycHUiXu7XGF
VcHpRlXpHPxnVUq7CS7L/VrIUVkAwuetNR4+VxSlelK5oCLVNcnYIIjbcilktqFN
pmm8bCsFcQFO+2fWWxpv3vDDUChPMsrenlgvVuOMpAv4z+a/pgiQcAfD9Rzmqkv+
V94mivJbhPNikQoAk6A8uD+XfXf9oXeZTa7aHmO3LznrSyTfnl/INYcJlh762SKw
FKTMAegBVOg/FKW9Gtiaviw/MkC+Up1E/fr1CJ79lNkeFSASq4StL8B8xQycw2hB
O4Xw1t8Hy6jBbGEBNLA6kMVcWkV5ADxP3QjHuV5Tf683kV7CrSEu3H1Yzs6C/Wg5
RWyoQbrtm5t6oLLAFbBvtmxgRNlHie0AbiRkNO9+fmqiHQ+VYdl3G3jJUP0aWqNy
fKoY8afCYRakE7F9eYm86CDQFtcLR3BitgxHAmZ65cJTW9rIC64fiHydHwO3SsPN
9/ePmcmPnkmjIyapcmKBR1632H1QkUlWB4ox+NE00TnegQs6ICgijLTS7CP2jBt5
A6DuD3lYisKEi8bHiAK/tHmDF8lpxMvcsaQqQPTxkcHZpcK9sg2dyJl37+ZvrsTp
i28/mWFzTuGWd0Gaj2TNYQlLj/CKF73zHjJOFqfUTwaFxNYcW5vaWfPeAjBJUK89
Oh+0oJCyyzwSn7LhgWWjiEuat4kX5wjhbdUEoVf4JkFLTHbpOZC0ZEl6Oh6sf/co
N4cLoBK5lz8DhSJcGWy7oFprxhYRM0q0ZeFF83DQeeqKdbkNhjz6Phq6YqbIP2Xy
vQ34DLxbcy+V7rvem2kQV5Unt5Vmgnqo4Va0rBYViOy3cKr5/32RTfWVKem45XgM
Zajm2k86uthw1P3XJqRqlmXzR4mOSnaOKeAU53gc4XpofPXi11ic8hjPZQnM/0Bb
7nD0Ydcsh4jBQdyPnv73o5ih1AkEXzpv2xcBjUiUDcIxiAFpS359/f2+IkZoT1pi
kgcARa5qksuNvDso5LgdlQAzaVbJowDPoeIGTVVQ4K3+rmpUb2Zm7GZeO5ffh7oI
++OyBKRSOMu6wBvYtGFjIDTIAWVh0gWen0a3OQjPpGpbmgmSN/x+Rt9QUAJ8Qa7T
WFLc4OShn8KPm7aIsOlvj+qxOot3gfVQL/wPy3f+JGnxtwQ4PHJxAoIapyLD8Elg
SRGA3+InXVkrMmrrPkkaS1lxBx4QOqKkRnxX815E7mGqN5TembpAr2ENxdMNeAeH
1xAfmCMI0SkPVsP+yZr2isLYa00qxw/mNKLhYZrWoB+6NgN+UK8q1GfMcw5QK03V
caQxSYnrnzjnXjduJY4P916jvL2bfruTZyFR3xhpmPpoF7sv31ASWujCDdxT9alk
9gmselJyb5nA5bN6Psit0ORE1Qlzj0YbV8u8++i2ibXhKDI/i6JoO/OdVJWyKeuO
+si7Bwj7/y57xDHOVyIUhIZ03T1V/cx9/SrYAUaksL7ANQdtYgWqCtftRyDqamMC
OkVbx5dWA61wZVDh4Brl00SpXriq41cR3NndDDsFpOdhR7QnHSVCyqGuK3zor3RO
x7BpiuFm6I90n4Qz/uUpjrDQC3EJb3o7yZqQo80ui7d2tWdxTdHuz2hSZyf4FQ+A
r2w5DD7Jl7fmIwu2f72tyl7ue25XXlzZl3wXKgh63qgmYvfxkHXvL/TnHgdhMOnh
1awwp7sPUuRlLM+0vMTqo3vcKZpaY4JkU7QAQm2ut+WiSNcK/ZNOWw2PnbSPDKpq
wkplr90BsW3t66KOMHbhDc6Vat5k4PW3yL2jytx5qy9sueKSrVe4l2nOED44sZri
SzGMGcl49QgdhKzADEu0mu6fbJoqIh7wCDyJwqu0cNN1vUc5xarW8RN48JiRd6oO
aH6dfXGR/D1wXeMOcdMYA65jg0sm1OXuelMLNZNtIS6uvPuRP2dMzdE0HUwzBpgo
zvN0mytXKLfcCK/B6mYjneUwIa0kBz6axchKQsKllL+iGMba6nw8iRHWyC3weq2H
O9pPe1HUBjKafm+fPv1lvzW2FhE0eHy0KwYuKiD7QjtVR7s2SepYTiZUt5qpMWc/
4xRZzhSCrxvJ2NV218c5WKXxzVmhUtGrJv95aoODIKng7rWtz9s2hpZohLbItKyb
J2+s10izX7SUTMBIJHSQd6yTuuZhtXNnrL5Tn1yu/Vu7GA47hSs4az5cCvQcsoAM
2NDGF5defoG3wL100UCdWDowvR/Fm0QUwoxjH4hjgfbwFSohoXZmjiMpCofNl6Wc
wiALyXYnnPHQgT2lMyl+G8h/BTIUiwRAHRbZYqIkQ5JWEOMdDbYBxh9WSdmqg1VD
lQlZzEoUEQGksQqwKnhDfRJTVVBKanESbCVWB+Hueb8/j+bvQt5siNmXAq4xNQpl
R++3uApXhpGnEQotaKfPXjql4TgGxfaz+crHsXQw4hShpowlc1H1kfySQ3/yFx1y
ezTak99jhRbrhJ11v6JzzeXrjPla/o07bKxCZwW5LLq4Q6jbAxipGNtXSI8K+8hg
MLK36tLUYd0iS0idXdR/R0HQUMU2djDj3oNtrmJSXZ0D71kOFx7gXAbikrkL+JM6
+KLWGMJwWBHEFu44hVfpQEaXLNOCnDcLjFi8h6S3bPCnBIeaTmyNcwezn9kuBL75
1x0JAS5yq2J2waK3QAO1yiyel2VfqtNvIYtTgR5OLIhtdfCyIE3qCyiBv2qNX9On
Vy5KGzjuzwuadXLgnRPh4XxyFlAEO2JRSj0HA7qxGDPhrkB6hyPV61mpiSoXXaxg
EmhO1gG75dg7gUenpqGA9NxqMnOyijJatCNJBuC7upCymLNyXtH+IGRXRMIF9j1f
9NTRfpIVMhEsaKRUN7GROrIOgT7mlgfiI4XXH+abCRcF/xLX/xC/AUUpiYuXWy5H
qGvFEeAjb1U3ts8YgukEfY7MwqdwYzCjpzYwz/GHtVjp+/oUcUvHtuFAta+HVBB2
HHNYjGODe+lMbdDiGMzfcBj8lzRmhIoocsvEu7xzcw+bXUh/sDciYmt3+AZ9q7Pw
SCCO9y6/5ryWiPeq6d37vcPCW6CiN2RFsDQzx4i8/nr0cACyAb7oS2aSaxIpGsXw
5jGP/7clTBqeV4CU9u+5j30KlQMSnIfEG5DEujjueOQ5o9ZvvGPNeR81oyFf5Ras
aHNYt1z3euy5MjYm3KDnc62ht5a8cRxhvKKEBLQU4mIpizzXQav0YAaUf5ctSlU6
O/UZtwYUuk+7wWyS2ukwATnl7n2LTPF1vTtupP2iCeAwVSOJ01UWKgHCzuPY0xaB
/lAo9RANuQeibY1kgo3lapxoUBhMuh/eH0AofMiAnqPXw07MM8v1E66goJjl0vjr
LeAGwUAFBbRoJLLFIGI0Qx6IFIkfMeTdZHt4mYcdzsa6GtDdsoxmhmNEzO+qob/A
ToIEGCaypzuWhinrBTcvj3A4Gyqm1w16lLR4tZKuTdnXLJCNcgokuKgyv/Cuyw+X
nf5sGWGRXk67aTBf6uEeHLX2K/e1aIvU8hagx3EL8lqA6qpIHJFn+wHzjEcOR3kL
y4faRTba/qtUxQpEQRAWNKpsvyJGeEaBrarqDTZOZldU/Ya6um6tnAy4aFYXFFRH
arxL8iOXt+JQEV5V5RhzDjVvZuzyKl+6nqh/OOi0SZvCWQbcUC4I9tsMCi4Hlzb0
q/z9QjPVp+3FjjNd+9sS7H8+PTWkNO9dBNaxBeX6gvWyDJcLIKtNB8jSSNJ2Il8p
vo6QVrbe0dF4JOw+Y813uoE9T08EzfFSyOgxgGIcBazTd+bIiAtDGEBpsto9VRKK
4M3vhKXuAYkTrxBJHdPRABcpuB96SC4smsvCGq0Nzv7jIRNj17HaIEOBjLUeRUy9
TZ6kNI/g+dSs8+7NM7T+ZQN801dYdydcxtifntUJ4XpYiUmnIrAEYPL/KXjOAgZ2
ncCV0YI2dTfIaIb3nhn0+wiPBwYauviAXA4/QBAUqgV84QfOIomX9/vh8HQoc774
Ixxa9Y00VtSLQMBBRpxPNxbvek/8h+CEBizXpYhn40IFTW/5rvuXNoCfqrsqMVsh
wCvg+z1g1mULKA7lH3++7Bpg+we9B3Oqj3J+imACsVOk+fSrY1+bzicH7spEdEgh
u+jV48XBpj81mbvHBsIgvW8DHZfTha5cpe/+rE9FMl8PHPXZxnH5YHoBLxF6uYT1
NBWQFiRsLTdjptGKLMX786S9ibg5gPdEAGlVaTs41TIbG8bQRz5cV9kPX6Xm7ISt
KOh94V6GTLUD/cFCC+AoCrN+aoxAQ1G+hIPWGEwoJtJmFSgIFOQEoCOOg4tVo+A9
hgyXa9G89RVjOnjLo1WpgnMjVPXKBNgK+WYdNbkyCtGTU+DQ/Q2FX9tv8WwuIilB
3/TXw0+XcDYBUgr7T8jMleuhvsCv/6P7ksfOSoZqXGrXJIk0G8cAqlCBZ4AkqbeE
IeZxfQtoq2j8PWdfPstYcx/Wvnf8E2Ne0GhJ4Bv/PUdCvDCOFwFKVrv2HqdIFFFp
CJu74jcTV9TGU6di56ui43bu8aSaIl4jXi3T8wYDCpkSh46IGxXui6qLBJ76iehM
5wRSCy5JUX2teAgD62uyvzFqkFqIElKzDnpJkrtWHPAGVTp2jNQbFPBWZo2gxRdl
8wzgPJhG9wYpBtdQny9OU6BNXrGVnvJLnaqz0cKOx2oghMfNc0XpJHS1KdP3mbz/
1eUUqYYjTDea1xV88LD+QbgKNvcx4mt9EntO436t3tDODlwMZ2LWNffEgTKTpMZO
bSQkVTnexbn3vCaby5j9jcGIbCuJAACygeZqAetrCGGPwSeckQzw9uxGpayvGgu/
e3UKu5rICkVgKI5LR2v3EspspDOc9gouhzC7YfnPzaFfGbm5Mp0uwwAMrKZi/OG8
714NkjMtlO97OxorfPAn/M1VivGd4M2pkCF/WEVTDsTvLpfvFw+2krbOnL+Wb3/o
Xgpxhy3rN8ikMHljCznnZy8wQVXg43r32Mebh9tddM6kSGo/KJf8Darp3pym+w/J
S4a4/KAGmtryRcZrVep/YwBeJszohAqMYm9nyifOP2+SlsQl7I6fsiHvJ/I/aa4x
LuNFqolISDqCJ3zdveMLdcrHB1epRGm4klXmOKxDr/VJ9UPw8kDe8Cusbyhgf7o3
PLksunbdLY+/hPA4mZGAvUSxkeqH6boMnAQL7Nhe7izLteLLeFfU4w1GQiTdiMC5
LCBDCxs9Z9cLj4V5Sc0JdqhoJLDzWXXsFk/8Slb5z8iOxvIXHs4WhZLb0i/2kicC
fsqly5nJtP4E+UZBBxvEY70REHQFcxlBd619KHg+01kWkpJ18XVgzwecssBIAzK6
vYvCFkQ+v3bq9GQbVZ1Qd96vvw/TAOOImIsIwGss5qTziW9eYFvZWODB1hgI2/b6
RnmlBq/27ms0IORr1NLUuLbvsseXKqXQMHGrxvjQ6DPbEtQRzj4QLhLHNY3aTqqr
j3gfGt+kjDL1N5b+o+UoMCxisYHCijp5K0VRIbVVgMjKfnon5E9eM9bhUW7hdVG+
Lbd+5V3HUSxbMKnJb75vP7tOVy0Pp3sTkX1Tm+BJM7ZXJZCV9iL+VAzMp9ubJR6M
9WQsHSl2vGg1ks+nX5yhF/ylcEMdhI1UO4nROPAGTxkqWh7TEcyCP7IshXyc20Xx
n8zT+WDdG1r2y8iMROcvQETzlCeWrsMsrMqcZ27vXqQ1Dkwl+6wTd/McE4rl8HA3
9wCbeuKgK69WfEdtVSbgYDZ99I3ztrs4Dyu1JT6SjeXnlLl5hencBxDH2HSlvBsp
K4kG1awgoNggyJVflyYWod0jkLJNSPD6N+dkzCuGO/M7wadnYAdV6qQIJj//3B3E
5amXkxd2X727zE5lT5y6vZ4KCypbqYGJVPfjy/iVp8tTe2MReKUYszt4s1FNqFml
WXeZ2mKItpbs5Z4BTYkBhtDs2z2iFEkka3tLNZkf+sSTeFzzY+9aRyrjBGDpwa/L
vlw5GwORmRkWzC82BfI/3QL9n33lfhe1CEghrwgCt9BBvWkytj+1F02wamBfQwzX
KJzWxALWdH1l3d3hfDbq5CnZC26zSLL99B4t+aj/IIONv7cP6jIYr6GvzRs3Jdml
DAcK1ooFfNFz034qcB9gFcIuoFoAlQi/pasW2pcEJdzW3LLIJHTXDsIcC58nf04P
rgtxkgiFWbNMidGbuRHaU7qu7hlwr7sukPanRoi1kFRXHD0sowA73qXCeAbObYEG
zShtnxyBLEaPT5fCiv2x80z71HjymW+F8jFQAq3jEASCLObVMLBQFSD2m+4nTS4s
ndTL/7TSo53EQbJPCjx8IkqZvpwILGrQFb+N3phJZLDbYQYp45g21p6xR7zlgEn2
KdDpKEoLQ2GDD5MEKG/j6wqbJM1o5lU5ng6rfBx6fjiQXo0YnCGlxSJaYwg5v3G3
IoukkFrx5OtShAdG88YFy1HV1RsDpFnPrugZZCZRCluuatOxgAfmmAb5WE8QGojF
p5BO6nbZrwW+EFXTlCxN6WajMJUW1AfEiuCP2FEufulB/WfQMDLwr5jbrcEclrvB
AKwRaeTVEQ/nlARKexQKMnhD8JZ2CEpgylqaPp2HqhBB3zsliCbTUA+/veqycjJj
i1g3dJ8e8Up3ktFBDlcoYILfXUv53PoLnesgBYiomQBGpGG48smU4/yBFTS07+1J
2IlBcywM8BsJOOLKMf5sF5k4maQeB5nljxFeQZyMH8tLdZHfgCxWTj1pX/tXW+mI
3wVW+X3ZXpdWPtn0nHIHWASl/NdzECt6Lll8GFYVo9YRMCgWVElciTn4dQDWmqWx
nQ2BZMzuewak16fXhcvti123imq6KvyNUim8rR4GAdNXs4p+Y/ms6n+X3T7PIQaH
gzrjyc/rfFjzWbILhK7XkliMoqlz2h9sZVBZt8gw8QRsnzbe4wlaw5AqunygKe2V
mSMUsEQBIdFS6gHAyU910bjtLKEeBAL3NnpYJzuFEO7JWcZmeN9e0FBnZ0CWk1Cs
VV3FspR2gYxQ/53ZdJTq/3lMtg7Kkxl3lqw5yzNNQLyqwzQ647uptj4ZVBdzKCXN
7gWNct3OTWxE4tjoaN965dRBg69S3HAq6rBq3Azhd/K18zX8DeETe/NH2SGde+ao
TGuTFOMjQ5o/x2Qj7qBi12l2DUdFD5MURXEWQfDlYDdkej2Xb3kx8NnbHlLN9JEv
x1zVg/HSgNi3LEPg32vyR8u2L70XYu4LcPQCrC9n27I0ayfNKqybjkLZ11id1QsC
GlJQb2NvchA02RmweSSvOxWnARQftZRTANXiSEO2FcK7+qBEdeEj9QqHGuSwBMY3
nFwYATw6ZwgNUI6AKQFKny+3qU25ZCjFis2684JdmIoFyCZUekAILLcUCnpPdc2l
cU91/ObPZmGN6c75RKxz4x6l3OjUGmMO0K35AizN3kGbLrhvRWDYIIaIq56qQJhL
3g6D9sXJqDGW8wQJlBFM6uujPxvi1n0qKtHp+c6pT1NkE3pdJKY379VdtDRwvIgs
uOoKGZtTAhsWFXVOLRVd12Y5DFsszp/MGVuuZpFagkYr0lBiMeGpksAmuX2EAqOk
YXcIAgWYYJvOX57Dkjot2u3WWoqGhxjzHO2Fn5P01fu4SbQDupXnDT54ShRKHB8L
T/noMLxycu7wAiTqJRSxHe82r/ziyMTqa1AFm72ZoO4iqnXu2j/NYEeZNc+Uk5gQ
11PK135xgtBOblHmHeqNh0/kq5tqKTduQbkYioWAqyu3KKeVbg3ge7Cq9VTL31N5
uGQvP4v+9O8Gwo0zz5DN5a+eqJVbswiyXmu/hc6VsKE7lnIqnGYfRmQR9vTLFM/X
yoL1zsWSQ6iXM9z2+v3mmdCpMSr+TAQ9Nanhs9mzYos1cYCWpp5G0ghBQRSBSR7Z
1hMPGekcPEDJP7oC+Vou5TrON8wMZ2Yl3OQ0OXek+cedkhEXZC3vUWefagJiNq9Z
h2YyhBZGJBgyhkmycOYQG6TmbfuK/JZspozO5qUFWPmvVFkm/v0ot2ECFQKOVwmf
llTJsG8GmQpDVCUePr5mS1k8IIP8YkAPwO4NfO13KLX4LvBfKcyHhpIU8lJuLYcC
f8XDtRybxvwLVkAdUqW6j5o5ETAAxT15qxnfZqnKJjDD+c9KLG86uG/o+QR2jor6
Fx9JqU6jPGV6+Tz7q9X+UOjrsI+wAgv/aYcDSAUGyXw1+QbDcjX6ZMZN6khew0IW
+ne7daE9AFoctBV40cxDeFNqJ0Vr3IVx8USxThMKkEdLJXtTOSfoeQQMfOtz+rD9
jQI+LOqY0LrWdE6HLiG/PDuw3BKTn/JqYLRqlHndkTVPV6d5HzQmAZfgrhNHUNeZ
tc1rVtBhua6CoFufs9gISFUcjCy0Nb7KdH+dwygZvv5S/iyJGrKsWZkG8fx7/aqw
GuvVqWEzJRqXHjWeXFT533EoeafkWxgDa0k46Snt4K8WZZEtmG0rsOscAGu+Fper
DjJqhp2QCK2aEULkdZmBvBt6NP5fCT6KKFkMMf4vp8OU7MF9/5JuMiH4dYjOUPqS
Vs/3UQtEd0nQ3KqhAhlPhwF98VIzP3elJifQ8Irt0+4pYc4lP4of0hGN3MNFGSYK
q6abJrgvInqi1OwX5boxb1OUiQV3ybH//wQ89c3hZhzpCBemgaxHif377sl1MKuz
e5+6m46pJkkE70jC6lW8cNNYaW6Oxt7OuZ7GcvtgrPyJ2VN8lhguKF72KcIMd1Cx
ueso2T1pnDcIwTmdltPqjR1c3YfZG/oZ4LLFFrbPUv/aE2lIAAVgPzG+joa8RSub
2LL+PFNteHsimjlMJYOtUMFrgetsXCMxYQEJEyF682zksWGqhQggZjuhajcc6hHD
8JOSOi+8TXzurfXKhHSki7SMZWrDL7ondVW+rDFlMtEN1iFar/Q52xD3voupHbpd
Ywk5ZoiDTG+baJsOy9vzCfROoHRTFJPT+Y1unNVuJMFHjowQRSuLfx7OLquVTdfI
m/7ZMKskKe7ZjrYQj7E/szRLHWHeH6Z7EQPEOg+Uyhhj/XwG4zCr6ySRCWuqSFfm
+wqtnQD29bA+s3QryVrSFgOiqhFdhI96JuZvvcKltZs9uZmyPBsTsxeyrxwz3qrx
naONABBDJ+g8nF5z8w1mnNdaZfl2li7eWr69uQJrE9Wf2m8kGMGfXcewpRshCSpF
O/ggoNGKz/w2/EiE7xtwgDrvq91hJhm4G7W47rcStLznaV9o/qfpsCs0/66qPlQJ
08rpTpXCYJQGgi57u/nPMUBChrVzoUchSF/OjJQxJgc4gZYf4Q/2fMuheYR7HJ1H
m5Rwv6+eWy8ZrWyNBduW2MqSOvDCwV884l6k3eBCasY39l/mxTdhYY/x8JZ9cmJ6
t6Ou0R3NHO+RLu6Hj+HzOLk3Z92QyGXnLdRHmGHU9Jv3OOfmx+37TQkXQffiXUbi
I6poMZwtDEMVpg47LPStQ6BM/3Kf8hZCrik3Q+mGHM9xyPMp35KAY71vc3tw3eHG
vONDZCDJb6dTZfaowGSJKYBjsNjF7HySthKyKlm/X+O31UnKNcdAOHCwr9Wj+ZAx
h7EBjzT3lNjUaIcHS6C5Q+NYrT8YHHBOSN71/Swutw0R5IZlZpVZWbwReo6Ev4b+
eix4Q2JqrqIB+ECrGZJKc1vTAScxgmholrXisF/7mkccOh6abiTAoan5VxPbq6To
Cx6PuYfz+R7C2VRJomXJJE7NatnaB4skBIROEvqmtCqbrzcsbqpt5irsX9T6BZWr
BLwnw6o6IKUD8tc+3ewgH2UuRjfNCu9lMDRmfrmTyYmL32su9lRG/s5KR8Rb/C6F
fUPiA4Lr6agKYhdLJiBHonKZGhPCmieCG/5e2JNkN8nKtEurPNjO059IXXE2adr5
ZsMO4a4I8fDNTWlm/wlIOo08hoQxMRg8+b1WaF9WkoqYRi7YYQPvRHv1BIDxCNy6
iN+6caVsazLU5quCb137ilUi5meaJOAEgfp9xpK/zZ4+ziEo1yWEWmKYkeQqo01j
HWD4g40aIBgPfSDjm6XudwmjOGi5jJ/3lhfLjyDgkzWBnqsCuRpPqDoJGHzlSHYB
TRSNi171MqmlEHj6aN/3OD+nmOxPBcjuzaZODsT6vMepRTSpW5N1jt3FtSF8OvT3
XnTFLWSu6dBgLSWTEWhgtdoNsGUkbndBlCFhJVlmWPxEaoH2wmJVvLI1zFOjKkmU
kpdVC89ZNZ8C98U88+1oHAkXz0VlWuJTbkPWOLKYRqSHqEQdZqwt2qOIWm9dGYYc
vSdWwWQK9w/5YP5SHxjhVfsYWwW0xvJgvnpaCdHCrzQP9Ez1lR6TXoVI0lAFhX9X
dgzd6ai2afwNQosBs9yatr2SjXGGzOIVHsoZWqJMYyYqV4NDSSKelO2T1JSDXJF4
i5gizMTcn217JqTj4tnGIz3s6a6FTfJp7OLT04iz09fNZWMdApxE+KeV+BwC7CEE
vtQgCNkfkW167dTi0xVVgeSMQ4BdvNc1FneRt4FbWSi+z0mfc2BIx0Ju0i54D6av
IRTEvfWBBoMeDNeBXipnmmmQ4n4s/1Ze/w71RCRyZI9XqIssS/2g4YbfAnCUcrzc
iD/tSmb5bs2XVM7khPNC5fviwWxGQfw19ybKAYxJO7XGJJx1qGi96EqFptjr0iSU
Bu0C5YEBugT8KLolgIyL9zHE1diVpyn+RLFDSYueCqHub2lbneSjPjicdvkjCo6V
t2XmtqiSWMMknKVGINAIR1kYnOZ67ZFEfF/50hATVcqPcG6jxBCrI+rvZu0q3OWU
FZKFW0dtjsBKH9Xp5Lp+xk/OCdY0QH+j4z6Q8mvMcfgHfZojYQHf7scp3itxSKHk
PVHb2y2iGQW7On+QaRbttumJZu1hBaRAFwBaAkupFppoMOR4qBRuTbVksjSH6b+7
FhDbxVQVRsouH5ScSj1CNZdvf2UeuQ9iXxFUhWM0jh6hW3hnM1xydyVqhOy7UaGJ
LnTbncvxXcw838aRfC8l693wkx4LnXjEOEY2ui0tatjPP4ZYC0aPdPFxZeV3Rt9B
UV+QHREnvqjSt1lW0humOG9daR3DVtjP6guYarHFA5YooyhjtdLG2zpiFQFJ0iRM
0TtDsqyb4ELArBW/VdRQqKAxkEbyVVD9Az3D0wSFh1hpB0ZNlmewl7cBWxRU7H40
wV4yN95OKShRtJmEN+4tWdWRnl4MO+CCQQzejKSP1je1GGEHSdz+xwA8FkuNWwos
O9uZGqVXL6qAak7igPR1RKOajfHPUqzFF+pNDHYCYZAnVSro/M7fJPQh0PU1fdTd
T9BUO3en9YYToZsPndr8bCxr9KJsSlNFrcv7Z9ZtI7KUqWGiA2XGiByQHW4OvsJ0
6RAdXbVeQQsnX/45FRPpGF+SSHh6g8AApRsPJjKlcQVCXgjQFle9SmZIVALRoIwi
+D79nxYU3zS4BUq5KBNUtGkAGhVIICC5hTfGDmKBXVHOGt4bndUqusVLQNF6wRBc
eVw5n8F+BTl6bERuUXcotGWaYJa54s5nYhfZ4GDpq5uVRn0RMkZ2OceJXI7PJQgq
MmDrjor0M0pM9oqk44To5UU7FWB+QldJVajgwIg5/pRcgu4Mk9qte50hAW9iHuk2
BC0KU/ysIrrZv+b8e57TuRf++4AlAKNcU+Rd9hG2HmFvAPQJiXO0uJi7Jgky/AoT
jJvkm7/tueJqxnf85gfscPTlFFqHFVsec5obHxIOdH9QFxuCBZ0tZ4dykyTYlWVb
cSLh2DLUr0qPTABZxshcYCQzdjepkZCX8VDnJbwp+Iy6C/knXEwOVQzTqqL5CLrj
QzUPrD+doHp/yOsSJhCEXUDEslpNHO1h+/sJeTCeDZJiSOPVNSM92XbgluFoSWjo
tHyzqCnCKGuEVrgWSbwQ8uCeR1v6IT9KgxyNlpoGbentLEDP4wgpUqzdOb2fybT7
A+73pT47qXFEywmcg/lCibrSHjEBkc6ed8OiaA8p7JOL4cHe+3U3By0ZmJ/Y56nw
Sfu1CBMQzxwHAr3H8GvJyqo+xOvVh8qZ2tOhEO+rGL1dl3m/eNM/RA1IaRW+cMCH
1aPnRdtwLWkYAPj1jo3gbBa4kAeMlwSVkzHjmxl5aQ1WgfvNnvHX4eGu+Elz8aN5
iGEmhcf06BAOGr04Ghji5ZjX7XcdGvJOhTcPxW4j99RkKnpzaOWZGQ5YHZMUM98b
hsMu0LozjjUFHWKt9nNAIzd4SXqN/66uzXTvWzz2tAeYDGL5+tBLxcAOJl/r98Fp
jwcxVhA2gLomNR16FHMhWIo0gMT7QZyqoyjSUhn2osUT9MSw+vhRReixMkQwJCAo
rfHDCVpGfufP9ZiYnWwyp/hEgIw/YJYhDKLjRpc6i1TZhPPlecGH2w2QO5NS4Okg
AHcNBqFb2rhByK3v47KfN9Wsx+RSs3gzG8jpD4cOv1L6qUrD2/oPvr1LOFtmxW3L
ZRPQDKWpTMq60LbTNAJMTWPtN219yyGXemcz9F/iUgISlDc1UGKpsV9i/OI+1rCl
9B+fCP8QRgsVCGEWreFgd0TZMN6YYaKmuUvQtxK7K0ggZjsfbhuWlndL/alR7ge0
tPRq40m+gyYnecVWw+sRHZT2aR1B5bYz60LnJoJLqkyOy8mQWxozbD5hscQm6UwA
u/t9P2yyKr1shbKO/b3uJwd4e1+OT4m1hzUNE4LM0FYqN6LyAh5ktqoKQQnULDBa
K5rY3tBdjuwTg9dqwVSx3ISRucX3OtalOGGSsi527Z6yFehRsIjhfF0DnS7bHf1E
4SQYuTCILkRlwXbHIXVHRXf9byuk1Kqkv3hb39cATPqAUHy87wVfJRQuTY8e+HrL
5MzTSOCragwJ/AeYLlYeepJuiWyowlQ3A4D2NjifrPWaPf3qSNxpsXPffayCxtpp
qLkeJuP7n7YmVDONVO6BF0UmQ8z+ly76w5VtsvQ1bjCK/ArWuMEqhYL5rDo6L0Bx
VN19mmqhGUSbgh8i/2b1pP3FiEy3xSqY77GbECloRFcUKn8XfXVB6FIGdrToQVUo
MEWGF4jjwYrts9qREhG78LlHzm1KRBnUUAWTfho208KCblBa9zF1bZywx/4Ynhfs
JVpeEw98VaGwH++ovKHtCxliFZkBF4Jk+IikoThlwF8QLC0ncykAuTJoNVA8N4xX
jvmT7jkn0cwlP4RytS3GCv6MF3EAFMwDhLFtrx9dlEDHBASnIZiozf8DXMY/ku4D
umUnAnCElpp9lFPlLUIzkc2MABPFM0vPGj6yRk4w6qWdqKCwtab8scRV11KrBkd1
49WNKmf3qim0+QhWUOHOR40+5ONr7jrONWKzDPCbYMMUAxAQDm5zNPzHto8fvNKI
yp7zmxXKZpVpZ7zPjKS5r6arMXP/urSikAvD5NZBxol54vE2VlspVAmScf1ewGAT
cnUhCnp4/594JY8ONkXvQLcGGJzrohi5LPA9xXZdMXjEy8UnlrqOHuEw/hRjLfLp
hQCEZA8zhA4FCTv9rOLVvkC+qyjD4rF1d1NEE58YOUrlb7gRn1Z3C4fcOrf0BAgE
ruAZwJ9dv3oTwwndM8LUy8LPzQxBl2bzxbrmoLUb8PpaRfVilR2iI0+F7cy6q/Q0
cQK+tZz9pJvUo6wk/5MBlYC9oHy79yIEldeW3v/hcaq3vZNvuwu1btK6hO0uFwpl
sVGJtZTXrmXyRdqLdv3pyHanhO6s9TrrnFzCcS6uXETHOdQHFxgYrhYkQTY/9fwE
VyOpGAXRZArDINAosznRfkzEZQ56/pYVJtaOI3idKYmh5EjhGz8HkX6NRHjmtXoU
j6DS6m7Cj1VMoW5ZrGybOZsiUyz5gW2GsfM+NuLSLcemsoHX1Ix1sNt/czuFoBVm
2P3kN7qMPUtjZoGwdtzhHSTormomrhKwql/PheTvdWKTsXr6ztIrfPSHurOVWMEi
bwOiAVy4TYzrFWpzmP+8MEUOSwFAEd5Oxu1Jrsc/y33I5u2msGhzkbyRtSB95N0P
mBxCcJ/FcabTpirSo8CXf0cTFIkGDGWOX+kOciwOCvTBoUMzeJCYqB752oPyeVSi
BRBEznP/PRmA9Zh2CJqYb5UpAWP0Y5OC/jqQrZpTkiCT/9ClHVNl7Y6Zy6qBe2sG
WHOnyEXBGH8zWDFLXr9ucGuBUDTBvKmHs7OcC3cr9iULmo4WP5kJVq++koFugywj
CLDpmsp6kt5s/402rRSUN0XqScU6NaUBwveoeKY4eEWTrQPhSpl4XFs7YhYAKrNM
A5F8Crs9RC4L8QtnzsgzuwF4TV6atAvd9SZFQRbq+bcuTBOOSuXPZSIbcxlMkwzD
q8lX0ltR2TqT2dJSM2XCQSTq1txjHl39+YZra5CyIEQlJFXElLHWIDE2IpSF4j31
2RyS5tVz9SvCXnLArcpnvRDwFG6RxELXGMU+Fq9Zh26BLIXTrbGwx5hHlLRW7Cz6
1XuKoefI+U3piFRWgwulcCKxxgxtoHU0PIhJoqGOcZ5qYw0F5eLT6Wa/PdA/eJ1o
CpKWZYyPQuINmcL5ZQknQFMZajLJnsrkrwRy7r5anq7H0+II4DVZYURGHdYby5ax
RxmdynXsOhKB8jetB08D+xTCIpNN4SHdZX5AaF6R23R62I5E/f1huMT67FBLt1Vx
rzWtV45KP0b+iHv3qPXH0Wrw1W0uafzmreXi/+dhHJTDobBML0e1tFTuTB5AjzIw
NPKdPhN320mGJgbh0R0JJpjwnRfYfnWReWp1Ol23cSs9svIB7pW7DjBx6TixSYxC
z3g1NhGAthdrUxNo8S1kJtFF2BqXA+n98xm17LLbK8AW5h25PtCq97osjrersBI0
ZAxx3NeaX/oqAjFzf0YIYZ/ZvtlHrisQzr5tu57ny8edLNfUnVpw41ChfNVQtROE
i9Jn/FVLdURx7O/KHRfAEITIiAqWEu/LLNElxRhH6SA3tGXespX7JaJRrO7cMuO3
5T4yLTZ26HigcGIR2OpNcw+26pMrIMTovMm/GDIp/g/6+TNAFTXRwNt6Rg7pPJJa
35uwvm4+zy2yZhZxbo1BqYBQabZVtAAZ72BWReR3thlpLRCqI1e9CIvz8wFzmT4l
2DVY28SPDby5LrI7RIozFV3oektXm8CexUfX6rOtA9tV6hPVL95B7IJJCE+Zvrmf
56id/CB7RdkWJo3Fo1IWQcOLbIgcW36CQz3srDLwRON/bxUjGTdXkGGQJF4PAF/s
QmR/fWD8C6nSO2SNb0BRbNVCBx2HNR2Egcaz3zrXVdsaiytJkexLgbcGu0P3qWzA
xz0IJVQlbGHaYABFSxDVtfafEJFbnWln2ux/fKVPnavH5wbP6tv4UiQ8DzWAuQ+T
AU3RccdxdQ209aq3oU2hL2avVCj00vfqxZ1HHzcD/Ga/DiR5wPUS9cTJM3Z13UqC
1iaFecIrrWf0nC+JZGQSnDNlHTggxP5LJ67ieRom6VhXkrgAbNEZKOB6XGzIh30/
aEQeedkl6oS+emNS92yFpH82n+gsq6A20hyVxhS+kU5/u4Y03z/jFSETUDoR3Ol7
GEbVmakCwD3SnQS+BGCopCbFvCiiMXA+CWi38HGgKVobVUddwpTrCZm83OoFK9Lk
kcw+9sC0Hue9NvOKkN5mTL1y0M/Gjn7JqnzsxGRKx5T/tJwsGjlmrJqveUsgPJ5J
1Q97UFRp+K8z3k81Uzjb4vdnkmKLEEVKteFO2TEsf5wJTV6SZOCeX2+wSJfN6P1E
ml159buFLa0gmR/oK5OpLkTVkn9NeVJKAqiG2h4YHLiacyvWPily3NIZkvkRdE9h
28YxviBXtz7gTlxaRh3q0FFWHpjd9Hi09eHcDmmY4qBei8F6fr/wqRpWbD5bPBiW
rzcYxLGreRLFcMLTOCWu+rLNDicuqx+Uao0QOTp7kbA/carIwOgkFvF7wEBHXSms
//HHi8Mt9Q31Xund/3cjr9DDCYP6EAdLMfKkFDtEkLyp7kjTwTsIn/10Cux+4yF6
NJc862MvxjQ+WfY9zQJF2iS1yqTgzDOh1QNhT4wDvJs5KWyg5csInqRUghyFDGiv
VBRv8OIeRtk80V78cYl7YWnTpxmVv9d0wIDSakavcKlupbw9t9XjxrplHK0QgY+o
80aeSQZRu3sTWdLRhqpVGc6siQuxa7xywr1pXgRT/mftzj0cvQMAskCMNKJBWxJE
oEVpMstSDJ31Ug62kxvujVS7yak+1Bokn40RntR36Ds/Rm9OOMYa19z5FDgEildf
g0eMUeN6nD3cgF8Yw7SL/JP90SvKk/7JsZHvMOCDD7x+lLxvjXLTLfrSZDTYXljM
DnE28OVd4EPAQMKTk25VM+6WisMU8NfL0T3qRefFwSQcvWGczho8q7fItdlVzLT+
DFAyYlftBeFmseTAt2A7cy8kBLaA0B0DbyvT7BMSXMMc5j5+92V6H84GZAkHPELg
f5VdtIf/XuI9DbIyKSsb9qUDxQwg9So6LkjPERzbOG2HXVPUzPj6eH7p3xjU/FTr
R/g5opT0kuhYH2bFhgvun9vAub5+G1+MO95z4wNbMAwuoekS1cbOhjC+XeAQQT4t
aXoCDyRFfbXmdosuPZWU8oOD+26b/XBOnSuB/bVDAQolRGVEjf5MWA5uHfH/1shd
HHQV4+hircQzfH2kZHsND/ekcHRdlpAAGm6tuXXaxHzacLEbFB1UgMydu2O/i+9v
1mY8czc+W2nWxRSoijXCJK4ks6GosWWyIG6BXKCvSwzsQKqaIV6X4BegA5sxja0F
EhgwWQrL4tU4YeEuLhg6BAbDuHMYuPW3rMeR13WUq5oARkfHSTodLomTJ+rmxCnL
7hIJQq6gIg/2KWdx6o0Xnb/LYFr7Hz+HaNHya8jQa4wtRs28TM5aP49RhH4TYVBV
8kpo9WM8glTPA07ISxPxrBbIoRyYjbdy4JwmKg6rSJ/h8ceyucUPm4rk/1NqPBGl
kljjyrzgU9Ibjqkb26MtdkIJVcfEEWDEBxgYEdktsGTuRpMLCl0KBNPFvRabzK4H
K/EB4bvQ6kudSwPD9wYOLjhJPwxkDs1KgF0Kr+NtxVpMGZywGUYb2G03lHxYrb7k
QrhvzKWX67XiX4tHk6VWo7SxLKEETxpfk8ZCDgCngnq3iQjk+eOS2FWJWJXgGGPu
3qM6qQlh3KvQaoSge8izBkvujbjOuPjd4c/u40CXEvc1W9NWtK29CYXsCdUmlHfq
NRIvNLnCLAByyvnW5xZAeQ8lFeEJEDdE/eEIVuE1ZOgQoFWbgHg/6lifh9nY+j4P
eQrNJBMnovBPZFqUJX81SFgP7c4UdQL97YzkI6Rp8b8+y+TIPqxZFs/sp0DGKG94
PeVY4LUuVKyRp0kqLh+AXGMQmVH4A91zdPX11YowGDBS+rHL+LCBlf+WBSHCvYVp
vgqaucg8a/xz0fpSzvGp/GUwQn+ChYk5cCYnOpPOnXykCyP4mnkzspPgWPHoMW75
imY95jKzIMlLDJntIooT+iIE1RrqLg6QMJ9zQ/PhWn+2dJBzqlcN2HUu0ievilEg
2OIIYARhRDcAdf2bQZg5cBulCWi8zyeRIJboMPkYZtHbX7M6zkeLKSMAiKv9hAZl
alQapU7UcHjkNtzjOuyPuBfNTZZX3+RpEVfuqgtN7KRXEBIJa0HBF9sxQpv81L8P
GTbYivzEqNHPgFUpkKJp/nvI3EqehsWUIaRJOT2bzqFClmpWbVYG+fk1GAt5U7Yw
5SzqOyq58sshlJ7tKok91Q5zwSJ3s1MrDvO9H9r+9Rw41C7f6oST+y9Q7LFf+cu1
+G7cgrFDRNnZEDkt0oaGv/37vGgl5bExhietqR80CMUNmuazp1byZ9h4pPaYA2qN
+1mDwljVgwjpNtq+HzFBbdxTQhp8SsXPHh9/7QCD3zGBmO+fqvKyBxyoxtZBZDo7
3aAiAk2kr4gAWJYR5cbk/+f88JvfnX6UXaEbROgTZHnUNwLtNYvspfc2thofOidN
+yjgO6ZlHl8+VtA/26ckMjeSHU9+Ue6GWCJNDRew3LoJKlwEBi8doKaGGGgqKQFi
5K7u0mrKp096wWcGMrZXVJQ3o72Zl169NVgCMZZMDizZeP+oxFGXn4AmYPCVj5GL
ua9BegBQOA2XmMP7TqCq2WrsXKqALR1IiKf8u3ncIsp5kuJMnmxyC1ziRY7rb9qV
crrtHG1JyvFb53oGmgGOF3tLHQ6XWbAjpRUS14actW9qPWLPYlKvexdDvXgLf5OF
x44Cu34xLELv8j5dPCKjMqTT2QN61PPXWFNhW93rsljED3aMLV29xTnSae+nwyd/
FtGIqVdPGoT+/j/iRNmrZp/sB3UJol6Cj97FYLVV/cubADym4enZ+BLPPFMRWLdM
1xycfe43SOBS2mnJSVnqdHuLnGCClnygr04hBGMDbkI1PB9mUfmD0KKCpuZkLhYd
zPY8rUfBbSvK6uJ3HrifoMJdZlrh4gOzC+FVuIvFzrkY+1eTQ+UniVvzFdELJybd
+E4SG5g88vCUyBsxLGooNpexTgbf8tFslr76rn7ced2mUBgPQ9AtNCGRr/NaRnjk
DiKLB88xAWw1Lwr+ULbOMeIM0jRehzrbM66GigcMxyzB76pHW954K/WcAbYiBawn
04vKRZF+mHFkNrwY9MGQ/jqT9tg18OkSOXqzyaCHRwSGK7b72FKla1+jajccmDt5
ubDio5INSZUAbrBtBi+7c4OcBc/opVKNa1U28McKgZtOnNurvjatsqUKIXIXb6kz
wUT3eEmjN9MqJWfNA1VWUlS+XQXdj9vODrfVvnJVjt56nirKhuYiTkojiONDA82g
/jOMrEt79213GmkmvAApcc7epU9B/5eVP+ZCaHtr9/1CBxtM3hOnilf2oagkUS8I
V+qSCAo0VScCBrQeHCftML43v6hD9hy7Lh0iN524tVTsI1JqKgB5aTIem42PCCOa
gXQH1K477Ix04NVcYMX3tozjvSZottBJ45BqLpMTMc05IvlmXKNKbgVQcpIm0sH4
F5Y7VTpKHk/yMJS4s6DF2Uz1jdsp4yIyXybiaPyRPFS7TYKt7IvMi9EnVW4yxPl6
YQB2O0+njWcg9yUR22VsSUJdB3f8nnKFL6IM5re9wPHFAgTssmY/Rh78slNUiyUA
KEvTRGsJTwPqgGWOcsZxaQ1bOfLJqsAz2a7597LgzimkqBRTySqdiGD2Xz7T4W1y
Ho4WW3NKWrAzOXZ7sSfjV8trSr7EiVtw98ktBwJx0B8JwocRBkim8hsyHXSPWelq
GVtyzftnsD0ihvmp0/ePy20GSrYuUHVfb28/hQFK+OinFbZYgippDkQK48fUKJRL
LsIDMD135BDPsUK5qwxW5zT2wgiAL8cwN/Y4XqG81Wi/nfAf4E9VGfs1YJj3rr6P
RdMmjcZ9R07otJvCa8pxOszuiBxJlFHRQTEti6kIWEWyX6MqL1d7HllKEkcEtozU
Pa5DdKF09wBlhwemaWEZss8zKj0a+5C+biOqpz/P25/nKl02FKDmfajZBAkCbtaM
lkyNtKK8hwU1C9yIociOI8iXu0cE1hUEwDE1al6Ame6eScWZ/pb6m+2Q7HtL8zZD
vUrPNsLt8YvM3ZojB1c5xQMitKLNUJNg3rmXPDLZMRPIxvnV80z+i/rCepJ70qFs
+4mcLcdF0HsEvtEsIsfQTWplokwQHLQ46hG3pLx22iOE0l2XCPQHsZm0CVAnn0Kx
0DOmevnOSr+AQAEgvovdBtdOQfjokWMvgFq4aWZEm9njQ1UfRNX1z9BgAR0pElxt
BTXBSVJXq6XlMRidV88Vd99uwQHWSXJX/Xl/5EIMbrb/mbM4A9Kva7KT8ocwXl7i
aiBtCHdevmq+GkX1VNECAzFmL7sQPlzOxMHrtPjeCfUf9NU+wJYhubnRjnCcsq10
xXJiwzfOC8ptbGU5RvgI9oR7MLxH2ySkX5hjRxgwbjWehT52+KutQMq7xK7sBaeH
x5IveNhpegInmuQxoduRg+Tu9bO/mXHJWW77FHOOSSD6KKs+U6vMFRNAqZygojrE
NWkDJt3O67sIHxpluzrboFMqAErtvGgY/GmYmn0QEdKtAt0LpnXTUEFdiFQWp9C8
bC0e5TYk3qGkrjp6mw9LoV3uYsde/up1cn2S9eOL8ZAC1B/QT3KxvcsNaRDbSnRh
18tInr+DY0ENiGML2Cxv8YhqRstOUiMquuaCkJ8dPsJiToJOxEIEGlWPdaxpN9qZ
AVCwjEs4qGINQf0Z7LUQfqZQXvQ/Hc7FwwJkZJ3rxbBbrStOsHD2+0WfJYbaXth8
yZ18omEXw8kmYYrRC/f1zI6xJh3AQ03oDv8dO/ybc3VQd58CX3Jo1vnnPjbMhoHp
r62wGMI7oSKgvZZ3Iw5+oKu9VPfj+bF4/JDFPppdSCHdqtFl0b26KhgVCALrsLsV
olodDghh4FzUSNOskRK7QscHXLzEupD2wqMK2IUsRBzkswbz3DhXn0911V5IV2Cp
ACDs9R0zFAyGY4Xfbu1rQrTxvnf9519qm7PyTUgusbed1gc12TpnNBe5qxIDYy0g
fgQoxdS+gcu1yZh+Bd03OtQbeEPTDzowuvibBvMoBrgXxfxmS3q9aFDSLiYFrpvn
hpm2h6Qi5BxBLebvwmxy7ppzk3xBoAGDze+nOjom+2+Z5bs8N39b2NKSAn0iAP6d
X4oGCVlwGvp6crLGgJMQMPMuHtlGyyCyRb1NdSYDECGeVgH76vTCOFxlvSQDxxWS
eMmdI0qtOvly/eRnbush7MXx76DobbBYBUgqHu3HQBmZ1Hzn1uZOEP0La3tYgWZN
pxoYFUl9Sa6vaZDqYTaODyjtRapI+d2OEgy4Vg/geP4fdgkrT08J7HmB1xHUue5W
no6h6vwfL9pCBcWLH1ZaEgc+0oyKNxxyDLsX1eG6qAcZn8UtV5OvXqCBFhl0ms93
XPBIqiuEllL+MEdxIWxHu9reGImyEj/RgePgJ3WN3xJCPNYLsSDI/5aU0v7gNAbx
zUT52jneN5MjZttaQQPZKXrBhoJADUXi+rcMMCNpIElUxY0EFCmPUc+rT0Dp7mUq
TTJZH0niScjNIeDXHmPKC5gCfMnQtPAaR1OacLcAtmEcgigKv5KbIx9y/stdW2Z4
ckSUMoXKgaiFK2+nxSb4ZXPCf3RRsQuOGOKOMr3e9jKWo3+nTKcDRHEEmtgq3ZBI
5/AFglQqjNoiEPvj6RmiWMwFFfGRzR+lC/W7EpktzrIBiF5X73b9QBpCYtAmvmdx
ClbAn9An0QVhkN/KqBZ/O+9I0oo7fR09TWV9HuIZ3+VjvkqnuumXL8v5R4v/PU4H
HM4bEDayY0DR97+GY73FFOvK3IT06ov/N9OGVyjDUmYvHEQOajMQeU9zA1hqxAu5
9FeEGJVCz4AyoLee6heiPc/rPgmdpIJFZ1H9CuZpqtippApY0pevA1/Td3VsM84I
xt6Ki2fEbAUPVlLfvMaKLZ5/9J36mhyu63JSzL+AgFnaNqjOFUDU0uPhxV79b6YI
45GVRqo/SyCEkGqd8JhBdLcwOJ+9JBAAny8b0OcTYO1Y6Wz8em0TZxcSb6EJNV2V
QRSTFZDv+EVNnCw/XwbwLB03s0daWW/yXQSVesndv409Ohu84BvbZifmTHTH1+fp
+yv39x6fp69hilYIUDRF2p06vQMV+MkzYElzm2AZBDXezpvOFDw9g9Zjl/Mx2fNv
y9RVMSQKwChtOtaln5cayS0d7NGkeW4dkRItcgeYUwBw5iOZBvf9NsIgTa1aEZe9
R6lP/aGX1YUwr1mvUUMB136OX+CEsN2a7vNplmk1bJmBjYU5BBzhe5kIwB/u1btJ
An8UjwvHPlEeImME4IJrfMUApl8Qv6KB/Bdc1FAN+ef1jXlbXIZlR0LXVbrgZhkD
0kSOLi+XpYWhbzYYpEW9y0JESnxKxFm5ClsLVUJxEu+KqYp+tHmd8LTJ1O0YOmFB
Y62VlTGqRewSn7WLs93gV+7PETO1PMGT6/lbBqCjqU6SZJTMmwv34ec/sc87AVxO
140115tk0QVqB3VSTwR0HXU/T+SAMUibo3WOu5SVqgWgOEdT9xhbF2IOWA1Ty5PE
XmZkbISI2WiteQu716vvbE/Vz91AydX9ufzMSu5YkYQ2GzLcrXO9zpJTNPSoXQ49
nlG7yYlah7IQwlZqsgQo8zR+7keNOm8Z8eeEKdx1eHeZQ1JA17R1IxJ/SaYhAYRZ
m3L94T3MlkvM10AZwo6mU1dss4Nidzd58mAF/zsoQm+j4U3WOmvjqzM46YAFc0J7
luX6bZF8vYmaiB8NezcHVgEOhcMDQkY6c1k90tMHAF+a5gzUrGeDSEezoUq1iAmF
V86Pgarf8/25TE7L5ohwL0feUJCW6Kc9wvr1FLAsBadaTm2GydakJQhm9IRiAIYu
p/pSP6jpzGAQrCjkn9w/ww3Y0dYCoIfsFs1PtklpQBGOVWqGyziSeEJs/2tsH82X
+RenEZbxRR6MAk1hxfdeN9SImp2x+akt45r5bwRaod6T2YiwLFMZPqRQVAYP3Pan
OsALME+V+aK/CHIFcg69MLlettpKeX85du1ZAf/tWO2vVceAO88gLjuc/7YvLyq1
PeR55LMYIiQKqssJ4jrq4iuX7yfsGVCUJ/dWWV89qVj2ZWce3C6dfcWZXYAxGtmE
2JsqnKY2nOJ81z5RdTbPvo2vi08KTxZ19zojUNhzAwAx4Gi/fNPj2oKYUKXtG/MQ
oPbcRf+nCyIk5hZIB7dEYLcGEGXpsXPpLSFrgIfLIRTZBkAQCIqPXUDtlbw4Ka32
GwKLhTSkDfIE2ieYzer6GA1rs26TXZyYcpLXe3gh7IISDQBMD0ocFpb02tgi++7T
lLjh7nZKj8AhDmUxx9IeYNcDzlX8HwX3Bfdgjzq+ywtmKUalZo5qHnlCIzSCbWZO
MFRD9ryeNh0nzXKpVEFt6645jLpEuNbVCbTHMba7HwpS+rv6WxG9UvDIHpR3NW5P
TPfGgGDYi8AE6gGicuJs9CIMOQpIDT8ivr1P0HjDJZTNR5BRvLRBTi8p1i8SAPAm
xbv8sGgWcJVLGfaa1jd56fGFRfsGe7wlq2P3g93sVhJ68RCX459oA8STnjZbhfVy
36wuPm5/t0Gm1Qbzk89jCifeD2ZMFXmQtNn4zR0JBHeLFBtW1ROLsNeamoS+twWD
PnUsUFu+IjpuShqKSIUNcTb/WlKbmyGLE4tTLzvHtyPFuu7lp5VNTc30tgZGulmZ
gzHZcAsplQN+/7hHgQLzeH8npRxntxknHu55UtAZuSLB9gNtj36h8qFgmGyMHm9y
DMBkiNxOi+jJHZtwvtJEzRjg3vLr/rJRHpjP0wgQsjRUsia38SvBZ28ww3QPzTnV
7FWOwG34BSyo8TVslP6xrj3t1OcweWEJrv5hoUu/8zoXK4eVYo3tyGTQtFeOn3sn
cw0jA/JDBSin/c+n9xxL7bSOOj3klEIaC9gNhw8Kkdta4IRDwIc1Z/pngUkm9rzp
eO+J8aA4VaMI+DcDqLVqdqz3tcRh0xWnY+Dw3EwuQhByCmXBu2MteBaIpNtr5Ekb
u2d+OyEYNGoLjAeE9li41LW9Wy2nNgtHAt4HmDnVKTAanUVfx1pAoBts7YjzcfSZ
a0EBct9tKg3O5fJKvir0li1FKjH9xkSML/Fomos9qhbWjQ4un45YZeY8aLPqL+ok
h1O4+Lnm9CZlFVVHyqmQQlnYGrgXjQfmJaL8CMp6sTi/Ud5oZhnp5MT6H3cmLGET
bMD3bnY2e9EGK2J14aoQpeb3l5HW+5eFbaV+x0XgHMc0jZAtsE8dCTEXjTgi5Gpg
sDulfDPJPc+bER7gD0JHo4T54AZreEGJQZOKGFALa5BjXEjFBu6a3YmnYyOiw9Nn
hgRgr2RlIQBDppSun27yfbrIp3Qe1eG1/KtYsfaph4k7rUeF3GQoc6gTmUa/Nw24
hzrYmmaJ+2EdaVadie3ifUp1Pthgxr8Lux89axHHRAAAz0XPFLyQkGu0vMeJGbWj
MDq3HvFxUERh1b5c9jceBPg4KOs7LnGDJh03UGqqm65EZKYWnKuzlovFmSiL3gw2
oifxCGtc9OUJ19NfmcBh8I6+khl60VBoIvVME9MnC6sCX3XlSgPThIb5E/Rip5G6
Km2gOrTmDs5MIJTtqv8ePQVdBloJALpqNeQ6zhz6YkztoiZTMi6yhnHl225Zr84F
guQ7TntacLSMjLdn5vNR+wyHu13iPK1nTw5oBLQBKNKInEL6a2styj+aMettuNlg
dATxOoTiHTyB0Ru7VNk/nMZT+BKT0UjOyh/7Ld0FUCg5vehJtPOR4DUvxt3UvDwB
dICMe5OJ3s+Zuosc+xs+ZNdxYSeid0ziYKz5c4HsiifZecLoqzQ2hdktgftinmqn
k4tLx9AdpZOPYECIF6e8dbKNqd0cpFyE+8ZBztP04HBmuhWMHvVyd8K661j1OWdE
5ZXY8RTnDpdb6Divy+F8lzrnsruCPtq9omdiFUD73ef49usY2oi+9NO6Fv61mPYI
bt03+CiwbGB7FhGko+TH3FFF8qhTeqtgsDg7P119xSV1qQrz5wl5AFtbKK0v/ItY
pxS6ymxD3Jv+ZSjwjVzBLBdzH3pNWfg183otsPA7k/KiqjUiYJpBii5+JDoXfTic
iH2pm3fMsQF0oFGo7aRmZ+GLR5M9st4TkIyrntAIrRWA5KlJYV6JNhUIB7qEsxmT
V8cViU7nqpunbl4g+bimkb+xymu3Yyc6yDetU7Dgu7gk4yqivl0e19tHaII+4MB4
0HTkfvwQItozfOlFPBpEPktrzobhRm7wQCVRe19Z4cZlbBuc7u1t5EvUjz6PHNm+
ngPAK79Qr7I2YEC8h0BkgP3XyCSQYKYxScLLQz6hHRMYxoe+ppeXQjdu97/nYH7u
17a3BM/q5kTnSCV9pqNEvG0XX5cEovSw2ite5qvL7n14ZNEvH8yqOY9wnGDwexfk
XiTM/Hx+SIroOm0APEeg2UlRn8EnjoRE4Bgq5JhVoZurWC6Hl6fYItW1vl/C4Nnv
tuHa8xkflMloTlO1DytG+s2jGPEp7EmLlkv1ohFY8ESSH2sgEezBSSKeBd0TI94o
p51cGwvNKl61DhtjZIlXxotzO+JEKuA3m1sx1Kb0sYGWoFrs2yEJhjS2ghwc43s8
huSkVDqe9j2FyVqi1JvYy62e/+SrtufAtu/bNqOGy0leYXCtdzIFIuQydhLJl6WB
sYAnmEpB3VveSaBiy9EoQYp/FveLSYnAvU5j2tJ3KJtDINQWHSZFmqRMlHgfP9r8
EXhm2ZajKa4u62s70hS0uNkUDLJgGSmbk1En85DnySJ1t/2k27diIEuJTTBgqeNI
TbQTNFsgc3tfuBFFWABS+Z/zF06XHWmmpYjNFJ9RRRl/87d2WsZfjdBzxdGpolA/
0uhrO+O8oTBWRzIszqndLFbsRIGakVD0LH+ZSFhDI90fDCkt8V0c4OlQLo48Azb+
xem9w01OBEWCYl4hwLgtjE+uubdHd5co0d4SJ1VOQXqwuSw8vsh22KiFD3krJ/h/
IlNdDu4uBCdVtbDRl4x4kI8AWKUwFBFce4SE+prlce+SRMXidDn1lQdENo8jdLmk
tUAC5CHOke56K7Gc9TG83/3ZXoTT+qXMtahP9xpW8jkR9ArcdEXfj3VZ0gWIlDnO
698ywwWFNuKOy6LdfDFLc7BQJLFPGgEzsDXMOV3va1zP4iYkARuoUco/yErNRHxi
WRgaF30puttdzMJzG/B/S5ZUcKu9SCtiGfzXxdzWGoaKpZ33otdrpkCptTD1ednr
GmERlv0gkm/40jyYWbpISq49qZAYmQBVUjK+NmwcSrRcoG3o9UxRcrBZyrwJrY3I
2wBrztap/488vWSx7o+OoJ0DT1HpUrUY125AieI/j9wZ48wCKvgjC6nLBIUE4VBR
aoouwrRBlIRn4N9003MKx2ESo83npRj1rsA/wRhxaI4sdY6eRElxLAcHbsxb9SGR
tpPpwxDBC4BHAFOvF3ObtrNXf1sM2gTm5KzRaFxoxDa9ZXEaM0Pt9ULvjsolHN3s
k3MNUcUhXt30frJ2lBAWz0pUFqlCZQ1cKKvf/b/WeLRNzRK0Mzb/gCr/oDofI1L5
FMTynMJ+V0jn2rES5NPAuWVhLZJvV1WG7g6HTym0wUpv0TSHnNCDzq1aAu+13YEc
sgml2YioEhJgVw4wnhMWpp043Ntf16FqqeKX0ya4VuAbMaq50X07LUyJN9EKvcnb
VUuu+XmPLlSrexMhkpIZBmRGgvkOfljqmLkEgLQ6eOsDAuWAsCrpYMxW6tXPhrDE
Kc12/ZNN07eVk9P8Jw0RuQMfsMsCpj1pd3EBp6XqBuN8MoRNZ3fdxKYsqmjDngeD
witKUu7MOzMtGkTNxcSYMNnA/6d6nRDi0okHoO4iHNvfR/W8NX3lCLOY7hCViUVO
wCZ9AETuhCQwgF35YQ4JVWMi+IpusQYnyYtPuTc6fEt4siWZAozN1C1mriHrtgKg
+TBYlbczc9Y5DWeugRqybOsGy9vIUow28UTSvVVMYJSGXwcfnKeQLJo+QebJP0oq
RkYttg0uPsptj0kPzFWmxHBthoInGoY9Ooc/tR2CM1vtZkHDSfJ1hdDUqd1OL3mF
GkUpZL3Teb4Kajf3BnwIh8ftgTdxpIXt0x+KDYB1w71S+bvnSVI1DGskw6djZW69
FCJvbKvTS4sU1RaL+SrZj7vY7sVF16dThExNK6j/iPB1zydqHJ/uTzKma6qPHjGB
/ZypofAhuIkmp1wwNgu0iWFZT+bc5Xf5oLOyZuqm2ahQnT/o+mqf/i7TRf0A63Cp
I2dB873CHd2ELNkwqjMvsryroX3it0WHycrbKwkUI+OqJnXvdB0QOvVv0UQrnvUN
ekZ8drpqFRiyeJBQByQsIccnF2bYuHoRzELBc3ImLWaS72XAtMBXXixrGonJ2Siz
WqYopPFJFfMh1XaqOIgmKtBW9IIywyfyRBHxMAMlS74XmPZnuCoFMGIQw3RuMbvQ
TGMFt+peMgO6uLD6EJDg0IxzCv3lpq+OKGuwz2Emql6KTS5X8kk1GN76ayC7G8sW
M6aaZ8h2mhV8guqAj9O44SQrkzgralk3TEBkdq30b/V4MqXNNL0kcr/SKannJLf4
rnUSXLZ1okCbnc0VbKsVxXxcgudXlB0QVbbzEonWKBDRgWhMiQSShs/EfOiQDakv
JVqW7rpngHS43ps0MFQq325iJeK2qHOgNywXklbKfG4QUYlsqRatVXWMdWjPRD/J
3R07e4dlCHDU/6WultecTeWN/9DESvGy+3UAF4o4RfUpgFqMA+si5ovkiPwApBDS
cgIirGr2qTJHOgVrqJq44nje/btdxypVN3SCJA3dK0c2wgb1dyomy9ex1zthpg8G
LZCk0xPlVzRWYkx4ikLmLxD6oqoZXrvVqJAW9JsSMH3m93vYJ6ovTlcD5YwxfMz4
Qqyto+5NuQ9qqqQOyVR+cB9PQCW3TOYPxcQT1jnyA5mInREh0yOIzs5b8j6CsxLJ
Ljd9SkfcDiTT8PT/xgC/cVURZS8F39xuVSddCg1dp6C0fRCvsbm1bk9yg1o0p1Cy
u5GGoveZ4LSZ6NQ0UmmRJHNn3dzpB+oeupsfbvh/BQqrr4MHbTQQUJLNLeJOKyp5
AYmPhsILTDG12sZhFBWYiaBgR1Tvwh1hgTk4F2Uw+Wbz+MKknlCU8iQr3wW/Uxkf
ov1OpyaPEJcIw2xHV9H2w0bYwKPugLlkdbCayVTttKAu42IRuKP5sZTRnjn/mamZ
sQfWGJff/R2UN0Slaub7XT69a2kEgxOvKrNrGmqH6aVzfCIJouXZe6N64AWZULYl
vN+Gka5Eim9ia0PTl69ZfQwspQlI5RqNjCDC3lsvjzGbhf6WmQV90aZG6z2NT+dz
RE8Kbyc9ANzrhzQaqM/vHtBrVY13ihBwTkfEYOyVqZs838fdaTcIgdHfDLVi6Ltq
UPttJzFd4GCF+E/e76T5NS7//RVLNNd3H59Bm7AUpJo6gGK6fBvBdRFvzky7MKtA
/GjPYciIBSV+krkPejc5eVzHN+HfUMLfwkQPESiM4wG06XD4guO41kQMz9e97bqt
7DF6brcl6rpptM2RJd5fJZu85RjZ0dDnphI8HTVPQ32KNfe1RldsqATBPnPMfIrW
7LcqfhnYPcEv5Wv8Qpfcmu8zlIgfFjtTXfPlHZJoDawbNlh6FwFsgxdnBEYkggiY
0uYohNoKf0V7Pua+Y3q0UQ0CEYUBlR4ewIdPWafC0a88YN/emK7AXIar8ilsFg3t
0zkix8v+4Q9mE2//DMe2f9h3R0Uv9FlcGikVlZrNjHw2mflWoepxUfy7jw3AdGU1
soQMYGVxZIpMjioPaY5Vli0cEeOcuzASpzwnrDOihzDGOE1Pb0j29TWznYuGe2kB
BYqJsUu7uXa/TDctnIYmTjmmn/NXAvCy1MTTNYk41eJXrJrs/wrH8qprOYhKB2sN
L28K+SrN6B9aVrohvYylyGUTMj7+VB4K/TyUdpCjzu/cSXfzdmBxc8xFyuekvjp8
OuSigTNMyv+zBld1Smp5zWgcFKvwvYiJlhP/TgTGwak2koGrBqsP2Qb76FODPIsN
CLVXrVeQR9a6t3896kGRu1m4OyuTztybm1B6Fwbi8a9nbeBhp6uJBfBIXB2/iPkd
8aOIfW1JUE9JCyv3iInOlxOjwaFoSN/ouEPgT4Et4dqM2ra6W2Ca3V5GwryGkF7O
UoFOadbPWuyykuIWr/G/bpazs0Ud2bAiOU4YoH/tb7jiYdtC2EpafBUajdg+YFpe
z9+9ZZ3zV1zFKLXGj/oqWrWxPV6FuB36uabywbqF6I3sPPqpJASjCUBlQTIM976E
Xy2ZVP6h/MMI6OW47GWqL4zTi4uuSwGJIgm0hy6A/yzbbVfUS2+DqLxlvbHNuQvc
Jy12bOAuEZuFnh4XRFm/Th+JufXuQ+b9jLypGVDrj5UORjJe2nOrlBvuXG6jjKEQ
Uuw0aNdlNM63oo1ocJaUmMN+QuF9xbNiEq+3f2Fs71EFjHSEH533Je+qx5WySlRS
5tenzaOz9VVoMqJw4MNQAfHYyliHP8eAUzCYMxVMOJmCU0m1Ckh+OldSBh+DuY5Q
mRTYWyeFG/kt7hIROQN2K9uWezr5X/CXe5qgV6D8Uq3REtpxZt+jeiILNg/wUE3G
x0hbnsyyZ9f3t+1/8YOaxFwkg0UtIaN9gpiZ+iHOh/3jPHCyMJr0sLyrjr4uDHRW
aBbbawI2VSTUqjQLQdi2oLk7hpK/NrKQwpj+nimaKuXqoP0Wqz+kI4H4BWI3Ka0e
iXi1IvoRgdeo2nzN3WE2OvZhMtcfRhSEClKHNG+X1gUNqaBVWAxutQVgrYPxXYfo
eiT4FjvLC7NLcQJrFc9v4Blk+WY8fWSE0hrXEr/muRh3A/sGuQwuU9+MKkXyEAek
ewYwq0BEtE//TwOWBR4I0LXUtYU3xGU/SPBTBW+/GSvkrnYghZ8c7gAPqswWJVCO
zRnnw+WMqUXiPX498pix+mXYi/GE1tdjveNr1ENQfppnnVNyUY0z+UQXfVGdfoS/
9bjp58VFZ2xPwjfp1OP0wyRw6PHLLurbFlosMkxft1a40rj73ixVcHall7ojpaoA
704Iq7P8M5EF+KjtEIpmaPYwDyheA0fllM5FPP6DvcwLWyOczvht9dwGWJ+JsWJV
c+s3T2xTS5DH1AFu4A0L4Rnmt/2cgNzOZ5YDlw0BnNShhzYmJZ/n+Ou/g5GPSzo1
DC02nBMdwi5wCTgk2pr/8tq5tvkyNH/zkJSuR1uNVrYkEzhUgRHfoWkNI7UmzoWJ
FTA5BPH3k9cZwO3fXlUkkPsHhvstB7ug3IVVIfjTOBfiAHnMmGUoUP2j5Lx5mcf7
fUDCMH8PDBko4ovFFrjh+bgLttz2F2UZstaBfzfZfNuT0CewsL8vfHsYEVZO9HKI
+R0nUUn9GK042F3bLAXdtk/F6lX0pBvtLF1QWXrd3XfbJcB4bmoxEazATW/Uc7jR
zEmLtiOGE66KKDfJooo5cDsgDsEgDr+s6XxAGXOE1lxNIUifL3ot7+1dkZvq0Wr0
m4v4wjfuXNk5iMADLR4aDUyYLRPrzL1ieCKdDUbUU9jDLMH8OZ5s2GoKJqRClele
juYZPm/Mn5HSIu0rraY+Eg9AP5lie24+mcEDDZHKcNjoSMnbkZsOV4L5TgGX5F5Z
UZaLhTW3+hRrF7+k1uB7BX8sHmOkRyU0fXnjhYQR+r4Kceb0jAQ+eagWGFvPM/7t
3vtyTjWnI6MxfO/pHs9FetmXsTn6uoiX5Nk56IqqRUqVvvUn3844Brsi3CxjgB87
sik4oKiK/XiSoM/Ce9YhzjRjfNyZk05WsBttkWbWMJomEvWWTEg0fsllgFEic9nt
JdwnVaVJRS91GZ1yJImDZ1faNYUonCpge3vC9nH/jNnAOuFlBg/4jc3dZBvbmrP2
p9epBgFC41Ia+6DGGi1t84DOaoDw2LN3p4i+VlFdV3iwnw1ljlIV2Hr6CZNaSZ9g
9HvPKNvhlTcRoyFNNS6ZI+7ekolMAkcIE7s9d59CRlZEvd4Z47AtKnax9HFV71cG
aZhs+AeP5bAJrnWVwjXgcBK6jdDS1x0DeNRqPd2try5oeDX/zMEzHu8RFkqlDlUI
VLx4r9ciTC9IuKIqwDzTtRo/F0dECew2ziNbUAf0rBN8j3L0nrwnu0eYV7kj8KK6
pGP+zVAKVsfir5fFly6zYOZTsd3qG2sWRj5G57H1+3SPVpTZup/d30zeGhz7TDv2
T74rLHPLOQ15Olu/AyAyTrO4+mgZ8e7LytRMIlclUAQm+N83TR0EmQ5qmAqzgLnU
ZjclaCTr3r6PNt9tMm6uuDBiK6O2l+v6BrIL5cK1cSdHlSWVcHWLvh0y5ECFlYsY
PQXy2fVGSL1f4hhH5FMeNvI2K73SN+kxaMrOZeCQ5QosK63JNTIq+UNTwAaC0ch0
jbJgo2KZm2duz+RUBvo9oJkp2e1nSLIqTd4Hly/qs04JImAx0d8N13Jy/TB+iJln
79NplJcDhezeUctIlNeM4Q8D6ujXpUCj75o5n2McxpuZ4SGQRTRLj+lJHU+Oat4Z
7PvodYOg4WUtdC1AYtkzvi5C0AVZC/SFwrbVMur1fPJme46iFxIiDfennYMFHMM3
mu9xG3wrolBq2NdJ+wc/xbpW1BId+ZLWARWZH5yvsHeaUqOZeGfLZu+k7J5L8kuv
AGiQTUB77qxeNizfj+bgbJ9gHhy7wMU+Pgv3QWreryvB1DRidCdMnF271IC1UqEt
oXZyaMhhbIApgWZ5HW7oW6UMbeScm/P9wiUCfHWazl5zmCMOrNZHntA0Bk2uPetR
NIcH61VH/+hMVgJ5v7K/J/WOa16pK08lCJQTiIjEdpIl1Wg2yR2kzXecYnfMnGFO
c66Z8XZkvFxRi30jsfFBzHg623pj/bAvmUSHoIO9Isr6MAPnR5dkceE8R0M6bkgG
GSObx0KiStejSntqIYTZE/BN9hrcsJ5WMHvmrjc6tfpQNHWKauoNUE/YHAllpesA
LELbmsyWSYD6QrxzBZB9k94w8HC1lov6c0RcjJI8ELLKpEio9NNDQPYUkFwQCh2k
UoEyHmyUd4TtUV/VvKU1UjZbb5ye/d8QlNJxvO0A8LOU1p5s1KeejgLNx+u7b2bR
OvUI8QJRQzhK2quxYTtOxLIGB4XG1Yr22xAjse74q08WUVvkXT5vleSwfwI+yXlz
vRwTesGVCRnarPt35pab6nwPMLUksxOH8hh8xTFXzTfWZ4mg2Qc8Rov/IwTTf0Ha
AwlzdJv3B9zI2BlON6TS6neSmFki+LV6a3TBcTEgnvu9kKg5Qeon3Wf+bG1DCDzo
o1qcUd14Qh9++1Mde0RZzX5qwfq+/+VqR9XjrFCxAgl4/1Y73EqJGTkuHygL/DSj
ATa7Emz++D2cc86nCBMjcUrySCEZnxAt55ZgFNVG2b/lak+5rZlxf+vioYZp2tRV
fxYIrujJTTnrmEbobDoTUhp2cMMkSj6ff3o6YBYXo8coSnCHfGDCCIoeXdLTVmQn
yLc46Cg72JFOAlsA+rh1qYD1lodIpE41jHQfPF6JsLL/ra8eo3g2Tll30n9ND0hF
QcSAJElRyPmaozih9ruPoJJlJmjoswqZRnQm+OVuQaLofbOegQXmo2z7OW0t6eN0
O0gk70JeFGGIxbIJlWC8EH07BodKLUxO0EMNToi1kcNfvH9JdgvmrKjLeL635CnC
XaRArEiyeWAGmosl4XWYtN9lGgID8K3u5Z3M4a62HQ0+RkCF7rmK01FLN3Rs0Qo3
tTH3ds62ycF3RrCDCH8RNKV3UgSxpnfwnuwxhMPp5wepZShNqlzKKULz2Qddpqh/
My2Lfve794tCCs4Onsdg5bV+dKaAgpKAi9a5lojWj2LjZmh4+ljsLrZ03t2/GhZ0
nkB5iAedLb3bRTFw88cxGgICnj4BDJUrsuOxvOMxOUI8FOVVpPR4ke3q3rM3zM2a
G2LunHlpbur9a92sRopqEkhF6r6G98Ni1NgkDtBKVlCtCzsmQ9IE33ADKnH5/cVy
XqnjfTHLzJM1HW0JzPX7tWb0Ei7teK5OO+tSAS65QI/p7FSWGfd2Tgzvn2ipr0pr
Hg5xVnbFZduXiMsik210VYJ9yiE0SVKKUR22uLKTCg4Pt4l5xFmwLTZzjKPHX2JQ
C4XwrO6WfkT6uEcQnknaOJE4+wn81+WXsPEajvqOpiX2NmnsF4mDGZ2OBCxpQGjj
YWd347iiIxezDU1d0bosTdDOpbUfsc38I5GzcNc+HobUMnqlD3VrweFkSYB3fPjf
NA33JuD4KJn6nY0KJSLwnx7nnDxbnHf7hPEqIGgYO2hci5sg925+jNFZj0nOgqkA
tsgL+lo6MCjjeZFBqp6Ui1ppFReLb/pgoqecWIrSPvPMA4yLn2VgqMwHl+lxJgBM
AdadzbJcme0UDhd+dowK4lxge6JBnzKo75VvS0/qU7DhpUoTNuKVI039T8D91PUX
X+InCXKA7wbDoMXmwtpSgEtbs45VzUw0Ux1TQLGEa5O5i9s5Vk72MJoyrGAG6lEN
qxeaFUwllPw42y6kummKLrtDVpq1pMac0VkUd4+iO0rkd2EaeoY/zVdptHS/YQmH
dC/v9aEkcjLWg0NdxESCZ+Y2Y2S6EDb895GeXPEQwILreg/ckBlnsY5guHkcC+Hi
m8OOpRLlKwSlLAPVQTm9X0bioCbHN20IUNeo4PAet0Y3M0AOiJzLanxIdz2uT0oD
nXSY/ny9jyLXwMtcYfiX8EUxTdzUe2d7mkhh/aMmVcFwLluenMNpLfvXT8fnqcPc
frnA1HlOEWI5MU7Q5xdkpyhqwhn3Hj+RUkYivUQDMjMO97s/yKRpqfD0lgkFXuR4
qJdO5Ia2HhQiMoO0He8Gp3zstVaCvKZpeEAxrha92AjvSR+HIFsZ0cNbFsNwX5n/
FlmjpSDCPBedAZdZwp+3oPpqzgRRsoFXe1KW7tTl0OxKL45mBkYgtFzQvgxcTDXr
9Xf8k6ohTdgJqIi/zKV1H+7uwqGSoN9iniMVl9/vB2qKAND0lGd0knEPZgXClguk
BliCpcycklVBGVfbXN90pZmSJflPtQ6Towx/cIKb6ZMD6Y/S2MJ1O66XKK4zcsZR
YuhKQlnZXLlxnuW5csLAWqjOzvJtU/azU7GGsVPOU+LsT+BN47d//hikhjJRYFb4
SjDJ7RU1Dw2POgebA+UQ5ofl0xnM6iR09XvnK5zHY5sDwaSBJaDd4+v8GbVYIRXk
ecJdW0uG3hHGuSWDekgtaoGKpe4amPy9R7507xul0c4WI/2b33rXnB1uRKa9jGMI
fvdAO3fRpCSCtW3vyGjA95Z3gmxIzazRs+xCIu2xzM+fGIlaCqZ2wc6KwF8vxa0E
veSwrig7MNl9+I41vH6nd5Ktd6PI7dCggFUS1vY9QKOZKvOCza8Fz2UGhDKUB8j8
uRSWCr0voTNHoFddj+OrXUF/J5uMQbh3RfdBizSC+SJI6q0/bB5HHHKgzowt7rbv
iHzONXvDC8jj3KVRhYZBy2Fo862+ijW8FMp1uldfcrR9pIMwCY+DBSnZ2oPpRJ1t
zFO0OlSr4QgBwEBF6l3NFOTV/Gl5CWU41Ztyho/BZHaTVIDTOmVZ1qAaHkOSHsCN
GPFdAQ2u0zisuN0Y5WmCd+eKko1+apXtm6keqtLXlBG31iqahDCd8CnIAMrQX7UU
QniU8xjFQo5OJG4c5yKUE5zE/DeTxP3NrfGz5AWFZT9y96mXgopYaHCntjCgFRDm
cNJ12wkC4k6rtIWc96eMN/sLfx32KwGi9zqq052axaZY9Z4XpQZCrMVrNUu3tlDe
uFM6yqr71Z2Kp4cu/hwCXA8u3CkA496taZHI22xipLJ9AIXcgQFb1C13ZifmvRI5
MOP5kNkhHQ3AJmUCPY2qnBbRopUbSiqwVQJrrzM19WRgIF9/m+2CJYVWdChBSFcG
jUb/CCfdKj5itkWhcjXqbfB8kxwdy4ivmNsw9kENvZM5IEqItNqYoWP+ASkdsuQd
hHcekO9DFUxn/+QjNy5+LVnJrANsiOfHwQ7aliWPozPE3UlvZh1yzPauzpZu5g/O
v3FqBY2MaPdyrlR9IATmG13dEx0WgdGuFnotGbZiTE/hWLeXlAkxhqsAc3FNkKyY
v3PbVR+igUY3PneUexQqJAtXNKLhYvrpl6MGtZYQ16ZQvH0v96uNYGCzjW1x+dDQ
yzb6egktBbXeXrP5LHdacpD6MFVl6REEWUD/LHiMi4/Si5HLlQhptiz+YiYYG5Bf
clbce+BNW/T17R/a305kXlU2k+NfKKLBZ6MrXCv/dF6xnv8u/ZKWB7HbzmuSQy+i
MZic1NJOu/V/U5bg26FZhCR8vUzaaX0WNXLvruq5b92HzgwFpdr0Qqn3+BdZHSzC
utDHNJNyXKDuvd0dy2yA1QsEEQpdytBddv93Ogb0iKVl5HV+Dy6fRn8DaM+IvNXK
DtHwC2WMvo1JS8HfAB9NAAhEy0wb8VfvRlpi23W/3qY1ExhGXLUbuQIWFTnA5UFj
ftGGjRmg5avmnE6gBzDMLnrLmWVLgjBEYDpw4TYAnKvOnNiaEXgHxAeHfZKC+F5T
TVOao5LyVKkdAswum13OAqAxyteAgDtkrmNz2/cpjNRxYmHM5w4BqD3cMQdP9dzb
6wfMZvIaWHuDqDq3pKq/2+CA1hRr/LCAJ+qTtivODFvvt99U4RVMboL4mLhX4xQC
rUpXXxqDMBFk0u5/oEnrpr+Da/HvSOiWIO/cEn/WqeyTg4x6bY4DBMrLKEIWaoz7
`pragma protect end_protected
