// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:09 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tPvBjh6tvfscEwPGGiyL1byWJNajJJy/tCSthJOu5Q4Zj3zayfdtnQB6f5bSgTCi
7saZ9lwC5sYCGIJ/c373owAPrs6Qk5xhUiyobtJtjVVE1qOtgC12sooJB7rtCHA6
8IXBGkaKgw58aoAgm4y92KAP3i4JjrXRT4u83mNsbno=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1760)
V33NsbQBWP8rE326z/Z0eHNfCqr7V99WjEOKZSUmTug81EfjFe9cIDaah5emf5DD
a+YJ0cxEbJCh99IM8jyDugfQSXaQB0H8F5Dd88Q3X7DY6lOxv40+xNhN/7ImKo/h
Ouj733fTrlLCaBiNOpuF+kEMPeHw50wjxqNiZ690wU3f+7+LsoS7wrdxh0/OobrW
Bh2JKku36T3KwxvdXnBoigrpAhx5PLGhfr/9gFMwxDXtw6UDcf6E+IVz6pq2OCIg
K8Om2afMYiBtOsjzHqviRkmhkU7UXqiEbxnChWE2/WEbNcfDZrG6gXRm/oU3lNSn
BDwBdB95xr/oSKViMvCghAtgNxGa0hyAQcOiWTdaFgel2yji8wJVfbvSsPyZS4G/
8d+XYH6afF8kg8WrJub8WNvZWcpO6sxZJ+mqAeDHtokUzbG68RMXuj+1Zq6UiVwE
jWyr3EFqNkW0PIhGslXQFgAa7zFvHEWfcOgWXnVYB43UDfZsodoiD8iowHYDJ7uc
YhCfu5QropPVARNSjlM/TXtOqXFnVlR98ZcNtIFjjNi6gm1SkXWoeiSSASIidxlF
cUXAZuNJlnPfoqokRHqTsUW67JUNxgC9Brfn9UFxrzdiLEak3kzoHEk0n6q6y2QM
RfNza+5dLuBGRmN0Mh5+Hr7x1Uq/63Y/5DSvq7ZKodfU0+eKDkJUk8OiwH4pDBvq
+UJDLLyQi3ZB7f9MeDf8ttNXuMdW0obcCngeZ6/6z8SUxXjZp6d2eroNPrMhAlIm
NGX/gwbz+e7/Ugl/jN7AogylFFu+k8F8+y0Rqp0tgFymFEuPuVjDhoWjT1Aqfc0b
8jz++9UsnYCg1to05Ltf7CWyoXYxC5MdvlocQcJjjgZOy2S9WtdyF3Afsjx2Ga+1
SkQyzACtZGx/wVNClxIv514nnvMJUH/VfWxVInVwaoE9hv9d6QDZfLDt3FWZ0981
dsvk+UJYYcsXDdJHPJuFVski70749X5qger9FJEKQHfE3RlNGTeau6o+NcB7XQC0
QFvFpLA4if7aabATOb133PERG3L3MdraZl3REXuhaw0aZzD3oHcV+kULAU7j/d74
azr+LFXo6ynCqFzgQ0kme9w/VTZted6N8M28dPbfG2DXQOnySPXFBwWbOKoNXFea
3xGIi64tdONechXyHNdYfjBQKSwxDnzQa9Ojr5rRxyehZ0M/2lWHtfw1UxBI2W8x
3qnHsDGV7SkrCC7zkSDVBUN2GByFwP/i5ad+livx6SlCuwwuXbeeOfDcsmeXU6Lh
oNVV+JnReCys8PYr6qhjw0t1AcKNJScVpZxl0oWSG1MbLN+Fj+U9Hu1Jui5Eb8T6
XgIqi3VYJ4FRVqWEiNU1WV+3LpQIRhHF99dl40eRkaGoaWJS0XBxtWNgrSLO8pmm
oVEfeywHpltLxWgdfsuyKNrnnNMSeuDkb4ua9wTlCikE6nbJoQ/voPy5d2vEyiSH
XMihOaiZlX93+Ex0Z+Xn8UvZhmPeOJr4OnMKWSwzzC+Vg5aGSsD6QC01ixqKRY8F
+M54J+SlgdbinqFXwtnjYKhjivOvRUl9NPjrLLsDCZmZOahcLVZKS6GNkicEkXcO
A6r9N+Bl0HNDHA5Rxx/cfDT4WGaK8rLN/qDo1r3s43Szm7LWvP3bRouNcfMEuiqu
Jfb17acytb1wniqn8ck6H2p5KFCmsMdICX6MqiQHnABy+uy7Kk1E5npOssXZYM4y
kZ58DXKeyKM0B31HeCbAGBfW9wz5veSDy49wr6Zk4WzZ5HwleBlwdSO69nigbcW9
7wo0rz1sVVVE3s+L5TEt0VQZ2sfneEgAHn6HqdtThcm8r17trRklxWD5yf9tR/B7
CevO0reOi6qcarpPFAkiEFJtW3jYnU9G5Y4vVcbpDUo/elk/R4VrZR0VVqNbtj2e
LeyNblkqWozUDSFO92baGWu3Z12iRZ332sSKM39wAxt+eB8D7bei2pQycu620Z2T
J74XGhqLLALJSVxQtqDpwJL8GY/WqMLBLIchEAlWv1paPCesepQEfbHo5w1QCoTP
l3lfCgHSlJjc31MpNbyHfLZ3/hFB84RDiQppasDGPNkxhSE2T1SC3RpmUg7/ZAjl
PGdkDSQdl9KX8DKYX1dD4DsOuLzRWG+WyZwWcQo6bNuzUnU12iAUpXTmKCXGqDkF
bayvTY3zeetqvutELxb0BMgUYnQer7d4nWSvMd0tSyKPR5L2Symnap+N+UaApr6P
1mZwiU6zG4uQ60utVxvTDerWCxd6nJruOewsXHObtUs8Pvcq9SYz3cd22B92kNoY
yn59KwWpSrZdQNEOEv7AHRv59ytO/6oJqv8ubfpM6P4=
`pragma protect end_protected
