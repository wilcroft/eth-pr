// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:13 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ms7plhXZGWGEptOkYodfV8i3mesFL6T5o55WScLp6nngimVENVlx1k474OvBOf22
Fwx/TlMJdIF98HTvdVax+dwHbte0r96PtBommZZLx4B6GWPlKYX3sjtgK2o9wG3V
wguriVZpx+i3ghOVVOvZBW0aKfta5Q9WcrrNjgZNOIo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 183296)
64MsrHg/jUYA6aGAWOKIJvzCAm8p/PY9kxCEjcB+/jL8hEW+UkUUDV3jZgoGJXDs
xRuDhpy8EbtQc5Nk1MF27qm+805W1oVSHQNW9QXvvX3cMKxMA5yb7EKt00EBUFAl
vn7i/F/u+hjjIGs58eC2t4q9h6JUTSuO9HDPMNPyYIowryZBpB+yRpoiknwE07Yy
l9y07fpC0lHLp4vyRkh6KhLUAyNAGXxn9BY/wwIjBwW8mh54cFEPEdCd9OXTN8Gz
06RskrGSWTjZpIj8Fe+i/23RbJ2/HhZBhVtr7aeZmU5hAYen22rPuABG6gr1V6Xf
Pq9gAobQr7sNXb4TBnnK5XV18Kv2FRjR4yhkhOkdQBy5CSpH5N0ktqtFDd4yvQvt
m19WU7DeA6gdn9BhLjymKrAEvJsbwZprh0k14Li/LWO5F/d7MWbFOxKl8p4Lv7wv
j3lI95lVgA1XUe5imJXcn24ypuWhyxhU125M9J7jgAAp9MzykvliVSwTPNGwmOGa
Ic416DSheubymSTsLGZREsJ4WxJzR2Gjg/rWzdcKrm4nGWg/kdm2HZxlxf4tZJai
RT/LCbODfcjrlF203jaYuSlsaMN5v8nvJz//9ikEXIlbQYCHFoj/Mzvy6/tXAteW
wlDtmuMFm+98iPmehxFVeQbgQ6x3vwfsCjhlNJsNQbqmwVcjutEc1yHEQPS1/hOM
cTnhey/CPAgfmbXmC6X/LHtjTplRkmwqwteB7giiclQC100yD0JxC+qNK+C1/rPw
0b8AWOMK0FfB/QeoigIOZjq3qeRmIrxw+thQvYKmedO0LxKlQG2Bbd6YntowexKG
509fl+ivOVYrwfZ1QlOGKrM68cy6csJTILVLOYIUq3QEzBF4o8JU5YsGoja1oZHl
kJo+32hBWDD7Bwh+qacldUEmtveRBu6cDL1cYsg7UOnlLqbzXp/LLfgsp97JBWbk
681ZOaZi9DzUFRHw0mn50ZP9UkbAfsKnONHUr6fVxNjR9yRHe3+lRlpFm0h4nGv/
C2MP+u7SdtwuOlG23cKGBX6AqM6+IgJMMjXAlIMa+W+gLwYFXcm+59qY7YFNIB4j
MGyyiVqJu5QxV1LzTqMP5vwbnZmYl7aUc1ae1ggOik+mgva/gurbrry1+nTBhvNe
c+LljoipFdrny4h/wv9NjctYAXWxthni0GLH5zHcJdOGngejr6SmdKclyjlfCqXm
mRPhM9CL4B+bOwBBqV5lLfkw7L83nwmcE2KlR4HRS0YWWwG+ceUU0d/U2D87/TAX
xPSG2axQkPrMUxYLP2UP3PWCY1s87oS5C/1bFW9WdVETnrq2fG6/3tkDq5y0PU15
FQt5Uetu/z2PMFPNnv0+DpFmRf19yvZKbdgS0wwuD9YMTc9eua4zx1u5pHe9kc76
VGKgB/xUgPxoKX9JHjeZHz7isxIghocxGep5uEnrqaKCYX+N52VmXDggG2qiWBy1
iBLgkHWM5T6vS2mcvD4jC73BsohqwJQ9/eryaB7TZPrT0lM/RdowVYn2kxF5pa6r
cPI0lIFRXa3DZySDeF0i0b+8SEsbKRQ8arxNug8yidy4XOWWDFSywUTUwW8MQLSi
HnCLhvzXkNSIPlOxMEh1qg95bJRNvq5sPk/k6iqm8YmYnzeDO4Om94o061W7l3nj
ulfRUyonLXev7y/h3qb8dOeJ7TbplYMPqKbqtLRy0rB2/xRWRqrRFOUA2s4yvuAx
upZjaSLwNVdzD6uU2Ml00Zz0hl0YRP3troG0gvAudoXo81E47lQ7/YySoPTXPd4I
clqXZF+X8RmqZgzznsR+ouKDAa9HT9QsM4V6ADzRO4vDm5UAzFsW29xDgeZp5HvF
EmYeLAy80ZvODCIdqxQ0pF/uIXK+ibN0JjGUP4cXKGSLPnR1c8oGInMOcXHxenqw
z51Zxn1lJaejxDbtnIESUFVdH2NGsNcT4O6jRRlqpU+TS9rLbIbYvgJ6o9PMdhpy
xtHkHJfQiZZ7hn2tJv9bJqZIg6WgG6kuzWFgLzeEOH0SbnB2I/2Qi6h4ag/CZ5cK
uRVEJ97+mnil+9SqPtvjV4indhpEFDoRFuTmiOszRHoCkvvnsy/3ZgX9wQIJGE5x
akMeblm9kKu9jdG90mgehXMhbSeETHQPi3jUbK58R03U31dAniLPj/gmhjORImqw
wM5AjqII4WC8l6OO0Z3NqL8FUQDe1bO0oEExXJaH6wOGW0KmRuJZlrJ6F/h8Fte+
z3c/zlb+VXcPIS3xu+9niOtoWW/plw8asn9GtqAFswmuSqAWEIKFQh9rWdOwLdWR
MqcfOYZsHCH8gTHFo0fw83b0DIgxEszPv1Y60u6+fmUFqS2nQEkMyCHBCfAyU3d7
ry0Vx8EuooSWYsQ0jSiiFpOhyfWW29SEBj/j7eXmpfc4gXYsL/U/NcXIlJQ8NF1m
pwcWAcEHhLsqHQy8ZlsShqdfrzKvLu2GxZ6IIL9jFvbeyulehQv4S/hDEqeV5b84
Sz2W5PIRIJxkq0AY175dxgUMH2n8zTqBkYvBhD+Zpvl5ZxCJWva8d4w3xoxVponK
eIykFyEzq0LW4r9JfWV1SL03/bd+NwiA0DZStlsqrN3KHdQPN2EyjP5g++S+17vv
kUhtMX7+znq0TPsvSWuhHJop5p3FcV3XrVf2eCceLHbZXf5QgBC0ABNJ40OnUxiu
yzuUpry6QORIwKwhYYWEl30YW4uv10u3ejNbYjqN1wsn5gzb8Bc3VznTmeCkjW+v
xMbXf8pSRH3XydCtaJlzMYmLCh3guHlc8Z5TaxejbAZY+22sxBGFz8iYT8lNvOvt
mzSEPJ5hvbI1ZEmo44FY0EVZuA1LJyXmZMgyrENdmQlQ125M8AH7eL9mS0BsiDd3
geehCQsx61Q4bfpxa+xpgf6v8/uu9Kqh/uxu0SNBMQKCEbB2icHGFmw5NdH326ef
hK9IfvFUfNwcSe4ByUMyJaEFkmuBHxsVbb+PHckfBmohyVcWnfBqiTIoN6BAbA5e
sQR4z39Skrfa9XDpJ4UusP0c4iVoHI7En9bnaJVAZI5wGJ9IOoZh55HofIrq0Gd/
6X6tTGrMppWDYDmyUmPIc36TmpmbSMNNJoq1SGIvIw/48b3mFqSA/lrfhZAtSGI2
14I76XxyRvyVWoq7EmjnYnkGPU/8jB2pPapjoNLKiJFcfJ8wGdEzmSzBdQ6kYq61
vRAhqMbhStxO1Jjn9z2iotIgyCWov8OZsADn0cnA/pBWuKy7IRT+Y+RUQoFI0L7A
UiFg1Ap3lb6McRh46gPPzZ0NwZUzpGfxepjVyLkLi9z8RHm0wO61P5zI6Lw0s/9O
Wuu9w1JbQQw94DXq5bUTS9OW/RYlxhXdQ68w2GjttC6vukdf9xPuGjOF29byDzpZ
fGmKbD4knZG6+lfQZUB88xA6GNcdbmFoA0EWgQ2QoTDBvS/MrixMKV4kI3/KW8RE
FX5xUFkTyX8ZeeLlDkKK7ktgknYv4wKUv0gpktGTHbg6VoSQi8c1TgaAypDY/ski
OiaOhEMdZ/lBhZZykc1Q4WRq/1SdgzIPqxQBuCD70rmzSVoPfK0JcxgdF/KmdEPI
F56wJ89R0ppFzJf60Z3xJ2lIMWSg9Wn6MaNggAA/5FCoI9SU8zfYKCz9F52d05GI
AinUX22X5vjYnMTF+76RgXoSWArBYWj/dbItr6aajmDbyHJxY/vRshbFrFlWS2Z5
viDehLUJ8TgPY8gJMXQxhelzNEBUsPJXiA1nco88hW99OQXX8xar/wui3dE0mCzs
iyAAsIz8AURkQbQpvWfHz+nImCUw/kMGLCZVFvorDT1XRLohJxFdZMrhz1/BDhRD
cln6sRYWwuifD0Wd2NcoHkV5krktqpmGy0j52+VwJ2hZbU8DAbQD9uylDcuLtpuM
O+56XCccbY0bRaBDrpP5LLHUFQM2fVHsVif/Sn7LpAzaXDNIi15RpHYdsnxybm6J
pRdNHE0LgvdP6j2EWpefj9TC44cIxn7Ax8606j8wtb6bLc+L0/d0eRMC0PrUhMXX
N4gcbi8um/sZWqt72RLbw7JlzeKbj7lFRGwVIB5VPrcJUVw789Xf1LUskfypVu0L
ohIIuYkuhObKbN3nOKNSDHN6ak+Oc1SHDQCjEAGxy7kPHdKWvAEyyEjPZwl8hoAg
Pbkg2y/gcuq2705f0eUH0gKLElS0wzdnjux8pFacjNZbgypfz4NUtUbu3nNy0Vic
Y/2WGMqf3iC5f96KXYO2DxFZ1/r1T0hnAb0BaGacaq056CO/HZaHXT6e2vx1R4gA
XcOp29kJ8wtXjZgRaKpHqSydCkSdGDfAs9bCCtNcTvd5IKSnc7mzspidKCJRLaMD
s/zlj04d2Yu6/SYo3QEl2fCam89ZhFLn6anFhpqq1muV2B6MDJB5Bf/YpWU/4nLz
TNWoQL5IyThNglZ5EFx8lBZg/ymfxMJC8ITw3UWif8qGrFTjEi3V8lOMWWbvlQmg
xIfnqmqi2bv9Y/hFIBE0EvBEiMbLNr2oWmg1KzEscHwdGqhDS4rwwmNUJu1K3cuz
hVRecP4Pg7+Eywumftn4dQQWJIFMTs0rnLujcE+l8GAtFMBa2XBSyh0D7DOrRRWT
Ae6bYJ66zU0hEMW86A8/DVj2sviQhIh0ZtD/7c1e7tkTdIatQzr9QZvqczfPd+8q
01rJGO9Azin13+jm9Vl3r7/ig3cJuTcgC65irOev3UZxtpNQwl7SQ1s8k6E7BsVa
rLVjYeKB7IEVm5wsD1V9xJznZBaN+DRNmyEdb1R4kWCo0nssYP1txIjewGQ+dSsk
/mhwVsG1FnpAnngZoiETf9fKPHCkXV4bLRDXjRqg52JqWYaJwDy12MyZo07hDefD
PmFlCSVrzKE/+2UNCfva1ZnlGxG1D3wWdKC2SuPTY32EiRLFfiuAR/QSpwlpWBfk
SVN9XTlkVWnMaMUoTbqk0mnPuOTEBZiWgoB4ui5vRsun8NtHIkCaKhmDMjYduAZc
pul1flZXZFCA4ksduj8RFVuRDmsdrvjZjBMI6KhtqiyBqEoDkwwV4w4/90onEKRv
9vzYIYObNkIV7SWCzP41+UKau5A4cEhCqNc63IYDOpakY+l9gSg8ZBao/caqU95p
+LJRowfAs41hnrv++V3/rLcip8zwiwRqPcHxxqjkR3/ZFIp7W/+xDJth7o9x0OSt
jlYlhwDeBGb0IfqyiXYE1QJtqvPyJ6/wvkQut5g1wxF0fopeo3T4FhkozjBPtKvD
1iD25XnHUsKDJya9EbT8CK+OP6mAixK+qr8am6r105A6XgZPv99s8nPBfmoTZi9J
sCeZTOJk7rf1Gk6fTjFfGqHEqjPiqMrpNjeS+cOaomji1dnU+NakScyZe3ST4xEL
FZzYgX4D5omY0mh/3nTsF5X/dN1ANvvfrPIJkAQiChIMriys04mArKfomqHPjbjb
qVbzwx2LSi6aCu0MHtrqUTfcqHjCAe09U0H94F5QZ4b3o8Y+jTnXnoGVp7DQjAfB
N10cV/DTvAxDQFTaioXKQpBCkdcX+q8eo4RZBJ/G9yH688rtZLIs8VVashgzdTfe
pva9oAOtVtzZCgow74dqzVtItcgVUBwB1ZyXEtnbBxnA+3np9c5b8EJSSWueAPmu
Tp54SKuw5/DT+Ws2Azs32+e8m7z9Va8fUWmmiDWG4DlxwyRI26c6JvcybUALHRGT
0ikGnO4ufkFpjDAsyiR+/elqOGZ0JalqPkpa4yjj+j9/AUrR159TyzCmKluQRuHj
G5Xb4tGREQdNQ15ThTsGmgZVIEReJSmJ1XCg93spwPCDvEveMGH8P16nnxRjjEAh
sRL2/TTaWl8Qc9JmpQ6O3Qr4L40cTz3b0KOmEWO42RNMte87VV9d8tSWeqEptlgk
5jKc/Ed4ztE2sLeC/RGEZSNeo/r0C1JG0XDkxRfC5Ae1AOfp1Wx/K4kCWM0bg0pQ
O7UivaLJSCt1ndU6gQXDV/O3HM/NJ+uDvmoxWEU60FHoHgd+qrW3MuVMPLxZ754/
Hi+ssIK6PUA3BvPtUvkygNYQ7UimJMsLxk/DgpbVUVVOrznuDXDYDRfzLd+z4IKi
07he8F7BXg2hg9EtLVyeZ+CpcQYz9gBbjR79krUuS3kCzGcFi+6xjwdEae+3I0b2
5OiBd9z4TeP9iKleg5P3Vqe0yvPMA9s3RFyMo4ZYG7WlyUC/8jAtlyypwMqIacvU
iPf+xGP+ic8eG1ZzlsdIXvo4Pjv4HEQd5lPO0n5HQ8mwAjN0LIlPZoS04Y8KMBYa
NeWG2oXjc6jvYY38sX73FdPWSkftEp4lrfFA8CAtAeHnUun+ZEfcJBrYdMXU3Wxe
7QXxgpGPdiV4pLIDuffr6taqR+Q6wYujEbWG8Yjrj7GgNWs/FRSSOuWdXvQm/K4K
2eJbcR5ouinEn6w/0mpF/S06fGsPFgtZE1HFVhDh7hAyTPJFaF3rpZsW3Uqb8xlT
vCm5GIMmNC9zjUcudAxqlvwfXETKf7w1oMVr7L5cB4/kt0FbFjdtRvsOdWU1rNGB
k5ECNCmCnxsm1UIfwiHX5VuzcDkrLId2McBLA7NW4KouoAbk0sEJtzAWYOgNiWRK
SgfaY5EkXWGa69oMdDdFnKZL7DtntUCFU3PHy4FNlPVyuMZBBAMgAcyXmnBk+QRz
HiPDFMRiZqmDJ/zqyrPzYQmEl1p33cH9nnhD7RitZg4hWouuQ+KetsyiwK9ZQIPG
vPFpZNZ1wPCB84xLMHfREP06F22Htjh0HhstRaQRnWrqwyLmr5rjWaFKMkueSYRc
1KZeP5EBWyyr+s+c0ArLaHLIeIKCowH1yF2QLIRcn/HqHo5Nxu1CVy/anPiHNDnT
p+TFqeIIsZUrJqm77xg9v1KOG4PkAD8/p0T2LnTUi2M+NhoM8J7u3vkNHUNLUl/y
eQdWgAxjoY5VIeFEburt0Lk3Gvz+QKjHwx1VhrllVbl8M1nqgEEjPKPaNdCV1Shi
gsCIT74A4XqJcg31ODpNEVvCyiGHPtqmQA2/kcs2+ts4/jeUnDzuy4tRiEy8/Ubf
ZzCoadkYG53JfL5vRuG3Jlw+6wfti3u9on1aiSwRVI4pEhQslOtU29capXcC+TlT
I2Exaw1zM8jNqYI0ifhZdBNhnQkWUGruenz20NTJzFb3fj0tTwHNseM0LPptwE+g
3RG0otyo4ZbZbXN/qGPeDRHUCH36YtukF7+s9Zqihq+PWnePSb+1St2FWVFDs8Nt
sHuu5b8//SaZso4iQsR0rDTb+dAn1p+/QeEC8NS0+/2aMEKSje+c7YHDF03yqok8
vcNgA1mBnaVXPVRETYmd5vvrbHvAMXyp6/q7rDrwSBwYRuz42BzZag8QSrfIuDfN
J9P0QG3lYnfOagvjOnXmd88NNqY45b0hO1pzssEC0FvWWOMlem7Y9MTAlUfT4wLb
a5+ozDupcpLrHy/sqQ9ZUi+mI+GZFEzy0EeW3KEIfc9XQsL3Z6m4Yum9YeiyrBbP
4BpEDRGsQ0QKNAMP63ufwitqqpFT9wOenNxDLBxHNWxgRDe0AOHRNw8l13MkD65w
7pdNhhqGK3WUblW0v9O8t4um8gz4NY8bahAw2euQe4ocx5k8aH+rUeK/m4+eAnpN
Rhj+gRZeYkFGcAEm1JTaXqcuT/uMo8RQcNb7D1duRhAEYcJyuwWqXK8iNtpdwtDw
QTNBt4H5AEk+kkp/pPw1ZMNQJ0A3NcR0SPP2ODzyJnDo9MiPxq1onj4MOAyxudNo
E/CPaewgYTq1xg6yVOk6iRBC2Tjc2Mlj0dOfWup8Cdem9TVANRXjnIB0K/LPaBeB
zLdrt1ZRSRRf8kBw1PhrAWhSUyFucR8BtT7mWB4pa3/kN+m+I7ZbQdOJg9wDsZxn
A9TN5LdvXypK1NX8+iF+bUwZ1HiYuI4jaiK15Oy8ARzyp9ZoZjFhn6j36ho7ZPDm
OYJdpdxfvJWBdVTx98HuMlwoMjDUsYbvHBsqyQIx9nV98qZ3/ZTh8ZCMoBG+fsFm
kAoifgBrtoUrea3AXQPfN9XwUq3Zd28OaF5U/aT40eNi7NkyhvFOpwq5CLypoVMm
i2wkT7CmWACro51SrHm02z3dyQWxuSUqhcEUaqDIn0RVTshWt7smAj1hIIfalkGh
dDokIQh9ErLIaaiXQelpLhrmaRLbaCz9gW9f24SUDHkRXfRfd065GRTQWLeaBupG
eFTn0+ppH7bNb6rEDDszquz3lyS3MYgtDY3YWootW1eup2keLOtngpnFS6OJh+t8
j520/Wpdq+8Q8f7XzFhJw/y3ZQRKgMID9opl6mBcVozgywo3eDFpiLBqDKOPev2V
L47kCUA5WNjyspL9qiVcgEPYvHObtrKBKrYLhWFRjEBkGRXCo0/GBWTyolfA1xhK
79C+JBgxo2uCY3RyaO1aEV6wJo9tTyM8G+z5FXkluD5rtovzot0uZeRPC5E009U+
A+1yTSPx1gBnGwu+wNP1YnvxNzpHB2mNzABu+sOZS1LaJM2sHV0sVUPlHOLidacg
B1/imEtSECkp84/w8d2Za8ETo71Om60DaN1qnLnwPF/Lo/3zNJ6ohuM9B4j2ume8
E0AVZfoGQZSSNSrDKqhzs+hrR2ILCNHBQGKIRzEz7N2ci0hfahKXi/3quroD8WoB
BfQV5PjXsWw9+7GdP28ylXRUs7/vI2btckWkYYcYrRosYf3cxsyLkGDn8y6HMQU9
Pk3NPC6xmQQ3hdWedp1cRhuTO7N3BV/94XuIiW6DLm6zYhT/qBUuKoLIhSz9A6Sh
HBAqe5h0DE3CXPvZGpoKFTt39arW6OvAtK39avLUIA8BRDuXwRTu9ro6LG2aY+hg
p+4RkUx6Wpk39yeMauysyxngTgybeFnuBQaezNPsBs0QHm2GWPuo9f12vGKvMcEF
ddFNf98FTotLbBaSRWs1idONr3NofDdauL1Bru0bnEqneDntESazNxivN8bz1/wA
TFXz6Tu2o6KOyvGB0jrhK+2IAa8ee6TnW3RHbsx//Fvu3YGqEpE8E7j7SWfwwYQ0
z/wNFQUxCy4g/1I02X25lg65q1G4SYi5YgvSSm7obzLLWolprRDdfpPsEK/mW0mh
TfSJadUUGfZviAZknqQP5PiNA2E+/kmRjbGQduvVWH6uFQUedbb+TiqtaFQAKMAX
QL7E5n0HMeJQsavOnmBuRu6bgEQ5ZGY31OWxIh+7ft3cZzHrjPMGFOO2R5ndf6DT
YuESz5mWyeOd/DOcI0AAe9peRjKjt5EHyYFC370HPoCiMaUASTFH1czk4KFivzN7
yqDrGlJnLSQUqFS64LiuLnVKfzbKaVm+/+RUdgQ+ruw+sbYC5KwUUAyvpmBMv20M
C6XAOQBZygY4hV767I8nL2aXvUaGpqFMXt0xxXp5TByLs19DDi+soOudyJ7tZ5Ks
UBsHpjkfn2zajQVPGlP19KyzknDzNKaGtjKtEqqn1Wqryab/mAaQPJ88luzQSLLJ
UjFrLICekrSZ7KXqo5ikjM5mk+n7XMM2feN4VO7Hk8PnZf/infGzfOv04d0W7CAp
5meBaNoZmcUaT1zFGaY3FR+/GNV864RYGyFl/61o95XX6/pL60DkO8fyy9FLRQVE
7dZ09eBkh4Ze9eLbCYGX0fpczAHvAD44DIA3tDB4r7n+h0buatdQI02Fz7qH/3ju
WZ/caJqayLMx888INuacZKrN8BYtj/tENvGN4DSGJZiyPvUQaqwhLvNl4cITlPNv
HKUJhrv0vwK2qAkJDqrPvQxDOrCp5qoLv5oJekzxWvs4Rlvjts6+H5ZZdGu66vqA
z4KswfQI/qdKwV4LGrqn88UVj3aqPH+wO3XTvqDNpetwxEDHBp6oednOsCiAauYa
OMvuL3qrerWRjF9O8csJftCBaw1+NWtMkU9ivyWjxPn1svp9MWPeiHrqFzt+q+XK
Y1NdqRi3eJfILRHFaF3VcCo00NI+Se4+Y3LHli/L9LEYAQ3Ln2286y+OWHIvk7wv
OV9Qgkbd8uyUMB6oPhmam/xjjtr8YQgJoTTy7puozV8rAmMWdFLsUN1VhA6IYnUO
kxybzoGTlJ20V3kZKcWtN0Uq8msXlXDEUPvDTlej/cUeMZZb9ljvwLTPfKfTdhAC
D1o4R7agf1P7Tx/0KjiyTeZ/Vx5YoeC0PRgehLAUYsOoj6QbYaICldc2S6xQobay
LTiwLOTY7LcoDT2M6cV5xbua+TlYftkSOerVSt3Sus+VsqrxCtdxxQiJB9HDnjln
5BS44XayggfePP0m7o+w2RA11LSUl9JJErD3yF7GB+hz8gHX5HeT4Vh9GCGJZ3Yz
NQv08C8ZzOwewBYAVVl+n1sJQrqzrp0c5O1QlS1YQjp4hy2arVs7+W5P9l0Gep/q
5vBEYVTtYs18nTzfLfbwcTsz6HEa4tHxEiwE9aVuHLu3kSWe67Es09wKyFE0jpr9
+zJ+uVW5SWH6NQ+wq4z7WsqKcByLGAN3o4nFEvWCJn6KStJ/EZc4Rx/q/6BeqSWO
q8oY8ywpFjF0CNMCrXBoWcWv7yI61TfgWcrDgjI5M2PNEL40qr0OfAZFocqbKmlV
4apyaJRAq8JCsfI9bTI9XsoDU5Pyuk8fYpmbA8CNKG6whKunay6i2WcHWu0rDeyS
IZ0mF2R9mab7YkpZv/s8Xip0kc4ElyuSVlvdI9QLscBkLA4t94gV+LYyoOKDz+fF
R4AczMCLCf9JXUnkS03h3XtSS8CRA1xkM5P6/rCb6dcZs6z4aI7RaWWZiltcW/fP
siE5AiLsP9JOqcKbjcbETtCbfsXvlnMdFSIngQz4NG+FyArtBvD9eP2KWgUXbMS7
V6XiBHnDLxVOBQcc2cTbxAVO42h4c6eP/vYmv7mF5aUPjpBqoTzLzRPy1iPPmvWu
T6AiMras77EuuAEMsb6LGZ1i70UxfM9Hk9QPCFxV3S9ZGs/roa1p14OYNE49Flo0
xtyHU46rvtLcoBnQffCMnuvnPWR+l4vm9SlJ6dBOFYpccOneBfkj3zF8gOUh6lOe
olSr6YUFQkNg4KxA+LfI4BqpJJRnqtrpD6wuDLTNDdpDWwnZqa8C7w+wUQK5JusM
pDV7RWHwrFbj6ZflnhKqUpb4cWoVfzpG/RDOUwkDk3otzfikeiIb4MKOholRbHbR
cOBOIbWuX3lfVNdYG62UKI9o0wyMhDZSQFiqCEYxx62RyLRm3/FHKNoVjQTF/QtR
aOowuwT4nsvfwDEAgvChd6llOxGKUh1eI7Nxwud4ZX/9wc0O2wSv8Zps1TYg7Bid
8fh7zESE/FvrmyPx0TKl9Kdw/jFAN/HPOcxGSo0Y2ZsAhG41slRnRstOY8DHfLs2
1GrQeUVxAWgglC84ZJ7uyOcrgThyw3dC2NTOGcHZpFaRzmvZLk6WaeRC1mHo84k9
FDB2489VNxK0Tlvcf/R+NKUqIw1VWs08+OYhJYJTYfEPJ2KNiJ99go6RquQU13Qo
1KTXKR9gmhXnFkY7YFjkFyEF3g4FckP/4X/1yBDC6CoedhVGY/cBjn/Yr/NuvU9m
v9d8hOLgF2PflvcLTNLUhNaaRNg6SUFpDvW9ievLNUX2IYLMxWr7+5Cn11nGqenD
LkeH/jlJ36ne3TnDwbqm5DHn8FJ2woahBAUelYY7YU7u1sKA2jS6HxC/j9NKM6S5
8lpPCgKmyYUNqQbE+NugHsMWdZ0+b1JPqE2wNxUL4ON4Dt1KK9kjGggOQZu43xy/
U9ZOhyEZsGaSnOTMITi1f2UdgJ2GBdVUAFyO2K4AEQ3Tl7Zc390psWcZPI/KzJQJ
GCT04Fgh9neKsJTyb3vllgrbLl0mPbpU8+Di8cQvmwtBGe/ysh16e2WQ1+qlSgIp
53tEqZak4ByW+ThrKr3RNrnTYHVXnzUeDPDTi/9nABvLCKFEJ1zM8tGpMZUl8DzI
uCZ0MuY9IsmXhjoRDBJ/d15ixgjn6FpcLW0AeYaYM+r9pnWVxVq3eaWlx1SycoTg
T2jmvHUTtGwOnjxq+xp22x4vuJd8kjmwp6zW5gZ0WpkVFuSMrdKCBei49bdm53WH
aXDClvSB1SefzCV4ZvQA+5846BngHRX3n1GKEZAqE19N1daGOxsBiiP2P/OJnr4r
w3bjpWxcSWfrXdEm2fNKz356QXTrrcxpWSSM7KkDCgzSPW4Il+0pQTXClC9/rvNk
IMo2FA0Ai706fEmq47vQB/gDqgePzwgW82PFgPJBq/pkJtD6KolkAfE1ftMgXPqn
KFaCBBub717kfCODWN9iKgJGepJBSe79KZmCIf2VNygls+ZNg8c97R4dmmH/yc9T
/ljEmYMAgoCkk70wQfMnpmC6tIFNkXo0Q9FSZRn7b4WNqBsZ08EaaNdXzDgrTrjx
fytRBPA6hVtSEFcd3u+OSeGFd5tQU2OfRMVwCpAMKNR5rCRuJaEVO6qcZkSewnoP
Mrl9Zwg+91Z+ULBX//9/G6rOvxqss+wrw6HSXlJOBBFXzVK57GDUdzilnmSo8FjW
VrIWPnRVQoCiWqoggF1HoZFwl0tvVydUW13NIkPx36Xskh1tUSH6tvrghc+mZNzI
aUiaWMoA2Mttaf8n0oteQ9ruODHxeDxwW+xPaqrAYq9r8VwYQvv3wCwr1SvYf08Z
/kWLy1oc0uf+t6ccSx+V9PZz1YNWn8tDySgHBY2rHtGP8w1gs1YEHQJbe+m+gcFc
fpZrMO5gzqGXUFdbD0U1dxy4BG14Uta/Efu1qeAgBzosfwXzRYaZng3CWaPrYeay
NaHKuDN63vePuh1IBR4JHBQrxuKuv/eYr9Bqoah6+npMP5C+y1VC0f1jhsV6GUOq
wSWnarxonoCudYaWS5QLMoFQI89ezlLMEgfhXq8AJFofSnDJsKHHyEwqQWVaGF1m
1PJ+jIC2tEtn5cB1i2VaRV8QP8LupPLQgs2pBnCndRlhM8r3KUt37bxulrGv+lAE
DVUYHOLqgJIllY5qK6aa748FQ9b2oBuEsfBHZ6h7frlQejl6WX0SKbX6yj2qjvzZ
C1fUqwTfTEUWBwNA6OOqHE9uNXoyGTmL46KFv0PQ+yaYmexEl9ZLlCqE+U8gOB2T
tzRbitVjypb0UaeJg6qFohG0wkrMhIcJVqlA2NBwvRr8Vif8ikGrPqRwil6YLzeb
tgpBlAH6rby+FfMsF7tXLxUF6wDraeFw030g5OoqmiE8fmihHViyfgdCaIdcicxp
yFw9hybycb4+Ms9VvUfzkVvIdkeXPjI/em7z6pUld0/VWWhSECuOzufxo9pdNMkc
0aCqD/yfjv8Og4P2stREjSkMUVgQKdN8W+gKq2NQKfVSJWSyrWpDaZ6QTQsaXxYE
JcjMVyc1KceLYPDpAyCBvzdoQnalbegqy4NmS3n/WO3RMkvAOhV9AQ26IqpQp+yJ
Fyi6DHqioUcLW7CiuBRMdHSkkwmZOQne27ul5ZG5AEC3gxjbCA5KtZH/uq96kJkE
r7SFPTg4z5nRLJOLkdexfD/isWaA5vG8MH4ZOOr2aN0jcAQkjSK5UCLg2/HSDo6W
aSDsm0UknBcF2sBnetYtALpkUUQg9XXrlOEg7uHprypbTtmXhO8a5r43mHDMcHAs
1/WiPcln8xh741DPyjLxqrR1fPn+W3UIBfnCn6h2z+OLEGVuLrn0HT34mNfdHhTG
hgQP8g9EbiNDoepXm3UyW51S4ERkSKmUXXgsouCIr69tUo20GLWjGMwurxuz43/w
E1eVWJyVQm0sdbLldW6CO0ZeXlfy38EWZuI1mOW6OebWFfsC1swW9lseNeVBHl7o
jD+SFEXlEpzA5c3ao40ES24Ehu6WeyRyM3c6g+b156cOKtKdE25bweBjNj/eTWpR
244HR9W4AxwEAwPVY10wMtg7fHs8Gz2kNGZzgCK+O5mP3csN/d1oYD41x29T7Uyf
kfsbRu2XsXtURTGF9fV8yIEX8erIFAC/ChG8IXyU/TzMDSmlSxa/SAD+e2KirSX2
7b4XnOAo3hX/KwZPT1mn2+lL4ItAhTpkOrOcqmY3TYmGm3QzYlXgEu/582faZD+c
/L+K5DHLmCWQbChCbhc2club7Z8I4MC49JpAemFOLNL0FkLhH+D9y7jtpIk6e5cq
+9LOITbC50LgAmpMbogxh2BapZ3esXwtUzzGDc0tG2lmyCxQkUDLp5e5m3Ond98v
iXM8HRr4C5iIMIjAcUw2EY5k+RXRxbdWiHu9WBYudQkb92HekF6pOWmD44GkwPMk
2FSpZlbFlXThEWVLaE1Si7u1sl09PymlpiquudjXdWT2q0wMcIdF3WOiJRfkgzl7
tafF+PLpJxrvDM+TkwwyIx+9aTD3IXCmI16IMFu3z7WpzdzuVS0UUw5Ou7b0r5aP
v3wTdkiY9HGIPpug+F4MlJ1QZ21uZUY60wBhFV2PObaEhruoR39FTk8dBZ/NKdS7
HXQpEmqI89EgOpbv5HlyFSySD1AuRCzHR8nT1mcz6lFRDrrKdET52O4YPiQc6KtE
RsCZGeLqJzFj5B8I0pnQM3vrvOj+sV/x3KKvU/bWMMXpgYnB0n2jUFEfQxME234f
QVhcK1md6Gc9B8fP7XQn8jrV83SCeXSngorbtHC72xHSCjV1JQYyxYM8OVnTDoNR
dNuCMD+pXywMD5IWGdZ8BOfIZOIqB9iLKcRJdkLmHd14r2ITSFSUyFu2eASCwQR5
zfXfPtJHCzeVrM82jcj2JPWAnTZzcN7Ct+ZZ4Ezekf+gxAUrgYfInUHSbbSIIhU3
csd+g9hdwgVIyPZxJq8r5DBlXuE6qotc8/Ie24MlJQgSMejVpljjV7z3V6elxd10
7sL6sHFEf0M6uSl+s16plsiN5/LTPeIsb6pEmlcxUl0PqbWVXOgsnyoWU4yEQYxa
NTzIvpVM7oEJce0oHWP+JR7TU54n0pegrk0Im5+HNQ2jFw30666xuL1+ArTpUN/6
l8XWqfWJWEZNR43perOu4lpMEdyE0SnTE7KOeh0xAIR/dVI2UaVyUdeTsgBYfmyw
umxtBvXDKHyf86YhJwh7bXjeeqtm2wSlr7kInrMGYDuvR0GpSy/S0/OFiLrSSux/
mkot2v/LkQWzISGuxZFJSaJPe8JHSgh6yNNF/o63S3i+6hnYMGxhQvjsfcNtIxu8
LgWJylycPEp2UP5FBZureI4nGgTqFtaS7EmLXQU9wTV9ixoIJHOumpGt4RKX2vBY
t6WIcATt1XWjZAfKlb+5iSgd8XtBTUsIJlubgjBub4+KW6tYR/I53QcGIrvCJ7VZ
dF04YtxyjoPWk8M/3rOv8Yr44n4nq77pNnCbrMTLk8LaYCAA47bBV/++o57aQl13
OHeAJRSQ7hP2TyVQttI43xk8DK5kxFs3uA9gj6zgYibaTYkd7KibV/VZ0S4Ov5dK
pcUyGpAwiP0OGQdTVVbg7DPyheZQlab3q2pS7prUm6FasDoYhvnBF0DdFDw8qgQm
OfdX9ITG0mGzoAUxiRYy60LmMgyLV8IJk/4q/Z2iaMnxZ0quvF/0eF13MqwjCffY
thzX7Bxl69jWhH9Sz2c0ZheelrvMVTL0CnlqPbm3sxRE4SJVf6xwFWx0Oc+52Tsa
7LSncIawiehUnBMnXuPtCxxp6y0FHvJJrcuJqkW3V5xuTt+nBR9qPZZFhKBCDOJL
ZPl1hnHcIqlC1yCGnTnICEBmkD3ujc/7Nfkf0o9m5EB9j74mSD1aC+lLc4hb5Dj/
ZbgnI2B02Wcfw675KtdGdEbyrlaocxnDtxa7Rh80Aqf4s0eaOAFvXD/GP04PBsEB
RAbqXcC3rfxKqP/4juASFFjCmA84s0bAn6EpnlK7UEOzX3ESRN8W2oEo8ShGRuqe
u5IAAqQxImbQTkX3/nqOs9dWR7OyS1bm98TRlL5ACaO8LGeZiLRTnF7xPfpo+hpj
uoouwqnjNRMIPxT6I0ANgjdUep9tR4VSTqcdODl+ZJMxwXKRAehe2L8I+wKOJuFa
xRU2MXHBSiTMmkviy6EZheBsStO/V48lJSRwEljEX3z8TlJujG0UyEgY4rkPtCKc
Qcp7At8GMerRGh20hkf3VjLe9yrNuKZ15Yawsm+o1BUPyrfAOx+aZx0bX+kzzhAM
BkT8YXzHCF8yNKPHedXd07OJUlklSC89zAgirTx/IUyAaXX39KKq5IoijQV15n56
sFbGiz52KCBeCNuyaeN8nKuEPYCsIKCezpt1YzuVceEfUHX5HRofv5gJ7T7ml7wQ
FVXBm1WZyXFX5sCkmQOz+fyM9iFR+/tsqtZqLuSXJvo6fTEENwlMiXAA6GsycwgL
ZrAP3fzIgK7Yc0Ag24rFP3BBmg8Yew5GfcP85gVtJrpQYZJCmzztplgFT+OgpHqB
alEdHk1ui2JoJUi79meSmeRZjspUup1zgsYCG1CpSQcAkrSvVA/aILXvtZroVFSu
7ODD8ELNUXXkRhqJ0/l4YoeBmQpoKELa6OL9mdhUMtYSsCTdIj5+q09yTNMKP4y9
Ho6H1RBaJ2buqepOSWRRKwFJTT/WLcnLrYLAJTYoe2dvNqHLU4DV1Wk1Yvc7I1Du
fl42ZKA8IXQWUuc4d2YyupLbdq+junU2/s6+dNMg4ug/0baHVT0FKofGUZfB5V85
mKnGQuW/hOdgnuSbqxx+tT/HVCJ8ZNDnJq2L56ReKZS4KvTWuTlGDlnu0GQcmRqE
3iUOELt3tOTVfn/6AQIV3j4lWj2uKFybnpqgpAIs6gEybESlF2UjXJ/VXJMUQRJO
yuEQ9ej6w8sd3a7YXq/xAR8NgpYdlM2uQKKbRixbTqAYLK2ntdHLQ9GtOaSmULmj
UmQhu5aLOV0NcI9ETLg02fwliBvi7p6yUER4td9oRhAAVmNmo0Pu1hxJTgikmEN/
FphnJ09n9d6HBgNmiyZAUahgNFfVFtw9GQQgryF0bAx45/sZdOStNd1JOpFXel5s
L1XVWPqUYD/3nbKWqjLIGEyDfsjG9sX+Zw5xSNDphUyrkWTKwJBe2bIM+u6x2KZ6
F450X5sYSllklF//95U09a7wC1NKAWa+RbWBvZ4t2xNiFcaZtAwZWQXIRGiOt/Qp
cvxuZXthFf11wXeHBRMyAejB0eCv9DVAbcxAPEk5HWgq313uFh1ZMjhZgC/pt9cP
tvXkcbgnjS8zcMw5p6MXREi5hxCoQVgLKazewfvlCJn2/FHXPVb9MEGXjzjnArdV
bMc6b8FGT8F4puOkenmikOfVzlOQcJucbvSeO32ybR/rXhLB53nmaTZb/EZUZ3Ct
hkk85hzMKJvbmzJWMC+E72wTLiASlgooCAawWVroJQ8yvK9Hi/uD+CbXGJR8yGs6
joL/HSTQuNIGnXou2Znoffq5xa64B3MJMdRfN2cnxuaWZgr50H4GRJAbTiGuaerH
7um0N9ZfF1AELiZ91If5XcjoxL3vgEyvwJb5HJPp5viph8LZ32MbzaaLKhElf6YP
UsVLUCpy0eUbrRLJdoWwUpH7+GShRzHTO4Z7t7OJ83qEiu2RC8TvrOtijzRecpev
YDoghB1t1U0FbXr0QcHjmbCaDGTY0KQWJ4ODy4l6Ot7iHv6NeR4Db6+sySLFNg2I
md978yADwV+D9k1yrEZDLffeErpM/ytMGvrVQYvm0Yj02WSMUcSo62Xbxm2TgPV4
yS6MPsmtAmAyxbiSDrJGzOlmIVlXks3wQwckPDsxczv9V+aES16C1c6E6wlkwtA+
Lv2sHaUn6b1NsnPqpVrIAIeJw3jstAJDFNfJU04cx45ZzISi23RusRRRsou4f8dy
Uu6zjZoaA7y/NrTqcghdDh8AbgHy4TAqBnE+W60DI8ZqpFngtdGcf31dE9zdwpqP
OHNnL+7ZcB1MjpSfFfHqDN/7RGIGU3GzFxzYNb4rOt0WbLOi6UhvI+WInf1DOE2o
cPypfWhfbrunlqvYL81ZszGnTpiz5JvogxsNXRNdqKZCtTqPp8AckCwY8P0Fx5+f
dATftFb2aq31XJf2AdztKKrBhzRgDj24n7wngm1MYhQk7NAm+1kvOT1h28gbavpX
7f04KsYlURAPcuUTzgoaLEwU83nZ5z49+Z4nSONPheirDppTZz9DTxsD2hwG+Ons
Ni6/THc2O/Vvx0gccQNuyiw8bbWe4bTe2JFbbrA5B7zVypeP9fmjrxRVqjzDDaoZ
imvAahOs3js0JuJXJOdpPNJrOrAyHHMIZ6v4zZtdOHAPyyh6ZnbekwzlhsXVmiKN
eQDghnpM1Z8LOJ422iDbYdXhB0m/t0giezo5qfk1fD00m47CC+jSlhYP6IO6wfX3
nUx9ejpKZZ7zpLUYFFHUmIe2Mu/o1/y/8duu0P9d2pp4CYOP4P357IgqPTKYt51b
mi1Ej/aOtlbQUUmtNAMn/4T0INiTgCry5147ufmVOa+NfYtl8zHOJosK+AhBPzLz
gs7WtQ54ZhCZ8NoJJNpMKSyFT3SmPS7qKnxGYfI1uu2/DzUyH5ACmSPvvQgAm+75
dqPqNiXmLi+jTNW9ojYgw9hOsQnLhQXnZ9sEUO8YFBCuQlDHbBX1Ze5gVkbvmlwJ
Xr0QPj+Q6pAB9x42cr+LRwskkV0aoVmBNLJlVtijgshkarGqCIXKHh5UWkvWz2cZ
w/rnhl119uLHX2DJADN4B5LT9FLwYHnC9doB9Wx49cea/UOSg4VDjvi5al9SUpD5
2W0ZOPZf/A8G6m7hw+m5W5azw/iZFMYcyb7P9Jg91rGE+x4tnok5mIuTQXA3cYaD
wCM2vTczRlx00CeiN8mvlvRSz6NtvOlThkFp4vMQTzvyFQfWxmunQNdpTctQ/RSn
LJo/XoZmPAXVyXjG85p0VIK7wEhNgKPcXNVBxAX0xhjPpftVaDRVytBtbXl/9E/r
wM9gvr/THStTCGmvVvRfyON8ldn00j2Aexwd4Qf+3YJpDjCC6ySJM4ha6abySJms
eitVyQ7edEIimSN1xcOrC4IbSVzNe3T7SEWS0w9T9wg+eDArbLRNXigWABNuQPWS
5SympoLe5jo2bdYUgJwy4I8CPBOO6lpgy6EGCQMjFSlLBg27oWfXDhu4pJOgVEvy
g9s4igBkQAzpG4zSgMVvfgYPAiKL1H9+JolfJY3jw7FvfLQWO0bzixeAl1aDRBgo
Hqtzzq/Xg3Rh+nE1vCTT4kOCK7UsmrEqiEZWKfaxw4YVFL1L/+xjjts8pb2abDuc
/UKw8QyzxPWeWhU7Jrr68xhb3iW8OYK3Y2wI7O3gKTL9NddNttVx7KvWCnf969lO
gPlUM6/y2wvoaeCokJnjj/HhjMPWvDMDHwd00zSeYuLJjqU2yI1Ez8M/mqATzC7H
zQra7WczAjFgZUTId2vKMFswErnoiF8jhT18ZN6lv4+1nCsseDNV+ra/ejCTSD/4
9DCI6QpRNCRnh3j9MhtxLPi54vXoQJohKucTQ2/b0senVamGJHNheI0R/UCbAUeG
VLnlPYZie3h7/KvL1VlBB2VjQT460jtMT74c088/EfWOgjEvQz8CSsCsQKkqXlBP
A5JogJM7+bkBrWNo1HA5Kl9gVBkz2FpG542FZzfyp2JEmhQ7Fm+gvdQ/urckZKGR
dQihqz248EyCGhpDB+EaHukD6jySGrbSFn99maqYl1PcCZ5RRf6euoYye5xO1LWP
tPsUlYXnDU1gY3/k58EdwWH3/sOkVmVwr2eHkIVTcOO4UYUl4PxQnZeaK3apAjSE
5bFHa4NxGSXhMRw0r0lBaCCYo7gC3edF2PF1Xg0ZtVLOnAQhJvkMvlFy5pTgPA1j
DGPsnJ7guHP01ME6sgelpZIqivhK1Cg8XzDqRmoO0YdInWULgs3YKB0iX7X9CpfJ
BJ3q9vgAVEQquviegH0xf7+24QB+OMWVHzv5ehDUxYrVzeUNEw9K31Pt0f5AGo31
hVzec8k9NtsvP/pURkg+5lLvLWCwyftIe3fnma76XbDjDIm3/SdHBkXiPUCfBgU8
jyaMxYFzTMGxKllO274xh96+6tO4O8YpPut6iN1CmVbfRycV23zkr1uBohX9CHDC
9IgCre2//QLeMZ3D59EPMe3chBERaGgt18JXySHugpUm1KQXK1estPX5xfqrzhtc
5czXawxQ2uXFIYwApO9KQm+hbX3GMn98/5dRgFjP2I24tBmrtrCyERVY6VdbAWva
gB6b4mTjjk15nQAV+hbrSI5nYfO4s60UmNTbas+sHlFI+SasZhbUP3/3Dqpe6DjJ
0zxpLhUV1mHyAUmzLhFq4OCSyo89kruDw7KdluGaUQswQGYynCDuKu8QAjDDz1A8
/1B2LXdnyeMtTG2JTHNkZHYGQ27pyjxfSfrYVUEZnnwFBbb4Xk9JiywkfDYaX5Jv
THK2wZMGhHp4wlKGZR6Av3/F8+m072aoZt/1rF1Cyr6OVvOndh5+HrrHTr6Lt1Bo
9gV3J8EHxSFzP6ptUT7LRgq0DM8RGMSA3+Uy4nTgxI1vhGM/ug0mnYteJqKz40S+
FsbqN6RUnk8/DjLpxEz3iT48bbKeSxWNEcAAjxke2aCbSw2XceDKVPQDuLIZBY4R
etqMRARaUgPP/CS4M8c5XWMevxsbJ8YbCEBFEgmW3jgBLxL9l7YNlc5mK56k508R
CCFUYqQKyCQr1M+CGtf0A/okTy7e/G4CcL9Ljpz6BerO1PJqnKlWdiPq6YpIszsc
iv2sjGQRkyYyXAuR938dCCGCgAAiko6w18KGLNvjemA8jPCnkSUMXulNLvxUAp4x
O9Ri0Os1utQytNr0KdzRXHKlQmIGQ7FAaR3FO19Yhauiy45SBY/omn0PMN+WBw7D
2yDZ8JtzHuq0buXszUq9i+nbP0MjdCeaeOC/X9fuGZx3HoBGAlr1GZJuR+i+G/5x
speQZce1rfYRsnhVyh4rQsW0Ep13o3qoiiF3QUw5OjRnEiCHeWeSYQtV7+pHAvgE
4DQKjGpdPTrt5NPmrg5ZCX6p9J8kgqf9hqbNMV7Bt7ef9YqjEMl601P3DpALu7PK
XskNv9+wtSn+OhlGYI/y2KQHOdVea/v4Lf0LbgjioaZv960BUwl/hDzlIpTLF/nT
/A4C+wgXFnVtZCtoONDAIW35/xlKfogrrFEHF5KBjmVsN7pgoxdNT5YTc3R0zx13
sHop37QH002YXJZls8C46Bs03P7eReTRR6DXMeMM5kgPqDBs+AzCHVKFrVIfW7Db
jQQV8qwVSfxs+Uhozs2jA2PB1Ab6qTWKXeFD+oTNRt+Ortx1DaX0P+bOq9UNnOge
hGNjQ1jT4Oz1Vjl+j7LK8ua/SA5jaEar2HT3rkaS7KF0vAFv2zAc+DboxXjpVC1/
xavKeLD9jkolJfND6Q061m4TiOjcfiS+np05yseFykPjVbzarKwyZoX8PUHVZBt0
wOyumvM7rOf8h2DkX/qPD4LetCLNQaraJhiqzw6BPCHLZ1ZK8gnoFhBYxLocqbrH
lqiz7559qcxR1rmorZIDyYv9qhdsR12buoLiJFUCLBDfzJ2D1TO5VJYWL52x89lK
eolo01/Vymsj8Mb1QDQ4lE+LohO/Cf8MROierYVFpuDLnHAuWJlZEu/DWXmXfjMV
mW7WZhDIfnzTK/ty4tGy+LQvuAu4dXWf7qWJNIdhb4ZexPNsS8QRWwD05bLao/AW
DcQCmhkP/MTHvQFe3pQhQeLnGlNplyO5d69DFZkvMCiCnQZdmlX0ztixCZjA0T/W
Gx/2U39S0vi/3uDpL/vG6sk2SPgQFXbIn+7L/VNIY3fgIEILVIdyK7Xd3U/ZXlV3
qI96OxoQq1BG+Ky1se8Z2iuLAVDzxquCpSOiavDK6AmV+uBt7Xc4eEz1tKQDa8Bw
k/RRsMkjMFqd1cb4fOGzt3wSmVSeMN963bSp6UmylJazm0QQuCm4zZjdu7lkwMnq
iMv0MrdAd149JWxPpfERcDRTaUMfFy2Rze/jyfUoMfEANhLuvBsSXGmizcWVwqjj
2esWhiV0Bc4rWSb4zSEXtFnVvVQqQ//wFlpiqCpWGtrWw1okQu5QSvxMa+txA1Fd
ufF4CacedC21KjsxESlE0HfBgGTz7MFTJmzbV9EwMLTDrt18Yxsl/aypmbeNpxaK
smOHhpcQIqofrmXhlw5FAGm4x6Yl6GibEPQ6GV7L2LsJlmkRKH2/2Q2MhwG1TzlV
i2j5FMZQKoESaJxJHwZ7LliwdwHY63QymXKTb2YJvfM2lopHWkREf1RW6Ij9Cu0w
Vi18n6hlmhlVI3UZsrunmG3tAXlI/nkyC3GOEWuJdeWfGkh7jOUKFJWgsfYjPPvb
e0TB6Ls9rL/f/8Q4rMqEMBLQjql6PGxR4c6YHcnz2Xt5XrFE/CiUFQtXuCCBaaXL
ws2sQR6+gDf3oS6MTLrJuv1DidFum9jZ6a1MLSYtHeE2MFSwbtN016C0spZk3kRZ
GClHtZodw23+JlRKoHetPdiJwXTV7qezHqszpWcRZOHnFiPU13BgTqo3vdPSrYNY
PGUMBGqlHpaB03GgtpvvJ7bVYKcu2ASgs3cApbaDtgsd9g6PMzTPpS+CxF6xcl4D
Dc8ciIEpDd9ZgLP4xXmupus3qcEQOr3Ilkp+FzbDTVegH2TgPJKLk/jXfdAcyjP/
kHiIRis+ie4h3g7r+KeUwHMyDyrPDJskzFOqKluZ/JvCz0/bMhfQ7xKWAp3vFrI4
b66UepwNhEWH2pBGSIa7ymxudkXFWESMJff6bs4/u2q/MRbUTwt0cyHcUTkJPMIJ
a8VPra2Cno31lwHRjoDdbpjBSMxB9r2wtj9umwgNL2IedATg0v/7UpfA44XQ8v3T
7A+aPHfJZ++goWBOR/WV/8GRp1bbmj2pAwTGjbftnpDXTNq8XDYTShDe90xzNjnn
VZW/mRO4UkjzT3Qti08UmCS1IvxrmfsDEdKk/K326wf7NTF9lXufnAl+RnTVcKPB
cXQ7ya8DRp+HTIOyTJtUAhx419ASM1f7FTll6m/3dm6+xsEFOLtaxIU0AWn6Nkko
gQDVVA0qorpginIItpgSt11S8tNg7C/J5D9nSPlumN6h3XQAz3Ic4NI52qxTJfX7
pO0pTGF32i9zAJblSU++1B9T0cT47eyx6b4ZnBhZiGWxN7vyMGQpkaYIqZiXpUQE
6xU5o8GSuzZOXH9sWvoYGU09QN0NvQ6hlonJh6RNSU4EcR7Sez9NHvSuhywXXcla
/r2dKWZRIps9/YZt7WzXNT55Kynq7soauDeObfZx1Rv2/nHBgtOk+XAvSzzzW38i
ASUsd9bvPRP5cHh2YnMxWnxWsahB1ePXQU5oZ5bFhYUoaWtiC4LdRWOoAxg3Psp+
JraLQvqzTDCYRZviwmHQepihe1apELA0Fcs4kOhFJJMMW7W+B7tOjT/1Nlm5lglm
xV7TFbUCfh/d/tTERpSn3VoMaIthmOMQX3706G/j1ex2NdpH9D55i1pUdBw9TN1D
uR8T9xX6oznktcdoxB+nEX6usE4kDeJb931rU1MrMRutq0mvxkbL06ILsSOg8fQz
80cnhR95hnZA+FrpTfVvyoswL3FMkKtzLClW8kG8L2X29p7IqFhMJR5RfWGvr4mH
edlW2OQjqyTGihaIq9sYCxsT9BK5C+Pf/k5hht/NGIwx19B/OnYDvAz3XGAoU/jl
5bAqoHsv8AqgbLMqv2EbGGIBr6Q/5etpoONCrem2czy1U74FJqxGXvE0VAsUsyDE
GeIs8xVoijq0YIwgGqd+T/rQKVCr4g9kiRpwF+rcBBhiBW/hXv6w9+0c/p6cNlRD
gyrIcUu2w1Gb/6pPXQPoH+g2UihE8hNgoyma7/mnjjyJFL3ARVad6bOGSLzGpygE
CuAi7scA4u+AqXbhjghM8H+GleKzKAoxVUfceAU8zZV1TqlTAQgC5pC4U6bBz+9S
GYuPOp9cW4UV83zFR42eb6V4KnpSrvM5ldJRMVn1Ps5Pn+hAmmNTO8BdgfnmC7jw
aLbthv+Yxx0ddB9+V9aNMceXCkFrA/i21xcRpK9kbUSF4nFioUzfubKuRIXu+/e2
k7/VXyhifE5V9NA/d3hQ9VWZZex7gndYKXYnyxVbMY1SM7PZs5KTkNOMTF0GOQtB
A8BNZcMRGPb9H3RUsGpNftWWPESWFwY2+Rl8MPY7VUBB9/O2JdsBcveOLVgDCUBu
PLnNebwtzQwYnY+32A1sKst2IYLNxzJ8EHgDv5hV4Un9Orwm6MJDmBoVTXYvwIuV
IRVimKq1a8aSMJc3MV2BtkB3F9slHietRGVLWUi9S/qTwAs5UQ0lCtcqf1CT+zWf
kRncrEn2jmuj36P7BbDrvC/blUulZUpJX8qkgCdmpcvipHi3hiA8ditv/93mmLco
KpfBXR9Of9xaQI2ZV6UeDDt3O7cdJyOrdkdzxFnQvY3+oybr9zgMIUIVIlK7YEbi
G0boS29L8EhxXmehO85B52pG8kZCBGSU/J2j/28Qfs944+BTeRsRf/zrpCbuFvkd
bur1/imKH8h1DEa45hxjtrpTK4DVWS+3AQLiD2Lg7WTtuNCCUkaFq3k3Wry26nZ3
BniAZl8DjC6Mog749lwDNYiHsKs9Gkc6Eqw7Y/L94vbuCTEHK8/8CK8ZAjlyReQR
VT3XY0uUd8ONrBBBIpSI+zGRgnFwAAtXPFnbIaFXG7Bm0yqnDxfBt1kBwmRIwjoT
FgDOPSDKM9BSsVY6DcwVtE+HtJJvEmzcNwEgXSVQnKaLBmviraESdufINtrkRRzm
7TgDhR06m2cIoE/yeH9zs91vvSEk2KRdE1Viz2VA527wPEGxTg4u+8YLwKCh7SUl
tLbAaZygvwurR2QnJ7Rmruv0jAOyfWCQnmLyYQCNU2X37uL85+Vt7hpahUWCXnxB
W44y/lr4E8fuLIe5oc+oaaJRw5vok3vfS+4hg4JkhsshKTB8gDsPzIukqWj/Ob2I
kQAzd5pWAkwcUrvJzSNdbeYRbH1ih+2oa8IUB400wJYE6apFLOoWfbnlVRcexmEr
ffRzdCcPD1G3QlrVkCqGjaOl2EdF1RQR2mYjh6scPlpLha5+iJPk0Kb8gUzb6LXe
UZN+gITVZqY++sErL5zq5a9tdF1Wpc4oGm9rvFG5RMH6uV3rpNtrYejmnd4jtOSC
aZhOGYiUNDRSsrfT/2n6+fbDo413UPL01WI8sLwvy1zDsD0UqdS7HL1QR4LiOonU
m8lXo5OUuGxvM8nITY5YDYzXCrb2z1jorTo1W5tYcvseJyWsT3kQLPlRth1jVu7t
i5DnQAyiuBl9gnXMVnq7++GzbZN5ybb5pfvFqm+p+jTrajLPYuiyZviR0KOfVjKg
+mNqL8SBgTteas71fE5/Qyqp7nLRKz+65he/U81pspq8eL2UVvXZQ7OZEfg7VzqF
XpqPJxx91m280nW/Q0dS3rQtP5lEZeRvPSfPUzRUD5o6+bnLCtAftZQDLqquTsks
1aegzj7T2hrL9X+FXXMprNVEO89uEvgyrsWeptsWiZnu4YD9ze/IqxXCDLMmUhWH
xx8mnCDtDQIIEcFfcldimZbF0m1Nks4GE8O+U2Du/B1BYqmi1XgNrT+1MbxvsOWw
yP98CW6dFNycFzMdFaXB6C07ZGo/oG8wZwzUsse4akvd6VxwDMBk03rfIDK5zG0G
Olb5oklpyZ11aq82XEl3wMysElEB/WcMrQ3iZLYCd1WOKCcRDj348+TKnR3Jl0a1
wWULPE+VJm42u28y6K47t30NtjM5tA1fCPY5KdPDkdRYBeZQbK/sJxcaBojl50Yr
m1Ku3B29v5CIPR5HLZCyjFaEmwhFuK0HJKE8842pW8i54vdU5HFmhdA95gW/Zdyy
5hZFCfh3e6VGvBBlQ/wRx1pZzVEJkcCmn5rsXBuVup/vZQN/evSTWHhAFswO2i5H
+z76WLgTyx8/jNgc2Ljxbvgh+TD8bBwlQi3XkeBQR68I/Ny0d/uP0Gr3+U91qyPn
AvwVzvVoHcSQIAws2IqCAL7IG2HrD4msdOqV+2h2dayMDv1HIZ4nQ+JJKqL2Ufjf
x589qRZ7rSr8zjPZVDnSLpKOl+UTahNl7ZSOVqyn/c/rC3/D7sZtcHchd+Gp9xlz
YIX08WcsfiTJAYXlBhVB3a9h0wd1220L89nGOvrI0npWaPpOPbU0fbNeGbRPmX/p
8KO1qkwDuOl910OZ9J9/fQQ/Y3gu/PDH4c805t6QFGHVd9NICpPk0KKHjZyef7lB
zT0ZTpl+Lu1Yfb21zxPbrIxFYBxL9CSvNMJIB9KcCrLdpZ8MvSoJ3S9RWTidHqwi
M+N3/aS6nge7Ipw9B61a6tV9JIHKsqGxxsi/RiEwheip1xaZj+UjBDBqw0/NYTFr
LWatBGURClHdUJGCQJyQU63+SQymCWreCxqGVeYCno69u/uvUBuuyu3GPcnRVmHr
+75fV3LkbrtIj+NIwCe8ttbDvdcO/TbMgcR5T8u4LLFrhavFkERsaRPa+q6er/p1
qTP0PutFo0puJJJZQWsJXJYzpz0kOLnwQ0uKLEyj79C9KJ37cuRX94Qd25Ey/5EV
TsdAJXUvQdZ6ufHi4LoQl5IHrEnD7RktA3KHM125OkVBZV3WYOflHiexw0PfKx/R
55om/f8WL/hoETTZ+FtvEqCjQ/JeRmQ+K+sOdPjqhlopAU5niKwzYtxySqah/ks8
yOVSlBIOf2sK346zWvurp1asrf5ngsKfL9ekQ5n4OdbLiNneyFKyZtenQ210uEdu
bifRlfn33w2+RTX6ZJvwuz6OaiibA0JhB0oit4ISX4HXzf3CkavNTHD1/yLigFdX
BGhfcbbIWdBSMd1egx+MzpzyKjVSbK2yQxguxSbAl5Wxp64ybfO2ilmSj41UEM61
Q2sm3q33uUJ7ZJE6bfJ49re08ffoUdC9GQ8kVXT/XCpTZAKlcQs3C7xSSdCCZ9uT
qT30G8C5m9Ykp5oNuyDnfYuBHhHKKvcL4GImAWHEMaEWLLgUgR8tAqNYk8X9/txJ
kdgHG2VBM39ZBVjPMmY8gl0q5IMeZFkG2GdzcLbRcC2WapjMtKxhtt3Omj0dmdZh
DS98UcMdKYUAxrE9W/EGROXL6IFB1mAzzriTcSX81ifLsp7yeMzktzzOZHwU30HK
hCgd+yNWIm11lJi4ajgkZ6CtnJ7jYWrxMd9q1v6iaqfPx5RC9SkTBxAEX7xiXKvw
bENnRSOceTLYhChU5Rg8fcKpTwoSQLNPGf4LGV11XFFqdoNBwCbmZkHfpx/hrjRm
qwKsm0KR8/AsfW8b1PfuUfx7EGvr+PXL4AEXcToLeAhzaL/ZVEG+XSpgcJwT5wf7
c6p9XZjjqJzKK0/l+rbDwQSpTN2v0iAsOcsjprzvv3LdjGT3ed6R+9wEGqgg11Cf
CmaxYa59LR2Gnoran+vrTsHRiRcQ0v35gQgSYzURe+2SFK6Hsz4yuUU3C4O6Db/W
2NSdS8bMuVUQ65GcOoxai6aKi4vRqX77qOikHYT73a6bCeBQeTpOGM2pkl5y3Pgi
HSzK4KqGc6g2NYrQDWRlPL8zRgN3OlRNk4OTIMarq0B42vC0AKHKwkBomiCbZaMm
nwAx1/tENOgiVjll8aBXUeaJTj4bpZQZMc71Z4vuidBRTrVJOuvnMP7WsbXtpyXJ
mr/KKMtNFVxYBWJJIJNzg2aJVLhk5DF4m0A3X4KJeDamt1c8cLbNDqEuuRQEYkuU
c3TKkF08ZpxjTugkQKa+DG3sgc2w2oGU5ArWVmPPdxSIAOqOJzrOIHyY2EIx84Q4
s5B2RX6AsOn1lVDwDbpY/DUn8yhgvO1FcebTsKZ/DsAt83on1k6y49m8MYUkgYkp
UdIHIL+k3Qv/CokPwq1V42MSCwu0kJHCuXXKGskdGZunOKf5wneBxRF2IRq7IJrS
SMo/O/D+crXuYeRmgirsW9XVeDLrMXdbVJJTo8reJy8B06TzINmvDKbXw7OwMWvF
0asYG5rXhho5W+p39sh2hHIJo7PIZdF/oX57pYPJErER+5fAtVp4WEbTwpFC2sAT
/Xg5wTysmBL8/3CxRAo7KPZBedtcZf8jilzDTLHwZXZAcc0NJjMBO/RTVLV6upKx
XYDjas5YDg0+0ZpHiZG1G5N9lCUUU3omnQEEWNFlC7mjpQWL7cUoPGB3d3hUpNDz
d/W5lHk2U/PXHehVKn3dvvO2/z2x5OLxCLzIiABN9ePaV8rDD8CNcxGsNpb74bRC
xnQc8NYW3GS101NKYaR9IH2KHAh5z5GMdZUXvMVmMQaBRSRNfxTIojmvYTgP5l8F
qzrGQpwnJa35yACtw6MhSIxypBq6NSFJgVBFIJmFcttc/2Dvu5N/NMvvAI97nyjU
6F/VcGngpen8k1yiR3LdNkJYUriEUWz+1+6Rr4cO44MSzSa2ENdHid82qazYH6Ac
lPB/8Auzj/2SwQ29HXjlcaGPAGc00TtcahDd9Tk6cmxmFVD4VmioYtugPuiIGxnm
iKMavunZ5lH6l79Tssv1oFQX7igYHh4YXtsTZyvNxLwcBpuN5OXn8FsmF54+LfaD
ZGBEXT22H0NsqjlDBnUDcw/XwAPDdfndhMClhDj0ndqnVBq02CcCJMfd8lxTxV7U
8Oa/Y9o0WCSAa535k7uK/VvzWx3ma4X+L8qGkNPL8F4LBtggV5256IF/Fu/9zYly
MjanG5jzy8eC0LVkNKqMUVEA1qiG8bo1z39O9dLIpwtdbfwHdc8eo02I4X0UC1Xw
1M3W+lSTRy5vzVymlK+DV9QJG2MNsA56mTrbZmY+aMwUOF34QM5kXdEhMKYTtO6O
ZCW7TkImrACEWQJDgtEeDgZAbSxBe51ciiDpbn3wO+4Aydwjsl+mdFqKUqiSsAqQ
F0FzFzoGnA27qezn1Z9hHluD84kSWi3ccWbfTcx3LM4X5Mybu+uam3uXURECQuB0
+s2tRrCqXGMQ+EIz9ECFt2mILC0y8cL/uSGJ6fbYO/1JuSFWMUDIPSXPms/JG3I0
raT7XLex9eRLoTGHDSqjNaa+YqA2O83Zv0LjnhMLr2fShcctpnIZb2pH9q+lsSK5
uKPrt0HTaKj6UhpuxCgA7o6LR64DZOSpMj0t1nO85NI70aaUFInnOlfGSh4NLYDi
v2yf3ciUSXmFs20Uwf1o19YuDVbQ27QvxmJkwz58Qac+kDp8oqlrllW2NHLdQ0IE
5RDQER+HX202HycsyPC0YK6BgcWZVONAZLA4vuJz89+ySFRB/kUCZ/YuW4E7GDx7
ZdOpTclUEltnAQlc3dWbJeGRkGEDDAPt2xIsS5PPTVZH+olfsd1DABbAPko4A0zC
4oLJIIqlxDmp85zA6OTKJsaOkTew4gPZ1hEwbuetpsEh/Rp7QSTPRfAsRPiJqCXR
/FjmShbvIjU0FUzrjSw063b6s6dqtuO3lOfTP/QHKDZogUatm0AYnT4HZi3QXeV1
c7cifoDkblMB6AJtNhp/2uP7Q5+WLJqpOCWI6NmIkKcTOm5Y868Yv+CXVVC5Y/+v
vgf0dKa2xqvxbm8shdc5WvCQVWtRoqqSOgzVwATn15xYZv19vndCf11J3a/Tl6K4
rh+NLn5OqV0hnoiW4ePkZ7pMYMx2N66HwVinDLYOrh2KFY0e0Y4myZV+V3r5crs/
0yNLKyCuutYSXe7N3tACz/6UwpmbSo6VAh2f5Kwlg2QXse+yiOt3nE/NtT4QASHc
kclWmmUI4hIUDCE4lMVWDkxoMVRt0uwRd7TOaxRhnIezmbgKGan4R/u5rK9hGmZK
AGi9uZv8pn/cjUBLU84eF4My2hv3sDm20W6wh8NWHU7D4JO+HaYiBamC3e3K0G1B
bJLR+G70am02x/QfI5qaHDa2aiWIeIafEl8eD31BnQptCQD1ec5Gb/+F8AA/OK0z
ijm53YlRzCmSsD+zJLPJeWHR51CEJaK4SMzFTs79W4/IT5lp/7EXGglJOpBSoKgq
RMsYkZpGl2V5S2zJA+nxG2pu/7C4tDpTYe4xB6UKG0nVmR8rQiylm/ddQhNbI6RQ
LFYKA8JQqyYmMjuE2PHgBCI6Q6ln+GDdi/xEYlZEoVGRb3C+rJriKTtUypFwnnV3
IGAqYWCP9YoIyWr4EBXLD5/I6RW9lPHrnKHfo3Xv/81p/tDLz3zhdxuz4rdDKcbN
xaYt/ti71sLsO59U3CW5iNjsyqQ32iAqRZwy755dw+K9TgOBcfZ75x1T6ZyEOS+w
hMvVZsU1+zJGOw+f3zq11ynTTPOoWudtPVlo7Sbpvx4x8bEFKrnjAfFZi05Of3mK
1B79vpUKow3v20T6QFGvJcDyddnTn/9BHQ5aFcALUUX7d7FI+s2+gAF5J16HRxC+
z6d8ePBw8+XA9ogzAb55GcA9oqZVqxvlWRVnLqCnc8bx2hWyTbqJtHMauJCjrZCp
FFxPUSD7WANuaC9uxkOesnLNBCHqJ1qSmQubWC8wItoJAxSgoKlWDik5N6O3vscb
ALTl3pblYI762TZIyAQOkInixqo1oBMQIknGeLQFAdGVXCyCD6Tjg2R7z/Tk/fNw
MtNaAs6JFLLHJ6azQBYdAYdeDMwIcOM35vx52nu6Fc+wN+xnhywHExBFsJ+Hitbf
EEDvQsnbj+NKAskCw1lR/lGbG3ugSg0GSKtz/I+MjW0q38YZqZPCEqGVDG6ki0Bx
pAXgrX7Cdu7WcXSNpgjnyd8T8YYj6Y9s+xwp5qp0PsBsQRYWpm6l+ZQWtV8E5RMt
Hd2MkA9sN+1ViWqi8lu6Q/ropPGr5CtYAAd41FoY5+4i2qlfD54x4wAgvU//xahl
cxbJjj/tUy0dUwMzPc+171zv5Fklis3K71+s9M7eje2xopv7gIV+cmBzJr8RJbSF
uMMF//Z0lip0LOISVZbBiuWQCB69c1eDHfsw3vOqo53K7xkWT3vkFuK5VsjGkKU/
QRa9uLo7x8NK9kO9akzkbkt91IMG/qG/hEaohiYxZSb4SZb9mvZwEUN1nMybGX5h
CPpUw00RXsjb5+iYCxXnRlt+PZ8cjsoP6weY0cRgXh/LArTd+tTzi1SX4ImasQoq
b33UAw8cUK+ehNPAukULcYVtil/7/8LTZtekgIxRrkh0FJGTZoILndzK7o79pkjK
nivcC9hyhKJydvmyg8zTRD9aRdXTIuIYS9couIi+9LlRlWhnjNS/jkB4dAhzzzD+
/Uxhbs/riw+Bz692aY5qdpEeH/MucXpbAgci2jT9FYI6+2WIKsltsHZpaHdE3oNb
oNQCwXRz1OynjejLheE0UQoPo8Qc2gazmrFdJiminyjK7soamA2Uy6ZTz4idm+ai
d/HGU3Z6zsFVoUApFU+9VCB7mkECeCXBN5YpygKXL7KrnMwSsKvgupUTeUvjhXw+
KDST8wsqSwSxl7vSH4nq8uz9F99WNyNwntrg87HaukP+ymeJGGDLNisJXRjBUXKe
/lVEIZ/CdKhKBhUkR0OivFBJ86qR78yXC+q/V0DIBEopWRrcFEzffuxr5Fap38a+
kHF7xAgUFGXfKD/qlK7sWYwU3wropvPSHXuChPew/KSGDn0c/ZYGmtu+hvaG7qWw
vr4wVwXPtxthDMXXyKvmdSsohpd9awncBRJ75J8lHYSTtgoWZyNuLEmGwwPEa4j9
d2JtrGEA/TRXELvEGzbM1TCFvoGh7ageUL6exyv5yKEhPi7WHpYyzadWdqNJKlsV
buNokTKoiWKCOs+R4bvHn9qSFSxnAmBKV58l602S66S0IV70C1C4mIZYduD/B/Z/
PGZmEdhhf8vpLHoo/GJTznEwFBBrRLCYrf5hOQ55eqFBu5QBQLP8S77VBgw8Ywjj
9oZPu78zo9pibS3juZgL2hQYZJ2T59ZSkR6QKKIsuueV9qWFi1U0T18LNcJpz2rk
9XmKNsnF0kNGiJUlxAzB+wGwYLNWPG3e0sQZq80brtnh/Qu4SS+nYBf79yPYKbCN
PFLMYoAaXRLZ9h1CIlHXvNX9763JgzujbuWTxsUUVqfpGJQj8NyLNl/W1dlm+TCG
Oz7QxIlFbI4olEH3cgcCuAJo/Q40aCEAcUhyRUMMV9lvZZq54xOofibBHME/0pY4
vvXuZyyRU9zmzonckxhVT8sTEFgga8NSiAj7WR5yaY4xOv3nsS630/eFOQQ+y2E5
uBe5lCGyp6F0kCwSrt8ojHoBP4sL4aQ3g3cj6fXoUGzjKUCSzq87ESCindbo0Rn+
z5M4859IcIuL6OIPPsHYC00+2FozKdoR5uFGZd8+OfEGbsM9djEhznqTjOcoqvhH
WnkRPD5aNvJIkjB5Cp70JuSV9lWZpbvxNUljvpuHBgDoTqDVctRgG78fTU4rgVgK
moFZOQ3bKYXKM5rfdM6LnUV37Z+X9+FJAVqcizhgHnWTCh5EJhTgsEktw/x6M8zD
ejQjPlQ3jv+D7ynztJ44juk1mDhShdzjOkgpsbCp0dIN3TmaXcy/djYN/Wa/E55v
00r6//Q+iEPqpQJtbxmS/O+W89LT1FrGqpqyvhwQBL4EVSKCJ7o19Z3wcm41RRMQ
yph7KZEAxkvJhBYsiyeik33XgYoq/KJfeeLfbrIPQUniEmbTl8YlEX275XuFU6Zq
A/k5AEbgoWs/4T4Y1E/4VXecFz7FCccVCmdEpnt5kJ6V51wAKZWAp37OY68dLnkV
G3BFnjuvaVUmIXQ3M12UimFXbCjm/csCA8G3VnCZ5AHMD0+kjO2HBfFJEFvdX6OG
LGwqL1eU9gYkmMsu0gI4OXlpWndyEoRyotZ/oQyYuBZTEgGg4L6rNHRS6iR1VCpW
zZ0jFbPUUh4OFGRi9njnCeKe2ycnGtfMwlpNhW7xurQWREoKAi0neilcZfjmU+ip
I76LeRUwb4ezGUCNS/DNLPHrDSUPY6ycHfXtCLhIlvbdCKA1r7RaGxN+5Qr9nc6g
vfMtx64JgGALMuyYN5WcDzTxunY6QCY9djiMvWyXs18mRXBjx317Iiw0yKZcYnkv
gHqQQejPsdG5tsdRiKiUNB5h0PWmtucqG9TkMjvSfirgGUSdE1V5VgMBwUbFn3ja
J5LItB41srefrIiedmn7MI6gaA5orgGBNFTWhQ12LezoIgD7aD/8hvWg4gINflLa
18W1cAji/YfLcoA2rpBFgmDTQR2o0mkkDlnqeAlY5DLvi4TK2RYKO0lFVadHU4qh
0EopQe+x1xor9CxbAcvwN4acqtuRXaVCHL4DtUElTVkamUTYCVs1zPR0HNN7YYTg
DddFHHAMaCCGhqe5uGGE9/O7V+DeWxaTxvbl1NPupvBdOztL2oChQduK/JejGwwN
4FsdUFEhOoMzWq8G9I8qMOqbsVmRmkwh5uEVhLFCn4h0F0HgzayH4JXUD+QmWd4W
PqgiWc6GU565wbKGEXGDAgKK/3YzGuLZ8pR1ksqubdgV4QsTh4uHqfeCbLBpbXz7
tj5rLnkUD19LBNWEN7R4oQB/oemW2/V701UvnJA7v/K3u7LxE7MF0xCUX0w/deho
ajUsr8Gcai0FGw9mt2wu0uhzVMyH3mdqByPGNckNEkehVTH3YIfvFAeVKRgphdea
kfnWRj5XYGIoHF+Je6LxR/D5ZEXt7tTkG8A/e1s2jxgfs8v0PswQd5Ly5oqX9KP4
7c8bFQlbrXZZhsur0/a3nmOx8f3wvUgXzeJqSMxoMWfHVOGcvdBBGeLXxv2/A0de
UJ1DBNFMwjG8o0pW5uHa7j8wIONXbNGJ9od9EoolZ26MRM5lLEcMCJbzlWJuyOrm
G/ubf+p9N8vW2DAS7HPK7z264LzoW1hS80K7fcN+CNiGNHSZX3KvyNn0S7Qxx6WD
tz38N4voistq8XgkK1/FwJd8dG6ZgvxpXGHDhEE+lQR87s0nADa3FjyF554YRdSd
MSQz2L5Oub7HI3//m0ziOnSS35gWyyNrZi2wX3M4KLrn6/JXWvhSkD5k40DoNn35
ujMz21msWnJ+56hHC7kVrW0Zfnhx++y5h2z+g9W/O+o5i+SvpocswFh2S+ZsbrYg
y2w2/6DHhg3xFTlhI6E6khHIKEd68BIKRnd81uamvUC4B7bPjUXdeFC2lJ++ykeC
W2dxPkaHUvfbnp6+rmOmaGyQtcdrwMh0iDhnhHBVECSUml1y5C0BlqbTzj3m3iA6
Li9F7pPwtubCAIG54anh3ixn9TSnoGh38lN/W+3o9hi+N+mLAAy+y530PGrMDWcp
XS+tfd04rn7Y8Nrz81/EuokQNJxDDp9pnx6G2uBIYbpFKTFnhhROlVNHD00g6/it
peKSw7BVNUbFJtS97kr2qpVV0wvuxMT0iDx/aO+oIL1GtvzG5+Ki/I18IrShkuaF
dGrr9o6sZQjCujyjTGCEb87OfhUBAFNs1RoZEbGLZjA/lQusL+j/v7Ewv9RQ2BeM
t0DAJ+/NGSp9/3H4SAwfPuERUjNsD5K29e048qFxrTQwDlxH6xncr0/EifbbYKyV
YAi7chz50e/WtHMt24FQsekg10iQuxZ0kl0bptD7NAK1SjhSiUs4mWYqMcP1AJwK
zTiYqnwiFx5wmiH0A346dK1kjKr21YRZumCAmYc18TQYs9QaLHE4NSZzIkvkFQDs
NCAHnnSCssvAJ57EXsHVUY/6XtxiHzrjpzAkUCFRZq83CddV/AshMdoe4elkG1uR
E1wXK6Y3C3MRZUh20Lw7RK+aBAjnN8QYiCgVutLdGUMUpYPACSISSZFxGgNxavxp
uaTEK8lZ3Bvq9wBLx+gvn4UNHDo9UWLO5kMw0Y4D+FK5xX3J1tE1q4Ma74CRP2CB
tAiohcA8Oz8Zb9blqqfvqDcryzSJYouuBAybKsj7doXuceUd5XZKrkiN00SbLioE
vFSwKPvX7K2KE7AfvlLdszopYybiLTMzEl/45LD0Ga05U5wBkqf2sJ6DJkQ6RrBn
eq/g/O5v/3cnVHZ1XV7wR+J0pwxjlum7WCUQxFOFdgkrVs9wZzYBVTHU+DQL7K3c
qkiU7MoRMkMyLdbg6dhZCCkZCGOG53/aJB+0luxo/dwRpmY4w8OOg909E1Eu9A/l
ouBRQnYfnOp3oKJW6OlMJdgFFvAF0aR9DvKLYmqlzAMYhStWEhd4Z0JSWv33LDPk
WW5UrgRqmboArBRUOdZc4k1A169ErCV8JCztntsH7BtaINt0ix/tF1wq7ZqWxvgz
lBJiKfmCA5MMaBqMbPmNw4UEyvGsG+ggY7EVDrPhoaWgRhiVTAe1azi2Zn0xx48H
HBJQZaLFHw93hQhc90s7iDj80OBkN062ppGHhZbn39cU8szdztDsHJR52DmLyHHb
mFKXZ+iXgNnu78QI83rxfwN6IEeZgLjPnUlMvgO0LWuTGiCJuT673XgJs8kryFu5
0DV5wC4I7nTUkqv642Pp1Z0v2lc4kc4E6uPwU9S3VVa8ik2Tffn+XbMoeYftNh3Y
3Itm1XY2iiWeFHIWuPCq3HfYkn5B3fdcXsMLqF471CNgL9IQE8TJNmoBYDwDOcU/
aqQYOiJHCz/Rj68cO5G3ywvMr5dtnK0Da67prbDidId66RqNSBBOKiFCAWXRYllI
kpZrrTnGBDlswPQsHk+/7/ZpnaK/vHa28XyKfz3iLcsuoTFJ8hl/aK0Mdo4RZxHz
6HiOabte0DTm3rN5aoeVmkJV8BO2uKVkefU+y9kHYCKK4LIpwUfJ9H4E3hitGAkV
IYdcjwk87ZGGEWc+90aeyBGUp5vgrMenUl17HFxQvJsHb/bYLL+NQ879+PAUZxpQ
MEI4bfrjyILGP64pMAiWTzxIJVXMv5tnlqLaTbsV6GVlOjqZU0/3klScb2dSADib
q+hDSk0X66DAtQq02pLgc/H4mxZQ7g0GOUk+k3wpInf6HBV3N619jusQuyaQnFJ8
5U80oVq4exmLU4r+oMVh1aS6glDA++FXtiwM4RSK3urV291/GX2hRTqxIOYPr+PS
VP1hpYzd2/UcNufrk7qRzUtqENvdEvxkIrVU3Hkhw9f0quaQW2VW/iZc5UxxIYtD
vOfHWkT17qNjKyc44IdYIKlh7VJw9pc+XA52QPdC0ZAsfUwvlfS2+ZDQgS42nUkD
2I72CQJq75qncdT+bX7WUXnijIr2StFpaVPe8cEawfwSVfAyhheEyYnMZgd98UkV
3ixri3N3Ld7DBG1SZPH9jmp5Jw3TpE739H7D9aGow0lCMgbCFu0Hy7oskl95+zaT
MpG4OEAvl69WNzk6snXh0GUESQgPvJlYbcqkwlqs4cIJ3Is5n8POdSuQOkXTJnwg
VapbbSmy4eyoqNNh/4rJy+HYDH2RVbfBTtvNdjy1ZMLR9mJ1SH3cFyDBYcSasVOs
ilymBvPAQfQ3beptbYlOadn+AZjSpEkgc4ctYFzh2GXBCK5hZIXAFK/7T5BPBz9V
w6ghQk5Ph0qXUKN9+3uwzmFyIIBw6JJLGnCRi2zhU8WEkhlI89IUfI508kUJL6UU
sDKCI7g3onb/54cAdhIy5AjRvVB1YaJ1gB4eN9tfWtiMR75xyq/55kTtGVtXcq9j
we2MY+vyHMp9aXs2Dz2CWGQtumJQDBh+J+zCmH9MIMO2IrFATSjJ+EWV/pQacuWP
HxoFT2TCPn0OecT++rNq9YJNfi5joJbKneGaxZrf40pnedJZXhEDj3y7bmI8tT9z
DVd9a7ZflHTzxpK+eTqYzT4KlIYt5dMpIoA8cftetNe04uruqE32pFE++rDEd/z7
qRQxS00KzKJH8jVBWYlHaL5Xb8BUexx4qIqAhMMj3jEDEfRR2LybR5bUUIK1yKtP
bvS6diTe3Fnv7SgwVbMAi9eev7s7ysWVXaHrjayRHm93ojWAB7k0Ss8IqlvEQkG9
FbDmdm9PVlRjIcBGb6QD1BTxANDlYSCwUrplpH/ADxGf3ptvSpRD+aEAoAUru0SO
TpO8l9zaPMH1rl+DTOfRklWcCfx9ZWO4GQ7IJyWlnoyoyG6buCvcMuXjNsqP+5JE
kd58X49MzrC7oLmEU1F3LBGMErQ0qIEGhQi4vBE5FKnE55SxmbS/1RqBz0bCMYhM
K73WRH/0+eQDLqNI+kkripK5wA3qcugeP6ru9G+xiU1TeGt1yfnDCVIoZnCv6p1b
qMe10X5WPd84o7jsfVObdCOCOBCbrayIJAd0yClPbr621aDvgHsezFGGpTDLY9AG
spyb77oU2b2V+y/CPDT5lxcIDM9cnhQl4calhMaa/0cB9wXZMcN1hSwNzlb/yNMt
iLZLYDXuSv1TFuu+K9vpVo1cuMk4c+YtxxQXpiScAd9sRQob7SsLn53W2MrXILJy
BF8Y4xULFZB9QTGPqJsMGY9sbd+PwV3Q0VapAv0L2hIY8vo6h9SS6PJInbPBd9IL
kzZX9nvRuJ0tIO5KzzCfBVFaMkHiENj1qc/rpllozQNnPsKV3PEJJaeGgK3nZDjy
ZpCRLKuMqxA0cdhwxucwbSUAqt61uUkDABYAiipQO/LD/DSo0PP8e0leCHmP1Tir
bViQ3PGK7mga+5ZSLFSBphIlHRCNO9Tg0ytR4xJ+LJUm5QtOb/giK+OLQV4gXnnQ
WhQpHlKgmrxw4XiuQy6++D3Uee4Yjlf2Nd5/Hz8RPGp6ALrsbyWicq9GiwEnhVRm
AuahmI5o7maNBJ2sP47ZutD7A4VvGe+lJdMYDrUbCk2imOFccU70HPiagDfKIYCm
aePqgeCeWdG6y35yw6Cn4+CVVTXkGh8BeBJ9gVQXIMn5upRsPEcRwlJglTPr/XAF
pXUOuN0tSnUlgSanKeWnKzciVMFk8wMHKyuB+O/XJtPbUEPpPr8Q9SlB22eekkNk
4Uzko7k1BNeGISTCsqpWM1ojwK3VioRg/47h3Jln4MDPegKSeq/3ceVo0oIKedlk
M/VB16AaWlWlVrLKB+nzFtE5K9WsHXeDpHa4SdsdiNByjKE2/CX9Gnkanfdad6ft
q+tyCBuSnIxvSIV2b2Jr3q0XH14Y/Hr5QSFqJCDGAnnqQSgUoe0AXJcZpZukD6G7
uIGR1PIj+ekSBoma+3stODmOm2lnfKyIKDmDqt5wSqYno37/xOO33O1nKjEWUa2q
hgfG0pM1/bwmVNEuJ7qEwhDeQz1L2ToRuC4FPozrcpXIbGgvOO3azaGvy8mLow1k
AcXgCvBiEXt2wC4/OxdNQFMGBq0wtQ5UxjndS9dIChM2RLInp/OGp20WQrTlYdLD
LTrY85GdfGWT6QzbhtK2Cx0JIPHoIuE3XeBKQaFYKukBzcBho68RMAWj0pmDrkE6
2lbMoI0aBeHWikH0IKylLKoYZ87tD4qDYoHgTO3vSdgxEUqlr/9wLLN2WbWxZRna
IJTNORgPIHueIrsHd1ohaLWESEoee/obsZ8/F5WhK4RQemdtdOH6Kqyko+ivCHJv
aonbQiGxiS634g6POxbJ5T/ciig6iAsRdZNwWkloUhduE5LIYGMH0oE6bXRTMEBr
hXowj2Jy7CvU48gA3/bky4NNieH4HdndR26cVFQpJ0BPCFIbxPdD6yw0E9XYDjXJ
Gg6XxPjZ6l9OxCp80GmkdXZM8/1VIvSW//z69/ioL0WQbHKhMv/N5/CsGlF8fJf0
UWXVN2tqGllLuUj2lxVhCR9asoVMQycKVi0eA1LTSLtg+Uor/wZJLJqH9qYFv7gg
XQ6YPeTAmPgIbkIEVFwd96XcH12AecY1XR//5A5w0651x85D4UylRSkRZVM+6C7u
MiGVvh7vqrNZ7Z2RtSKIqqJyYqaG0fCd6Mj313Pct3DtUEsg1VwJ/qlVmLx+XPZk
YjkXucO/cVlYw/26lS+ThOADFPGzWWaxwNCIBp1CKHni1RC+zu3kfrMKv/XucfKF
E/iplXo7znZpDrnjXB3lsL6B2nTEUD3jnfP98HBlv2IPoQMk9j8EgFhi4rn8L/GY
Ig9Ai5YydCuwI89Y/0VybSapxsHGFwHmCPdYL9euf73BQqezocPyZ665TXnlZCyz
5A1Q0B5CgEZlXngcvj9WpaI7oHNzY2EbCPBBtkVbKjjvLaomDg5XS740JOlNL2u/
Z1wxM/q4A/aZSvzNbIoKvwkZax78GqnLKKVSV9uid43mohGEx+Tsp87WyDXrJJoM
uDykcEKz8yDMiINkjbZg8y5Lzh3IVoJNFuORKtXZQY4AimUhssagmi1IjSqrDMxX
DiuyVc6Rr4n1/tga1ZJI7QF5eV4pnMeuV57Ueb05SVfmbIN1mZrOu4XrKs8FZieq
uH11hr4S77u6fg9MPCIzmTJVeQBvgU0s69SQbkQe94H4NkUXoQUp2MFs+3ugKQvd
r52LgvBEkRoBc8OAjLYEY4idkLVaTX6L0vbCBuEE/LJti+JoBlxRWOzcZbOWcFuG
ydoqJ+xxxUezGU24TgcnkOGghYp1SngjnMaXxr9N1IO4vLhgEBekVWsvomR67GPH
zKr0QOGGo79m3tozWUQShcBC2Bc0Hq3ltlHMktfZOs5oQ1DFWz0BXxcyY82ClLO8
D8ANNeFcnzRMDiQt4XK5kQkdNw4eobYKATD8B9NyBfZQf5Lz8QPRtoOUhS/V7djR
JXYqnS8QpxOKWsrTv+2CINo58yAjJyxuUqZWJ71H0WIL3/xsNu16IsceKlWAeX4L
iI8uShMo3OBIKl/tDtNeEHEDaWNsDgDqjIpv0Y/ewZtXl4pmqKbwjaVzJmOh3omo
+uMGBD5uIv+UDTem4m3CJCQDycQecNVBOZudKxVFKs0ie0Bj2ZEN/yd8R/sm2bJJ
CZnlLUq0mczrPg6cX8nvmJYCTrxdkQiguCL8T7wlxlzSaLpGM4+ADofICUsUF2Og
hiRWtdg5z+F4E7liEuHDw1D0KvFkPoVijoCzKO9OuB1/YUYuq05XsPzI8AY+r3K6
XYjP+fbWektyv0mYnxuoo19KQoaQxa5T4bSHtmp3i6lg0Cqvu6ax1mIfCNhpqN3A
uLPKjKDe93CaArFbXA4VBebmF1exEaKPdg7KBryYX3iXQtfNxcVRNxGuL/pBYbfV
tb7ZD4oIq+2Pzb+P6U8LXpA09fBkXRZq4obYmmOToTlPbOjPQ/65rak776+L3u0r
Yx5D4zAqkPTHFJndUgh5z/fAr3fhaaME1Q3gzg2UzdsEvZb9GYkTJbeo2xLtgrIH
OeNgtXrUVheFKyhDuSGYSzkl0gyl7pzPUJLC0AWL2biwOfxdJ59k8sMNBwOUypn8
J5tGZqXDp3EUHVTQg2KDGYkPQqtEK0eZYcZO62ZhSg7qh3K9/SYOKwpjLL1wlqTe
u/3Zqyv2M+OcKJwzWqVLzAGQ2+x68NQ2rrodTbp2LKUqh6pJ3RHtFXCeyN4JMBQb
evRhlCvcHXxjQOODNBiqNFnArCZgn0GyzYHDOXSbBLQsdbrHEc0m7k4FRLYnFvD0
jaBZFi5P7xhNoOZWdVMUv/+8EDCO7kehAlKrhwbhIQNlA39YX3FheYojLZ3STGIS
N6NR+LJjQTBioLPmuEf8yUuVymRLgvNQNCLjZcP2CbALpzQQuWVOdgrzKYqNcP1j
U3lOZSIlHY6va8u3AThgs3Z5Z8M1jqFaCj6IFXV5Tk1k6LaEEARrmlTmafBKarZR
5yL5qSbTPz23esMm0LBwsvfXK3EmMO7a76p8XCUuqoktpaSE/Pep5wYG3ObGRB+R
FEztrU86RwkZpLwaILbAKA3IVFgwcqCYMtqKXaRcsxuWt/tQCl/PRof1eIVd7GJg
hfVgG7JX0mnPo5uXbCBoyZ4esDvEQodx+fwRjtYnW1ehtB5rERk1hsyMOtGOw1UD
V0dSwXV4C8YdUdqpDLsCLwrFno7qYu/Qxt6Ce931MoGrR4BtucDAvjEESt30aG2m
ZZOjcBEt4xgHGJFXiuDcRZV/rWM2ULMkyG8HS7q8LNLUApHX8EAsj8AEFEq2Dbgk
XnpkcWP6TrxpwC1HRG87NZPPMBqwhMhkUFi86vXvRi1qsLFxCbJuTSWvVxopmOhs
dFtAgn8Bib2oOpgwcBUIKhSZJ/4GsdC2n5H1FYDtQShsgwA+cqHL5oBd5I4QScu1
ycHF3U6BJXuNlh5QY/6I7LRbzDesKQI/Ko+fH2w9aKZEIgv7U1FAiFLEhhNLF7Bf
1uJvkxoqs+8FixVxiI9lbgIFM+IFLGCOQmXTJDmhg3Le8BKfEONh6yKXNSpwkW8f
zaz27/CCyyrTeyeS29ha0v+eF3I+mqgwpkEJI6uwOEl4WfZufScv4hdC3KvNJrye
L0xUCmavfRITaqD70vh8ZmLLpzgDHs2XQkBa0lMyqImZT9ErHnBtH1ufJkhw5SEV
TWd1gvmbM0i20ztkVxKj9S3aGoygHndlovjA3ipTVKKZpePc4CfE1oYvy2xR5pdO
EJ8F6VxzeNXTcv1VPTTM+12aUv0BehFarHx05X/w+KPFka8/WIMkJzGbFS4KWs0d
arjznD+4p30Gs82N7rKlXHHCv5Dko42XUmMtMHs5g/rUgxNkytuoDBFeznwjoIK7
9N31Kq8+0x15oRGcjHheYSg3ConZoSuXnn1H03NsZTmObAgIDPNu1qAArR1AGyD9
C2DOBnFOpCIjXJOtDEdxe/wkDnPnKTV9Lkt4WyoFkmWw941QhcyRoMAIV/ox0tvu
UCil3rPZTl/7BEliPWj7ipXjRyOcIoimtd3/E4sLgM2QG8eHuBx+weA8ARFHPQFZ
wCb7DBCZ9m/Yv4yUDdj3OBIcgrLnRiHOueXblhcdxcDTZka2DTfilGzfJDMkcv6c
TCC1U9/pDFjWY4Vb8EksPr5NcoimdWPvjeLjNFqhq6q8BhgZrmImON7noGbBRwHZ
HpAqPU0Sqmunuz6v6HSp79rRvYuUUogG5uoS/D2hkYt3IMOpd6ptZWbYdERLlp5c
XjCpyluQmRlgZzSg4DHm6idfOfdllFGRi7NT2s1GKXwyqssQvXp9DMjCwZVZY3eb
yNTrOgmo5vTdOH3BSWZfTffepH/GkuO/vGqV3YHBdpJ1WxdYlsWHHmv6zzQ2By5P
YpBUtQhMHbRA84i4a7CvBjFZ+AXJU7mXChwMa+NOph81IwXr/zyfSD2MwVvy6vdi
S8x1CtDlfI+tvUIwFGjfw2BkIFvIdZupM6w0CKUHcx8HtmtVayCOcY/SAem//4Dh
MUYz9fOjPig6RZezM5NWHvmY32LrL6OE7glVQyGg9fCcSfs5kBwSpVSXUCtvDJaO
astn83zVz0rYuzz3tSuoMEuiqSNI8VRX6J5mcS5dpeebBZdnHowkztDhGJZmZzkP
+a5JuVmpO8Qv6l/9OcN2x/KMYBqcSyRbo8VNrJWA0PPe7PsShO7wv/v84eW59i2y
vneO9J4+jUkW5l1b0JpHFTVEdWVPDXmJXLIrS7etZQ5z0eZNJRtQjU3WO2TsLheX
mAf+JdQ23oWUH0CEDadZGTHUQYjqLqfQUWK+9OjbelV/S7Qw8n/esy5La0dONtm+
FMDjMw91d95EM4XwxLQnk0Z8Hv2HYvAwx3Bb5wGMy8Qf+ljyZlUTTV4yzH/rKTSr
QV0ISEuFciZofxKST4kku3O9kNc/zotE7bmPlVdMZaZ4ou8D902eyIX5CMUodvWT
X4QdCvezdTCeftqhyg/arxnocwnmeAt4HQGUJCbOQ2F0Fd/NrosuEpNVheUBHSC8
az8c5pxhUUvotgiSkYKFfLMEoGNuhpaHvgLY5VHS8nLxXO/9cqK0Y26pC7heyxvp
9AOsIGBqja8wQ+3kBGdSL3LtN46pQOuOM7HslIynQYnGgjl5OyRjSmvmZjQHHLa+
JqCIlQDE2vJ/VeohsBd2q44YjjgS3BioTOORBvW/p+n/SMuPQpKlBUdXRr5zKL60
0uwElywM5jxmGHGcTLfJr1/Ce64Ri3cnesnv0njPWn3sA3MR5C4W5ycFTHTEDzaT
cezaMwwoFz4NUBPjbMUC586ADKMriIDryUWIzB6RLPZAvRzvaRjSMtcsHMRNtlql
heU8UC0NKvly4hzhK4pMmM8VKHKtxkC2YP8yCyfAp3x77srjNsgKemGtlVYEVMfz
NOj6NVhu3F/7KFtSDJsoPLrtAcs9PmZGZrRSFZ/eDCXppxWzZ4iMulZZhG/Pi1SE
eh/4Et6i5ZKuyfmVPqKcXeGViTz+9ZIUP7PqASoE8iYtZia/Bj7E2OAlCl+fT+pq
Qm1iRkRjqyYGrG7ZKo3qfxxR1RIMwj0VFYbS2PP8O/BlKI7+qCRWS0dUVQugyE1X
vA5pWIfNdiQx3suKvXGowHNSjyMX3aIPRhyTNB+KymL6fD5sagkI3aZrRfpMwdW3
Pj0tmhwtiubblUUoA8V9GjsIfVoI+9qF9DthlQSlTJ+GHTLvhQDZLoFwdIAifkNu
bfn0dl0To4mNHF8WSto7OH9ZWTCtgbkALWmiT9hx/nG79f60ZolQIyfH2gkIzVIy
8fSm4QxNIOLPx2feXe8nvhLjQdwE7cYIwb4tTKmA8rEsw/I4ERtgkBjv/27RtVie
KcvK3yZZTPxR/ZiK8FmauDCTUXtuBokPv6oqaIXeUPNfsq1T/7cf1govS4DaSsfM
SfbGf27csT4AzLUXJMhmkI1BxSkmiHRB/vR78Kwe8PDr8Mgdeu6RXzmSJUFDpejL
KbWqaBgFQqpyLyEXVdexfycNQN/j3U9xP54ZJEFbf7ZFb9kTjB8boTtSq9ThiEtU
IcLEDou2dADxdnQ599FRX4ap6hjR08P+70wGFvXUjEfJYb3L1BhBmq6vrTnNuoaE
qTxlwxvDfJrg0J/1a8NmrLO+/91rYUwNii9553Q2ROEU80EZzHcDtDNSan5qaTTd
rQvPGcmtw4dbRZZT8Ptq1ufusoJtLDFL0fvVBGTml2He8d5LoaVRJrXLJKSAOn8T
xeugwiwumJV59danh4LY19s7a1c5FDLRI1B/UlgvQx11s4aGvJntd7Pa+tuQ8gQh
tKjMqjo8Vd2QWsmYrkEPo54ayqIbNVZtx14gqk3DRVxElZBetQPJUSJ0JvEVCeWF
9nRLBfslg6W0gjOkqkPib0plzBuIkiiG3Ffs1ax4WmrgMpfZ3eD3mfFDjaIgWM0r
d0IuSHgnDRd8hiJfiIDwhGykT8G71qyPVKiIwiJo6RfDBiEGUhZic10PHc4ZnUeo
3uDDGS7kdDIgD8Vgdarzs2gRTbP0sWpUjmKgcjQfAWrAZtpSzlv3A52pQS63SSUL
b3kfQnhRwGkSHqFGq3XEnKXG2YMepjz38QT+WmsZkL3mit2Af8VgX7mgqvCNbAJe
JX/2n7AYWgyMeDCYji+DhHp4VxG+abVZPavzLvltJpjObBwIWwUZTnCe/jc6wxN2
YmErgyRPaiRgwnJ4W40aHM8L7u9FjSJC3ApDHbIBRPt/JNuwmBP5O2O3WF/Jyn1T
2YMoH0apCvfgbpSIsrdaP6SMBnTBtYHvYnKRWcipLmB5IApjQjCigr0nWvYIte9b
Ht+5ksyNEF+vT9knttetLjAbIEqQXpdlf7hEuI5l7Zgz+PCV448aaeeb+irW3j1f
TWtzQsVDFROcou5BOITo7shMvHaLqE3m3y68RyHWpxerwbCW358rVi0UP7uMpWdW
1IJS5ZVPzFQL/WNL62nHS3d4/P0lptn+61jdt9AnQ0GK/1KnkKlHOnYwBOi9Pj5Z
6dQtCK9Lxk0d3EiGVH7rpirJ4H12ffcgTS1yT7sYCA3IaC1m7ciJ7WPoYlSVykad
gWt7cShlImwwaktEGUne0XZj7Bmk7EtjC0zI0iu0rSfk7hptDIijedgZ0wi2wRfc
9uJL8/hDIXGvVUQGld8SL8NXu/J5uyqk1g9sGAW4b5nys0ZWtg3ms96N5ccNC5vY
ayUFf0OqFuxKNyxaRad6qV3WOwUfn/uNbWDTps3mMi4FIHxWi9Z9K9aEyTS36E2t
I2nOz4tElTGj7/PDq0OOP+Df1YmqlQ/ihuIpMM7vBl1zd07fLfbVBwkLFH7kEvxX
QBmyfPWN3O92SDr7RfaMmpxWfCivzfrPiKvUjj9N33BUjCp045YrSKq4kAO5cRhc
lNsWGwvUFfMaJZpmkA4Nrd/QbvXx7Rq25MfajSjZrgBnnFMXp0xcVOJ6WkabTYjz
YYIKhOdXe2vjI0TAecm6iriWi9RU/F6DrQ7oEfFE/LspORuCLwFKQOdBWtHRSnte
+ZKEO/XQAPo/HPXlz+WBS80qc+hYa3Wx8QljHqp/c4KLT9898yLGJqVHUZ7SFH9o
/uf+R7B/1KNfr/Pj0EqfdiEBV9uh0nZgssqo+I5WQWwGxfBKGGmliKPgDUqu4cB+
+uu3qH8qNd+O6gyOwEw2LwqhDQr4hKJHHJoVZ/L7FK4g4WWd6geJsriNqttBaah0
EWDzYO0tPlZ+zf3uBJ0LFiZz5+MJ75PVWHpUKLEOIGDJL68hhSIgrLGM7M4jQw0e
UF7f2ySEfZklEYHj30/1ae0SqGs6Iu+Of+vdMRyWt01kB61RiH2vfZScWqvkNfRU
vsdGb7AkgXIQiQ/RsT3bU2l37lpraVthm8yac50FM8ljA2QD2BnmbHEXddos6Ser
bDg9A7W3QsuJug22k1dg179pSkfZfi5Wddz9vnNn0bC4I9pA/rDLBS14OfSs3A0n
gHkH0u9kwRGuFEkLfWyqXftFAjvJgMz7XMBvH8WX6tSPDeNnbztFB/DTnse1CfuL
0AisNKlgVKTID8y+145pdV57wYyYSqLp7YTgd4IZaELpaoxOH11m/r1JPaflxbpI
TD3bVjJ6gzKc47qiaz/msPNgl7goh83GOzf25bp5YTwBPb/CfumMdj6pvANCy3Fe
FOLaySUM1w5Vtk06NJ/AZyuhOh2YNkVqEBzDIclYCdCXhyYXr6jhNzKLkQiHBOkI
Gh4vIF71yn5vKNz7PHYrRmMm8AGlLMXSi4hZEC3HNydO2jBIpfZemOTcYl64exUm
wHUxxmhSDEVfYHT9yZomAGKd13Z2uE1iXqcFpVU5uBgfJWDyX/MW3pf/hHujWe6u
d9mTyTmgyrT+aidrqVPssWBHmmy4ROzH7P5PWan9zMWR1leJ9k1IDPSsNpjXCdx5
lzoDsdbTKDoCHxscCvuiqKiLH/+YhKSt/Q7FytWdXghyn9kCxlUQyS2CAOO3bXsp
PnKFjbN0osYq7ClGN8CXPzBzMp3IJ/chcQuXqfs6G9ULFPLQaV27GjdiQmXeuswI
iqq1jPZdQk714Oz8VhZrCDClr7HY+NjhkKhmdTKjCp/icrVDDaBvUPMkjjdBb2bl
TqcJsBC+lU9bkaxPSVNYbXQZX2YGyBZL93txIDBlGmiAikvCMClWsyw+PDjaixjv
27oUn1iYS+IjeIg8ig0rPY4h46GVNynD6WpVJAuL1SZ8wDxWp5RfPm14eHYQuuU4
4Xd7iq93pSpOKXs4Tz7calSgHGlY5sgP81RU/DvP4yncK9NTMy6q6bQXa5LSjr16
2ZQLFiir+zSfefGXzCUMVi4qi7ketHwy1ATTrRoY4X5Y4emQCrqWB0h+u4Wu25ig
+zuwJUireQnTWSMNohOTHq2/2J59/yz18ed9RnvdjMn0YFu/pHCZs4WK4iPQLrWy
5fvGxIVF/DEdxmM08BH7amdULhMv1/84w08/NFdSNkyboHwj3g7w44msE/+Zkw+F
czGD8vXg2e9KeTOVrMrWWdItPfUXjZn+uRvCyUTxRkWs6XiglNBa6dgKxdAaQeUr
nsNS2I/HLgErUmF4/zoER8L03jXVD/uPERF77FGHx30I4iL/A8xKne/3SdAAmM0o
QtmaqABgFp+mVjFWlIrwj9/dGqy1SsT/Npr/QdLfscuJEZr+w+kCpnWW+2muIv8B
TVbG+OTL74Zkg/ocG98t7hqliNFF0Rb5wV4YB2mX4LLX1gHOrx32Jd4AsK5O2Emi
r/fbGowEdkg8ED8vOByMANKaAphCRKiyhzFKHdxlDMI1TBVIoQa131iVS21L3NPU
5Z3b4H6AT0ShEueseRkyLOv1SJPTxkoU3lNO8bk/hqjLlmVQxoF94WwcTbMIMd10
sY+5zUL9FYssGaOaOdP5mh4z63Y89LIZWe2TSvdMGzJ6+9FfaJpxOEcxkTki/kSx
gdJVrgYXZWsFGLO9C1Z7Smx9X0q0OdXH8EbxKKlQbaWbT5zvD5ltelkBd40kPUBM
pOsAScyJt9vpUY3ThLMY5NQsrl/sq6eyFs++PlYeNe795CRe+39a72Q1EBkf7oeN
sEjI2W0IX65kxtv2jmfFtC1emYcZZoh6VebAs0qUeUBpmjgkei2r3A5InlcN4lKq
tvoRXSMAKSRDdFrPIWVeG9A9F0W/psGlDB6/XMpFia47Udpgs+r1ZVxf2Un0k58k
8tdkMkfe9iZ0Lw5//6FOcWeJj8GRhIkzEPULIRgqj0sg341NEivd48CfVw+qlkSR
dPSPxT/JwxZtSvfur6kftslk6ftfBM4wgizI6Wrzm7XU7Kz90knrPeW41ZhK34XF
5eTnMFo06j7SS0gd22vPY1RmWk/5In9d/rDqIYthgUYMt8K9j2RAx0MG1PGjZnZn
BjMHFEyCQPEuOY2c1qd+qcTseef/YHK8v1yo9lQGhoqINpVFcnQNtD6OJ2JD8lp+
QWZo15Sd0WsNVnXvdCUyarqcrVF2BFwzFFVL9f3GemO4FSMy7yqadZAqa1lFyyDM
jb+DiNCnyqxS07AUA/SzN04dS4qteLgBv9G2pp+5X7SPEJDFPeIDBBEo3cPRJIjT
qt7ERVAbGaWDtIx/HbbDFzeBmD13CH0hJZ96FT9KCq+zHRD77cFie6CAvq3n6fQ5
iXGPI91P3YS/iENHCAC/ebHixkYWsmg0gMHbQZoM4f3M5xj6BKRNSZHCWggClHbs
65r2v0Y3I2/2qm6n0HMds0YR2e3VtZwTGt/daX3N2mQnlAbVNG6rFSx4EI0Dr2zm
YoNBE7J6X2ET0Ia1jJDPp7dF92oVhTvJR+oY4ZtMHTsyeTQoA0rxJdFO9jrWd5Vi
zEb8wlrRTcGPCkSirsN6doQzeiePThefOrNrd4rOjGn4JMh5IimNWg4RcbYTw/R+
2eDdJy6MCwEEPj7w30t9wunC3HNS6zqYfdTTVzYxSrioVMwx+TOD7sRugwXX+Xuf
LJwWAxSKbose04jXNP0p8ClrlEKAM+qMq+2qBX0yoSAlrbzuJAbhfamJopRM0Kyb
yexq67lvP3/112CpnULFatDu+014SeNwBciR/MOIjB8p0+zaINZociyocrojNit2
jiHhAhGK0rW34A5m4BKpP0Tya+1Qy1DYqtxb8aAdEqM9ojjiZM7FCKXh+v0V3VPh
NuKca+Jm3q6I3Fxa8q51xHE1CZsSBxzWIot07s0iZIWa+gPxxUhku/7b3PyYI5tI
6Gn1d3MRjJO2x0JEpnkxyg0iHx+9EgCmKyYyovcsrP0ZiSEJy6bR/MUsA9Bce1+a
bX5m8Mysc2NbBYpl8r7+9pgnCPd8JPZvoanXsy6NMDVTSXaOM+9eOWBRNYFa5y0x
5Xv6N6c5IjOxCUpeLjwyQW1CnzjFC0aWHQTzBxN9cqah/gIXqgUuAT3jBBf6pUBn
tf4ZpzP+mY/OfLMk1EZ9ATGvRu8zESEDoB1z6ccw3j9x3gx3galt7UU1Lmg83Eab
QuIh6ziMBhImNX6Xbqx7MW27/5SLzntmiNkbVTFBsC0mqGCGHB/wfBXHG1Oy7LIE
IFh0hjXZ+BzTHrzbsIvAPl4+MUZNjal7dp++z43xc8iGWz8YCucZNHSTVlVJksK8
aWrD3qq6w2S010exFr+ZmJs3jK9ZgIpDUjFA3u78MEwYqiN8xc6nKihhi0mPjAzF
wh+3a53B1+V/yw9rq6hlxbECpj01tATNHBoh5/+IQINQCeIjP3LzRJ+L+c6V7F7B
hPDVl9OYSge3pkUH7Yt7GyerBD0jWNOuqLpL4ED4XtZQrqg/bGP9xqLy2yKKreQe
wurf8mQK9blvGWVrIDwsPrL5b5N8Kym4oZrM9PD4ZI00Gd/vksa25pEiwyd8OJ70
Jrw3O/HUGQC/wRD0vqnKXjm+xxOYZzBJthUvDcUE0YtQFZmQ2yZN6IjB3XqTiT2E
lJL0z7CVQBN84OePhkDfN+T9yKIuw7hgIpaDPfMQ6EgZt7oofOl2lZUt1HsRu8SS
e8Cwp2mLOdjZD3f/VPXGUICM7kBaGlqurgN3gVhPUJ1gVNfCV0GgIWRjohwOSjZL
ZZ5nXrW8/yiwvgVbkue9ybFisE7URYRqxTh9Gw4drmxtlfZ0IpxJpoaYDbqMD1DZ
xAvkiKsQXK64WTZIOgr3mJZAvrTkGaZv5jVn+JHODMD8DNOPwFlUORPsUlXFqZzA
nsld+uo7GpEVu1x2Q1ecHDdoMoRj2Y2EdKpXe27SMd8vCiqCKwS+GfPCtXmosIYg
BofNOZsaOGQqaxBVI252BmqcM++bm20jFYvzbSyTp114arR7JTxLUYiW/Y7X0Np3
R7LtwGZsOMVNmBzESMfJuQZXoL7FImZgJT+0CbHOiCosfVckmme0XFl5VKNEElnK
ZS8yFZYPsYLtxhfSyFPRPPPQBt/VeXk/tmdAm1UydihdkVyX6ueAv40QPTWeXLqd
QKnoI8JeO8H9GMHZjpVZ3+4rKeNQqKVuP4hqDirJ6kDfie5FWgduOvn/747QLZSx
12XeDuAbzuKKyhMkVmUxt2l8YlhwSB/MDBzBryvvmktSWnoua6nmAu9sH/8PZyXO
dcqjAsK7rOZpUzXTPnKu8ckfaTcByqvHXsoROYO/PLDmtpdMmMbVj94jDIaMRb6u
nIj/bha5h24hGhDIQBndXZM8ffUN6Ec1Grxiuw6CkFx+MOtiWhGOj0rYeOoZGwT9
ICbbpttXbZo/gr0ldB0VCGFQeMSMaIDDWcXT+4k2EaDYdKhiaFDadlbT87dAcdGq
BR4MQp9zoVUXWVJEEEjhRqdQICkID2yqmq28E6fIpkts3jD6cVTHhGnZxB3bPPHC
B9XsIEyKDVRNHs3ixdOzCRFioRG7x3b4ef/QryHOv4dyWl8Weizl0kAu2SsELo/Q
0lEpup1g6DWgQo1R3v0z47Py6CvRfL6oBcy20p+OHUQ/OUr6gCWoB/StAg8AsuHm
siCom1rekIpC4aj4ubWdyjgclEl/Zzzl33TXvW0Ah128RpKMHwgj3W5CEWjzAbn2
xCqbg2g7//zDYTIpEdE7NJpVak6Xbd2DGa/JQ9rtkopMHSZOiWfGhqmup+clmTOS
xLIR5xHzTnmZYsdaXcJ8gsp31Zcwa7JATktAbOROiXb5qqUE1qN3dPPFcm4CiDw8
pB2jB/UWK3mSOITqHa6nX9HdFxe9V/vEOaxVV/j4K9s6iMiLwoY76wVCL0JSyCha
+aY21wW8m63qrFILh2gEE5AjZfC72Ud38lucYm2xtsDt45qi7pb+a67HG+Yw8DSd
yiROoFxVrjrQ1K8N1KXgOU1/CWKzEciiuAZrByuXkPpKAX5037h3dozakAw1ElSh
PNbBOrueuhl9my3AhHPcP0ppV3ecmOom8F55fB21KgAtZMdEiYu/mRj9/EnVqcAB
qbogTE4RpNuCsU5pXvTrpZIaj91XwD1AGCWwuf6nrbfa/Sh6a3LXr/GjMkLI4gTq
we5IUevyibKDkTiEDrXCPQzzqvrDi7zQbZ5fi8RwyDKJDKyjQprxnNGhsAkBlXs9
DxgdeeqYvesdnDZx4UXSWBNBkNS7+h2SpJC91hyJTYsHVMUysOVnsbdvhhYQT8tA
4Lh2FpG+4JgoPcw5xoVXJGrSEWnujLlscTJcen2Bp4YFlizSw4LBuXMtsQ9ZIiAv
bZWyqFpLvE4sKq25aQKcZ9cRWezy3GtUZQRtqgT1RDWRBtXolcNRFQaY/6Y0YsB4
8UA8EcgpIkXMN/m0/JTsn8YsznKtSEmT0pVmfJwgSgXZ9AAmLMzSN+gD2Wno1EUT
ok35/4AXoY9DP6c0tLRlDCFkmHlzmI7OrVkWdZ6mvRKKb8uTkhpimAmz4i4NZREL
mDwwy3peC8RUc/F2nv4XbgfUHxoAmyEuKJiZaIg/c/OoCV/1uVeL16dcegbG3Qdc
PmRxtRySm9rUTG4yZ5A6mOp+TrGw4yltvq2GP2VHhIhAZMAJT8t9AUCZ9lDDaA+Q
xheORW24me+5mxtDZnxHl2vblxs6VUiq83+Yq+saBd6jD3SM91tfgxkl8dQo4Cba
FBd8AGj3MmLMOS0dyFCFQUWYx7P+zCpba2eOQE3bNSs/buj1yKGDUC5VkJ9XEls/
trOZjxgeg+CsQte2CwhYpqKx/emW56X7oUyRdkSo2XxZ1wWok/+FLA/fE45lysT0
T2MvdF2sV7o8UZqp0ZxjwsfyQuFDwaWU5is7sAVmarYP2q7sP1/DGq8HJJKOofEc
DsRIEKvaESphr4Aky2sve8Sk9B9D/z53S+2UD8rhud68QplAu4KCGU0V+9Ckw3+5
rVA4V8OYb5/y75g5jSzSjLbmoHPGIAn5VpiXSHjQ9AYCTSH5vjJTo7iBbQdYmEd5
CqCItQODYTxHcsIPYXUwEYXeBlhZ3UpOZdsy99Hb4rFm/W292rCCC6OwKOxABVXY
NoTqM+LDbpTdbVZniMpnKo6tw61E2EHLJnkiG/Qgea/uun44ZUJbuOY87sDR++uL
BhuamkqkiYbDMH3m3KdTrZrUp65TUFu8Cpny7vocoUFEIKUuiu+CT8TgWZm0yv+w
NTjvsRy9SAEaoCvDFWIyCXXFHSog+pLqswZxfv69WoZDb1hxU7dqyZqnY0NMMsnj
PDf3vFqKqF8R92WnOSCECo/tsO3mkcMQ2okxOIYgE2HNTEh8E5MT4FQYAC1d7rRA
C2UA7f93DmUa+9CQmXDWNu99Hmcl744R+ei0aIIzCKSej/hVpsg2cA2zHOK2BLzy
SgPSEtPeNgNrmeJxccqUKkz+pBGmlx+zmPGhIhRW8JNJDuBO9zHS3u+W27np6lMg
z39GNWIKAME5y9Kq28Djq1LC/Q3o+eY4tyEjY/WDrMPNBqaH5kWomHDwPH628RbX
SN9s1lZ+UYInDYYCAuUM/hwFh7ZcKkXoDYfo9pr9mfsNdUUL6tGJNcPM5NhgYktD
k7UbpKWbIKUp6qa+sDSJwjWuvCUirRUupQFc59a3JC6gacHos0JRv8GG41kOZ1De
Y6aj+CLUyTXffYXjbj9/DAqw3GMNp0HVuoTtk7sqoCj/IlmZkAUHU1rA/hNJdXVm
9TFjLf+20ZIeUAUkWa7zurz2XNzEarQ/PMeTT3isSjOu/jjTSaLiCxbgb7rTeVnB
b+BLTz/nrp/Tc7WHpb0iwhzY56z/8jzoaDPEvXp3Hx6w0GK9Jiu/kx5Rrmvwvyig
crX2m+orKz2rPUeKB1aS0heV1CLtVGOctUhbEo+/yodF99PWcYmYQ7BmYjGfDaC9
LtSTjHtA6C2i9TU+5+cTHerGLWvi+Sarx/ZT0hsFhC5oAyixBaKjwJ2QuRGMjTxw
dd+a277PFFTESz9HcKYXJQ1tLvKw9+RP6tm8+9rBPnF1SaZ77Oi6WiKTFnyVuloB
ALyF3+NfQCzvSRRB56TREKdTDKOU6/MXOmRhHPrS26pF5jwJwGimCftyemsYmV0f
Rugg4d7/f7+6gtZx1F75HbL554kArDNpAj4ULgAeU3cr4B6xARO3XtqTOT6ZxBEL
zjuPFXjPCvFo9EFqwoVjxHYEwlOpzcWhzFS3qQ2J0tx8xTY3fthSzorFJ9FCV/ZE
283F2mi9W2f69TM9zljIka8DA1amcHxejWIIoSxDrJGc7nYrO2+xhsWaoXu56yln
f7RET6rGRZO7R6L9gp5VKW++YxU6XOuPyHCyfnJSBRtgXCM6cN2TX/xcTSCQxrNS
uc/y0qyuT1tzHxozQo50U3QxsSWBn9R4tvVvZf/EmzYZZ5ikNj324ahEzYJ8LvZv
cOOwYApJE2JLBiMbWI1tTUJhWfdnuSqKB6JcTKwaQibBc06WFxcvVR6OmOv9y+6i
y4EXGjsHRUicE57Ld7Csg42ghcL9tLbIZl4IP3C7JdxPilmdFlvStASuNOcMzXCU
gy18gmLOMbQukgFIN62Ag8riBlmysCgeptN4vHu0NF8fGdTp7uIAI78SK3QANYxa
R9FlxAlRxPIxITO5gk66AAQbgQdTEqNBWdE3oGLfzVfyghv1XwTlWjHEnFwGkhLY
eU189hIojo1iY+kR+saxcX/AyHQ1+INeC4dLABY8QvVZuwNGZ3h3eiGFAbbeEaFh
/PVfvmwqQwv8TXYhyCD6SgTILg7UdGKE+WsQ2uP0uXXFn/Tc6N8vp1iLN7RmN1KO
hM0GDl74edQwKdYBIWMMps+a3pLU8kFvzNOmWv2mTxX5T4QDzfIfFAzEux+Fy4l3
zLUXvFjOWFRW7JC8VEBVnk3nDTgMUrqw2fJk5Tvouf/+L6Sru2GLZ2Q8TMvcpcT1
aLmhDXSIK9I43qZulB24eQpCTfKQvs8DdVTpTsJFdjTzfxwNXf4kL4xTCeOd4mYU
Scy6hAViy9YcajND3C/sMiTI78kZ7WhE0qi2a/s3pSTOmBRhnoUjYSrtydRFFDOW
PM/HHm3sgXnNnS/TgkZy7p5JhYuPEFdSyda8uTAOLcCFtp1ynybXPPacccRsKAJD
/iUuald6RVqaKsi42BCFztgtVO3S8NVpvJpcZXj1bRZJ5la1GqzI33RfLN7mGOoZ
waUuqsnvnsq/Rgo33de5rY+Cso/K2PGUsfe8wLHwx34BDyPtqIwcSXDGUnP5fpj2
bf8AI+B+9BeRkRz9fPdmL+7aQogwx+LxczNXT7P4cf06kG6c3qF2aSI9ns3HtEHA
iZueTkdJHmWt7leLUL5QnEP5bL09u7ehbVwv/MC/oRA9ZUulTMJe0AMrg2F+HHfz
33ZrJstgFAMgELjv8s9qyiJq7jZR86BybxYevipnPwxH4GiP/hVG38PXriWDk+7N
US0YcuEDU9BezoCSzVCx80RdkF7Altuly5k+B0L54Edl24deqZy49J2szmQ/4X9x
jqJpaokyzqFjnj+Ir2h0+yADQwHDoHV2toXIKRI/OrOOr/NNJZPbLmQ20fIUsm+s
EEKMIYy9zAaWfePSEqNlwweG/Q9DX56L7BDKTNgU2j6hH4I7x3RuJENauVZv+I5K
McdcmVXDMmQrJSsbdExguRCkkMKUiIKAmC7cPe1QOUrqp3NRXD6YjL8oD/W8OrZl
eBertyOLYHrggMv5ljFIoKbAuf5MH64vd5g5PuSEtSXUIAlyHUX2rVjblfnWdse7
ZfVtQkSjDsfRvlMY8YCvi9yi6HgRbly9Dnvl7zrqbKRPjoDg4Wqp9m4GLao8qrdE
GMMRAOBI5qTPu/CgFSDHaD/qpTQbZ/Y1fiexHGWMO7xbzmJ5Sx2j+XtEU/h/BdtD
C/HbYZV8zNklLWsj8Q8bhUDMybZp37HyPnXjlMVDrSv6mTXBtIWwq6dQBf7sOpvL
ln/S42FRynkIT8SEl0oMNBb6D0n9erZm4DTKymRtpUZ6z4LAluBopm4V2kA3LSPD
KY2Wqx09Aqa80/PdR5JsS31h5RDM2hQV55Kf5V0/wPlV0GU3g7BBCVx4H7W9CINZ
yhbfUUfcY3bdugjNdb41yk2LAB9R8xMqo9wjFQiusGCVGHZS9Xbd6KgIhWeco4qx
iIKFjcVX9TCI1kQhBmt0nY8xu+K3frghC13CRUcTjmdhX9cakMpLk+u3oLt+pPgk
AmsYfSwGaAhBKZDaadp1fHXneJHlwezEtIH5rWeyZ6c6udNV48zRXuEKZ2+7e5A6
p978Ho6mCZQW7sBDME0aNsyAA2UR7AIF3629thobGkySEE984gPszuTrwvGAB5Vl
qzJkKh3hIoersXdamCR6iIeGLyswihnozj56EBmfT0oz7SXtn1qUERE9Opuu/MeZ
4slMCmybUKArdnCpDzencXWoWj1zXILDIkHautOMYOTAQvo/2IPxkP39o9zZb7Zk
QZP+yJ3LqY+TD+/zbIB0Fp+zILmTXO5GZEZBq1CWLFBerTo3rbZVofT0NEJm1bld
WHA2OLPUtcoboHTuZ32b4ZrpnpwukKFLkcu1tfmQD7Qahq9IO4Vu6ebYbfJtqv0O
MtpNIX1TT2xDkqq16gl1dgKuXSaI3E0DIUOqFhyJsa6eP2+M0TI/i7jSbrxcA4Ck
tEoPQVeQL0ZhbI22MnR8Zu4QxgBIauoBSc4V6T7urGWrXEGTzq0ysvGKu4HmwqIR
mEsCuqRtg8srrxGvWXw57NciRwOgw6sWpPBxb4T8sE0WCLayeid0qQRIOtN1li0H
fGtqw/fCxtU7eAGCfaQq+0V6T3wKMs7NSfD7VTVC2gwXsA7mnVmF57WRZgRh4XDa
qYDn44XyPDP4eI/aM9ecGIBxKSOQKomfva+BXX+rzi2Nvo0Kv/l9UqNp63Pbi3ev
/dkLPaXagaDv6aRf6l5jPfPr28XCx1OvD5LeRbU79678U2bRqAhW0OwmvWk9vVsq
/7JClNKzRiqBGPH4Wbce1B/hRT23mg5xF5hTyCYbCHgrdOxg1F4vKrpsfB921zUS
D7TG67QmLKwhH6m6WCPoPB105xwcfcSx4uqE6cih9S4QwPvgJH0rVV1wjbbUAW0m
SQqwzNr/uA3r8LNCMIi9Kj7vRv0kbE0gnEePSRT20FfMFrcxzYrS7fAFXzXgPChk
256KYXzEDNKb/zqG094WkGJ8mXy4TH9pZcc+dub4CbEZUA38tXo8U8RyCslWozw1
8l5c2aeLq4mM83ldxnEqx6A0wlZDOb2D8Hs0JjKHF0Acic0Hx/ZALB2VeEdWz6aI
n2kQcYDDSBqFNH/vKldxtMhBLDZpDuQgt+R0uKwDLhtgaIJovsZPRz1AEWhrL5Cw
DgAkKbd7vRu4pEqI2mnrz0OjkxjQg6rprfx3+3owICey9zjSY2Mcb32W61nfNW3B
8hDjN3gVLe+TPxjNfIi8xLWljBhOA+FIX0em368e4ztgPKynNwXfCIkHBu6Yo2lP
HWSDyHKyEZTs6ah1Q9f1JDBEJXQUCIlCBL7G8HSl8vkLWWzr2QUKeregPLDYoA93
BNUYjRZTB+T+ZFx4VOV7qAArRjkzhqmSQONWiE/bbHv1EG5+p1scABuAvUbhigSH
dqKQt9cCwPwcLj3HLYLlNs7smAWWrlBYfHbUCVXKSzUrH2W2YKgyjgtXQhiqjlkS
kXg3CtFxPnz4l5SbgZN4Sx+M5JngvJboPPBxRQSpHA1wDMTNNLTlNpp+8qi7uH4X
wFwBpBdSxQ/8DxxCoByJEUiRG0y/ErkpCvWf6+6UgcC39Az5jeTSTmDVJsF4hQev
km04wFNr7QvramxyPWr1Y3RlZcTKB1eHP6c0QFtf/cP+PvCXe7Q8iDH8dtEpBVlr
8LZIpNghVLwADRaR+MvD8bmQN7NX/GaFIr+rz7sEDLm9VzyWPqeXYqdOW0Gkdnuk
7YJvFVKA9Z++XqHHFt/loszbtXSCW9W4HnX7ylMRtzotAvqO0erhZ+B3Iy+aejCv
ZAkEV+3t+PCNmwhEqU2VKZDepw9Mf3xK2IfQ+9GzKwwwPpsqm8ueZYlwZmoEMEeI
iDvWc38aAYKX4K8N2Vqu5XHCCO3D9JEtVGIAGGep+VGtYWgr8lEBRmUkZyB5rn1V
71t4cjYKKeZyCb0Gtet8RvkqQ/SJzaW1quBut3WSu3gd39y/2VxodRcz6/Rj8FCE
AQzGWK65PsWOUxZb2v1O9sDPTQ/PDWTzox9Nw2MxJ/d065ZotNt0FxLPcSYMhNi6
5nsqTWRLCGFdgRCQO485g4+IPHYVAQMYoi/k6GL7Og63f02LCVdZdm5oRTQ3WR9V
o3i9zLzcqo1k/iOuH2Lkm8NWOyWC/aZD/sTp5zb2mluuuowgElXN7LubDiqmtyEg
g5hj02l8yoqnyZlzy0bpDAHATHwMm1uiuyaUA3BPwUozvVmYqcQted+ocdBvO3o0
A+vo9+uFFQgCZkPE8tHl1rbUaULJVRsuqU/dw7XyxpwGMY+WzN/ju0aplwDgJla1
M8StiVc549ev1Y8MnIpVU6yEZDCV39Z34Zr2tEhtE2jciahXZwKrqRKm/ijCa3Xf
c3tQRqW0XsfFhmS6BM9TfEmAL896LptRmMHXkV0X5a5RuKOvbiTQHZNMrFucspfb
Vm+TpQcmbFGiWxQk3ZGM0SRL1ug0M7+9h5nnut9hza/k9+Mmusfh01GML38KD2Tv
YG5sm64GFSsEup2N2/FReTWYkbE+RThppvy8RLmsifAHhadwdlOczPZ5A9oTtpJL
R5pDtgLSuQLEBfpUAx8eqBfUuTED/Tq+zEcTsQWwRsB7NeDv1kfnzBVxxnilRl8N
789PofVBpxDRPWtTMfNY8j48zeJP79TOO5mrJVOXipzUQGMdTeUkIhEnT+8EdAIy
rne/SpJWnPxVHizp69EW3UR/cGiCyJ2Vm+W2uz3d2KeeVcx0gzX4QZUKaA75wovF
Y7pR9JeVplKH5vNwZCQjnUnDFz/3whJPoQ2Fl0sQNQa4vGXsaqdMmANTvbmSe2ID
+Jr49EK1y0uyaDtdO4b3TQVuxQ6hRMfxOLoN1XLxsCtImESbrooBwoFojsOW85UZ
oKcPAaswyPgDd8KZ70ODK3XCQauAbky5V+hNdzI7PjasOseYInW0pfDT6HvEeIKj
Btsz86EN1mcK+OM8f+9fKjQJBlLSgth0dZ483HCyiJCs1657ziRRsCBcf3tC5SUN
GlNk/gZvu0soL3yZox5M2NU+cvsWYlA5/1Y/OLpxjexNuHnTuR+sw2zCX17RC9VP
WUOefZphmOMmhOXAowmi7EG+c34Xll5fxL7c6Lsfi9sLtpuXIT1d+y7ZtFp0FmXS
H7dvYBFf4hWvkdbaRCTOaT4IEkt1G6S5yz14Gv0G1lS5e84Clt88rPdKTkj7K9eg
Zv0bfMC+rT0kmFadKFqIMSLfpbZVPu8YCpbhAy8OthnO/fgeRMI3EUFLHKdIg29T
elbbmxqbz+Hsgj2ZE13s7FgBykaTjYl5C1uBmiTUg55nkw10/gEApvEZnOD2lqPg
aLJ6l63xqjND1x8Zoa0QtBT0IlNKEzcK6EaNtZLATt0C3z5Hhtg0+xaesdNby/mN
zwaCujyl/+DqIj4lsZRFf5LToq5H08jVdBQdbsVybVs7j1kNiSJf5lLH5Cj/7d54
z1uz/bCz6aIRQ/CLIx13RvftehxfguctA9aIBcl97uA948UUWoWdD5U7AfLOM2uD
D/RFHHrFr2U8+tAGrFpARK2kwW2AxAZQhFb03lDHyv+RHSHbpU6a14laXMGVLWNO
Jih02zN9/DimNO6o+lCMo2pL5y0kW9DZP27hgrWEYho/5ALKuZpapgjqgtuTozHf
1qpg7Lj1GB7DdqSIHMwypd0oUv3T7gcrR6zxNWDFYjN1h1Zb5lHg1B0qSo366/vz
wXobh+TsZq6GDWO7wxR4eJaITA4C9AP7jrMUxA1Y89uiqpX+32KhjBHSrubyW9o4
Yxb+CMGLeJVPi/U0yFoTDKTWl7d6q5hskVA3uBAawJ9NvoTh4gbBHrpz9nCzNFUb
Y6USTLtlNsd3/ubjGP8nbEYb1GpXBarWjAyaHpymXxd3Ae24dklc83tPjkmtB4zi
Q8YEr0WNktM2dlkACmbI2/KZtdqSv9iWjNww5M8VfMcoFvMygJTFXXk9Jhea97+f
omAAGhyMVWuAnK83z4GBUSMnw/EZ8JbMtmO+NVKlL8s50VhE+IRPDPcvtE7XUykI
4QHsP0S5dbgx5IZXDOY5Jsa+gNLRJQntKJ/OVmDBx4gk3oZvf1HMhPiaBUPb9nC7
FO7eBDxRR3750umqiMMJqBAAyhgnHo6wusSvplaf/1fWcvlGX8O8dIgXdqtl0mvX
di/o59Y7BjNvlI76C2NRYajHJOKWOxUu9VjX3UCzrHyO8g03jkSIBhK0wu08pVMS
omB+qKs5zHESHXM8fc+frI1NVBJzRd8s/yInLoDx8U9G8rkWpenDSY8Qs7X4Ufz/
e3o04ObT05GryYIBR1mLT6A8tzG5woZtM4UpkugZZXhutR6LWkZNLmen1oJSrkC/
MHwEU1gOOMnnyqiG+J4kBzW4M1ckxTkBY4FDIn2ut42zn96zxPeY4t6uIFeXk7tP
nqDnRLkkEylOUSUUXQY4Rn2sBVV5rFfrLNkpSVHlbC7oe9DQdz9eQpLbxgu7VDqx
FqpnLL9CMxkzHpyg/UyRNKSX2uG2nCeNiThE9oSsGEanKxgKSQr1wjiunBjEIkr7
x2PI3LhVfgs/qR2k/QWgK/lnjuHAAimxcy3rZRvBdXbR4fZ+yj/sqGTU3kExc5qZ
Zywvn8TJhf1NnyRVT+qdWiNXHrJF4dIYeXaSzu0KWgEgXsMd5web7h6o48PuapIN
G4VH55iXw9WxyJrk+uJhpWqySV/ehrgBbYEFa10hAJOafbXSnSOG+X58qvtems64
xVrcMipyDtEBULl7hDezlxSHl0c0GtmnEaRJP+tbpmGs//d2C1DinbvxQudVuYCP
JUKsGJ9e93Oww1mA4JsJH+rtUox6ORt6twktPBjdcHKVT8MAOti0RQMQd8ozDV7z
WaJn4EcvCl1RVbkzfCc4Hvn+ZJU8+rGhNURcYVrb8cJrC04nzJFoSqe8MjfCP+RI
5PbKQEclGlMq4a4TYt2UgbIOntVBaYEmnJj2Z//XE7oCbv6saN4Jks8ThKjQMEc2
ityyxiVO3WWCV11leRhOkLVprmswYiu8dJB7apO1MSq7Nx720kMlEH4j6k78kP5K
QVGcuyoNoWBHxKYNRU2GEe0pgxeYpeOdvH+N/x7EPhxs4uTAsNZla5SEFgLAheST
DzdoBa9t0VaIdm8QHF6K6+c9Nsrbtr71UcJfXEQ2SXNOAWOPjgguJDFGvR6ohasW
iBdhdIYjZh8nGLu8qikNBoxOZ+11Tw0k9oLjU8fI6byca3OklUHxkNjkO5Ilw6IM
u3xsPqXc9BZPwfubztvhviHOXMqfgxq0SEg3bswRLKAvIpPeumLDzQNZaSLx7PpL
Fw/LynR6ZT7IuWkdotcm4Jl+jZwwACP8YeXReXUItTgQtdtnNDOzT2o4u/JvSPM4
DCIuWcBaZVQiJBqDKIn7/k4/NsNFwbisJlbSXUjb2Kpi9ZiT+CQ3L4FRYmr4F4N9
CtJwZrLHGADfxAUYN3ZvkoYbn5TLYLq6DJx48BQMqYiEQbCOmAZWIougSiro4vtb
+rLXC2f/ngJnZZHhobH2qhdZZMs/iElJX18SwAWtCFIv/1t+6lGVOoRwnu0X2oRL
XSH1txjQO8UDdZfitJ7aCtv1pybDOzdUTyXPR00YiSVQu2mECjYOTSHk1Z0T9WEr
MDT0ilcCf1qEovNODZ3RNT3wH2e5rkN5B8xT/TPv6i/43X2avGOplTUEIr63xThA
yc1jP7Ou2T80itASqua6ybUMKeJVsvdK21AW8pkOMk6qusL9ZD4M3DkYM7H3SZhl
M5SANS+KneK0jbzDstclXQtBLKKMv3CeAo0XY6o54eJZdZMdwxpwAnz6v94kw8RH
kyRfPadTZejYx8mpiTGZAOzax0dwbPgxHhCjrlyC+Zs5zQhhIOJs1u6l1ArBZvNc
wAqEN9O6q8LlE3VLNokSJM09FC8XrUt6G7PWW3X3eYcBsOaowfAWWSl+GfmAykZv
DhUAErIfF7eyf7TPSKQ3EQJOo6OEldrPqBG6UR5+ETzkN0LP5ljh0muCmk5xohk9
2t4YliyevbQF9Ma64veDxILis+4j8jSmcqe1kWxyzIIhvRU8+/19DhweRHMrwTIC
xeusQSOxb7FI+cgzN0ctNS+kgANg3/HXPfJocd7iQ/z5FNdV/loOcbkmBcGHhPSZ
aPy9LPKB+HudZ0rM4xKDS8dlR63OFISz2+U68mtxjewJFCE+bm8vx5jsLgEjbnkC
qOqRJmA9GCfWV/iKjLY3P92N3CA08Oc0/AjF2FnbpNCrAh9JsXOSFmsoAX0l+Qcy
xVl8l/Br3hTgnun5k+eDzSURmCLG33lDca6fHaEs+/KK1LqYRMn8XCem5mC8DSzI
PkzfhqGQXm33Aim8KL4gdkOyPsSDNoroDMo25mrwlVJH9hu1d15/P3KzJ30SK0LS
5W59OUkXfSv0bmLF5U/sN9icX07+CcKN4yDd4uV2xtTqDjNL77fKgyg0qFKVNlv3
XwEYpDDjzm+05rSR0WtvSpMgjDDZdVJV5gg8mTCr8yCxCLnjfuCJNBmg+BsjuZ2q
9MyW10ibI80VhiOpmKhokLQtQzR8ZD7gGjE9gfCrEw/An3BXUsBMKCXmIqEsk8k5
aWJN4N4VC9swJPHY+Ve27OHSsdcRElmyUvZfA/2F/WQtJj+z89uDW4DU71GqF7sn
ej6vULvAt2FYxof9Lw1NWsK9F2kUvDZ45rJ+ydbodbMVO07xei7O3uL3QSWotE2u
qAI3jdiee7WhUCcsWlwv1aKpbO+sDUJjyhAtx21avxYBfBmnUIfOt0iP5koESRt7
X0KhiQSMghK9T1M7ixHewMRtDOp5aKK12ToKlHDJrT7MDWAT3WpxnMPr1FWwGc74
X+DlAzA1fDaFWiMrGeeAVOxNqyIBpxBqFXEUNTbiEfvPQiasRP2cK6QFK0TEgj/B
mc/1rzCBxdlXZ5pDBm07ooRXQ6g2+aKMxIDrZx6tGEjHrv/WpSfN4naSWbZTJ0Nm
O2BwDTWO49G2SorE28D03e9fM3xPHQWa7X25Ecy8HwkhkNigHBpAwo32sNkv4nqp
iTuagv/FkZ3DT6az0Md6BUF2hVRP4qDEmQACNfX3ZpVZBb3APSi31kqgdk9IJ8Fl
EwPiITw000nXr6FvhIKiOBe2KHh2sJFh784dxGqhn/DL85dufOhKsVwqrbcSWV+h
dBXV4G2RNfio/Ou5DHANqBJs7tAClXd3pl7lCoedoDam2DLpmdqDLRWPpQB/F//4
pMazPKXJdCLYPu6SpP9CLOwn6MShWVaq1QLDGlGSFVHg6hUGUB4aum1U2+69C3xz
FXy0m7lRtxnFHfd57LCwLcOS+3NCiJSxICP5fkW712H4FGMqmJAO5YqotYpVo4/z
1GnLIkKOpPKATZgU0uFPmIBdCxvElw+osP2U5z+eCDJzenySsSV2iTGkbEtOCHHd
TNTyoLlPzM+H05oyC+IbLv5AJO+D8SJ95xRnVm3+mbs8rTZD4bLkN1btVv6lMkkF
G9ndphijjucySk30FAIJfDZCaY9IePFhz7Qe7Basdj27mMfq/gxqgNKQRBBQp+oo
+uXAKCNL8A74JhsECRTlQOrB64N8pplqmyAC07me9q1W36KMv+azyr2UBNTsYhIm
vHN7INtWzbKP1901uR8TmqD9CNlC2PIgK08PW8yl35lQmf/sOyqEsN4Xv6YQNjjW
mR2EI9wGRBOpk1L37UmDv+EfkZaabbQjdIq8C/mF/XR/vbuApK9YslIZx9HQwtus
XpABcWLVn5xF3oLOAPHwMKE9LWzZdEBb4HNtYME16qkMTOpm5+y0GB5iYv+lokJ7
JzZi8LLkrrpgW1GCk2sAGdC3RqYQMRdXROnN/K5RUFFH9HYi/rMQI6LIIIbXzsmt
5V9Brg8jk7/EY6qaSJCibfDDO0PPCoLDLun6OKkketBrLk0ksvXwq5+xCBhu3feW
9IyHN11XPbdI9l2RmSOMbplA0gNWpNo0LdcoQCCvVWNLInhCh2SJOOi1T9iQndpj
3Y1ARSZIXCK8StL0GQQvneH2sQWodedxUdvW34QERUAuEN4S7nPOQIekuj7TAHg7
BUBIN080qA2lCIt2WL0+05e3Bz/csjb2eI7X8PTiHvW4IYboOEcphFwS9bfcqyfQ
79dLfCCj5++MYStJCoL7xYiHECeAqJU1wWB1dPK/kpX2PI+I2trO5pN4PJ5E5qPc
ab8TPRV2Nk7LFRlg6OF/Z5H+4quCSCj5RFRYhsArj611ec4W/Ve2J105j6Z+FHwZ
N1edwz2KMOLq4wC1fVsY+o3dLl1og+3tQyW7uHGZ/kXmvBVa/zhkODLM2lY8ihEJ
ExJLQqYenFsK22xIpxtOfkereNyREVkEz+jnNa7M++6BYrriSlwdrAMb9wem4+KR
Y8+QMTB04/t1/Gjy+3snVi6rMeFgfpCvKwQtyrhHWUZB58yeoARv0xI8nSYdC8rX
Dp1xErK/6EZ33asGUBjtLqBEwsM0+bP7uSaU8wJaYHs9YatPvTgYfRmkDNJxbRhV
w3nwHyZMwEbWkmPfsU9BiADaXjJPWbdQz2827EE+dNDFqZHYpgohosog681c+f40
qKN9y66Mu6X//7dCmvzoqyhY9jI4lgU7DGav0iAPkVhrYB6M/v+l2oQcDJK5wxhb
90jgV+4XUMuTq0WsEB39JcUjUYJdbv7koa9+gRkGmvrQzV25u7fSzF/zYXuwljQz
D3auFsm/g71qA6K+lGXOmO4hnCa6F5MAUMOvjdx/FFtet6yxCPImc5qeriSbKjij
3E6naEs/Cp2lQ5ks1mr8Ll9jTTj6pZjSHzf5FbJGHwK005AwSvoydX4yPkmLpeeR
09AK4lxr/nvnCX5TnF8wdxKiTzGpr2tbpDlH3tXkg/ii5Qo4DNnCBgDbyg7kqNoE
2WUOh41GhN6fuDtNccImmUGANpPWLGNZmMVGbAuIKAOxmYHt5tiSGJoD18D4pGhf
tmL4DW+XfjY76CucxmcM9zgDigkaaUgtn3SwsSzfInz1Qk+JNkC1EpvI6An4UFlV
vbqi6QjDqy2Q6ykpYOC0h4zqj87/lDDUV2TSx0IvdsLZIBgcTH+SPqL/Ay55XL51
ueSY8TgpzjxdsvU3J0w3doW0DJW5pIySBjiwdAgPwQC1jr2CxvlwwucYudeu4nyw
ea1TYf7smGPyVGjLtZhaQA8Uk5d6glFv9kzcglOR1bKEos26Jk7ySk/odgixPWGh
5DLaBsNkd6bpKH3r/RG2em6tKpDCI6NbjrryoOhPD2Qr4+wEi6bV14ioEKAUWGu5
2nAULzGr5faCapKANQXGOE3h5A+DZ+CM4KPbqxtwAyXQSymJwgykkXfTnkIz2Shu
2AMtQJPxuYntr35lKK8NqCNaL1hAItZAIOqozJOg5i8OjZYZYOieQLBNuXyzFQQd
CT1H0krRJITKJYsJGBZ1na1TOKMcXTFgVmeR+N1IYwA+0MwkZ0b8uAqPqQBoyjAI
nRFEI9jPyIp1L966qkaeczONdmmmPCYds8muRg8wgAVGDYIDHy1+5b4RvRBkoJ00
nvdOPLtZ6GZGo6agkeDIq7m/hdO8SwWUjclMzyp4n4v/KXawDEDSu1OkpchGZGLh
01rP9Hq0F6c8Bfhjlm3f4b9O4/y83WXBIiE+UiR5AolaH0sYtAKGuxsZWGSnKOzc
0BoJ9KMKNozpdcqXesFphgA3sL5u6aAbNPr2Ad/kmTMJLM7nRwfDK1bBOmulEff5
WjW30feA9VFFVNuS3oD9blyXrWQ5VfFGjP4+He9SatYn/NLxg73IOHEdpAzlozcl
h1xW4+DWnWTAABOz8AdThDJJXFc94/dzpzezDK3tfc9FO3pfhHAODwrrxIWBrEUy
rOhPRCQ3gdsp/eRBpLnrARwIvk9pP5VfxQmxeIJks0aUzUqzD+Sk2J3IerSoDw9P
OEbpEy+rWjohvcS4l1UO/5Cpf8UkPdEM3e0GI5UTjzFkpeFTpzs3xY/ZeiNUEbTu
ci79XZdPu/kYt1HlN6jN4T3/OkVR5y+9of9K5NjSkgslvkKmMHmJG6NWgFYOofmm
bvw3Jys5YlszPt+OQsOf93MOddNGUJXtorfGM+cKYJ0/luflxO8z+GYEVMFAK9Q2
K4vVCPdFL3SiZVVynXuAj+/D2dt1aA6Egx7hnLhUvjbOSzs8t4BY0DvDIWCiB1CJ
6/k0k0cH4FUirsJA7g9EIuBpU9rJ38pbcFWpTyuRDanGph1kPbdw8RngV5q1+BFz
OqzE9EZPvtE0eByCiwpZkPtdyXU2Jz6rNBU8GXJ7w1JdegRl4YmPyzReX4JkMQKF
+UGzZy9vA+xtR58kOSFkItMmUmjBAon+Vu+0bFtZ3OOtROCtqfwjpy0eSvW0zUfv
VeaifbibR6SZAIgP/g7SLWdNiuEiAkKKSphMfmr/dg7mqu0TvFMLeaF8r0huoXKQ
8jJUGIkRrRp/3o7YmpzOHn52l5ty05gEoqqtrDWiiu6X/sUOPxIzJUpwx0KNqdwb
Ii9fCTyRjr4t7B5+2D4vXgJufwnJmv3w/hZypjA5GXAOxNItnp3lROd/ofCQFlbs
BL4T7VQjdJ/i8GzQTqTuLccUfRI2RSjdQ5P/aG5F88Y3a7LbyAADLa8y5SXSZZjT
/XsdiDknaVDGNr6SnUNr++kv06uIOIWl4E2riASGp2bF8WEvs0a1kHTtXK3BFt3z
aVNUqOKF3rznoMDTF6pkQ8aLnfe202kPX0Y0MZUPCExD87OXaHDWOLvk5zc/8+YN
ia6o+gJtVEvCaS92/dnX6JVujy+YpxzuFlzKnroxK4Pgg+lnH/J+SbDqMm+1bf8s
pNqiodsBQQR4me/c43jzXmxpgb9PMQehwv75o262LEzPY5gAg8N0/la/ZxBD75Wd
SxUwJOfQ8kOMy62BMKcOxgX/uVB4HtWZUmsunPFAx6lL/ouqJc5If5ThGGFWigDs
J80U2FjZR7lFDCorsFT7ToW6GVllnvxr9dbPW8ib9lEYeiBIUmLWpiuquWqKsqdc
SPhAxr7TQcQ2Ca+aszN6axzMyAabL9IdTPIMSSszEkUKCE2WXh4UyJr5Bw2aM1T2
TyOa+LjUx+JtsYZ+Ej6COxOwNTueMVb4Baq4Ok2GwF+B3zqVRgqi94DmENNw1fmB
ZluSvu9DoGyVKou0MpApOBNKqM8/6aB1NfX5zKiPjDanUHk761BJlckd4KzKmiO+
IVinrqMwV3dhksCPDHclNueUYUOdTkQLx06NGZ5bMpsh8udFPY2DrE2dkVTAfhLm
bQgGRosTMVy6dxNj77MMVluGLBjLz4tW8awkuK5bjbP1H3MCTQ42430KWb/OIbQV
Mzgt0UUfiHrQSDaNMUau6kwjnWoDHszbaUtkOB4++WkK7KjlaVcOntvZx4r92jxW
PYaGBehQ9weKjLHzir/mN5+MItcS6mRMEtvQ1pjhzs7vP1lqIH5UIsmIBsZ2Xh8O
FZA4H8i3bf0h58FR9GYYy/qWlR9Skz7n/BuDB+5UlWncwRADqwRhl/BJyxK+09Hh
8oYSBXLxEnWXBQdWC9m1olA7xm/4Trv3Lr7B+xkBfLHTg+eoZ1R2eOyuWSej5SdO
RQngnXdNBczES3a8zJ0PaFF/kbPzl6QhZ71ZKPBufrswb1Tr4FgKPcwnocevt1g/
wA1i6EDIjaPI5IKt60xazGTl25rKzFyMQBM1SlKxtYLA0LlteAJuJkriId4giRSQ
33ylNQqkNrW5rBkni0kR1jbFPXWWZTsp9Z3kGKpE+ft4egmnwTP/elTLCiPcDfXH
uDLlFWeS3/suFH1wTUopP4QSMKi//kauVb9nlsU7yCzYVK3WhEu8tuzOfgvLSblr
4Xb7pC9+cwBJwU6bGX/SbYEHuXnVDdISD6vcQhmLU/SPd8HCJAmg0eaisCDpBCo7
VrkwYhoK2oRfMpirTs7oJwmw/Qq6CSdCFMWY81hS0FuT+J16sGd6syG9Gp83Uc6w
6l2nSUnsCDDZTYFD9myZC5U6f5C0q5v5LDG4/y0+buQCRnHQetWdzK/EX+1XVmIP
ivzvirrLjLilGrbHqDVxIkcu5KAzPtp9UMbiDOq4cfhMWbc1LqhZU/kcw0kJUz7n
F//koFJwnt7j53hB/F6OUQg20noCxmZ9O/2M/Q3UyYyuLsiSrhujlEEWVYODijGN
GBdq0nEz53lwlgyiF1yV+d5dLvF5GTNxZ43exWayyOipXyqp5GT5TvZWWSGGS7/k
lNtoaFGjiZt65Fyq9SHm/1F2xMk1U4JNBW6yOpZPnXs0W6ffVMCxXyhPHabiWJw4
2UQiZdu6R130gHIH7fJhCuu2rb4nS75XAz0gVqCuu9fIwStvc9VQ/NZGi2S3ry/L
NBmnbRVmGDJL89YWnQo4WjGnvLC2kX6cTTpBtOXEnX3ukcwJ9+6eLaO5+ccrL/fc
nvsT4ft/yyeEJzxmPnUwrIM5YobyK7jjl0Vp59XO69byzU1qAW4BGUVDWgUcEPcs
ySnGf2zpLDhH3ks7yxuOfSutDFaSsRRq8U1Kb3bjhn7xmXKHbgIft6ikYCFupV3X
sRr2dnTzfQmPlwlt0DdTEqDVY0SfMiXuiSwfIyk9HMlzTJOoFHHilwLjlOorcPcn
vzpTUk0hAjDkYY/C2JD/YMHvWjEe190kXqP9S3izgEVxS/FERO+ni4tcVpV4lOlm
H/w3vmNUL4jZ38rvsbqfFEjlRLOFxIRnxvU0yEfoIFr/c3hTMW5sMmykNn2jXaHh
RUYeGLBJLrpN7QtvEirsws48BZ7n0trrsm6+iRicpeWoIFL/5zeKpR4mJrlmBwfl
YmpMWAdSpJ1pmid7zl8RpeFJrL3I8CwuqkCt75X0BA1GwDZPYHZNLMaCAeh9s+pW
P9JuCJbnCYBkSvVgYEy98zqCmf9LqVLH/iQ/UGG0iOQJZ7oE0jG9ygBTQn6DWtcM
JQc9KXA/oCcUO0xeAPvELemsQUrCLAd7qfsVqE58V+BabKs6Bso7LRpj0NbzfPU8
5LDUMykSrAh2Uf7ojXIuYxV2+l6EfNKfWt4TdxqjITOuYKwKU3UF8lYIBReA7AW7
ELl7C+QlYg5qDOPDxMO9p4kbjcyC6qSXA42EXG/8MkC4YKVSLtMdPSOGY3zNg/WH
dEO6Fksitt1adHBldrJRYcxc2OFbbSb8H5C5VkfZxip9J/W7anK89p9XVfUE7A7n
reyyUK+HnszlyV9zLaCRg5pam0feARLjD1O7E6dS1WYfHPT9J5Q2xoe4gOae+o08
5OsqmL2XWNGVFI1u3uZxhSGaeahL5sU/B9bkQw/xvJcJAmDHg9hi5VObR9uTQZtA
zYFKSObEy0BJX2Vky8FOGB8Z8tqGJeRHHtFs1baTuJ7+pke1gPJVxjD+ShlAxnUl
pmJ8Bq+O8u9s1ttiXsgdPMHER2SHidPV82iJ+J30w06a2mWgmCbGmQKDdgtMFT3c
MOJHdjwYRPHB++CG+u768ESWIDEWQXc2PXZy9jKqUv7bC2f18Ulh6DMrWxxLnTfn
aYkystiuB3DT22YWnaKS7oa6HZ93APTgue6ivTo7K3A0KNE7q/RCXK6HFt2wWnGc
chhu1QYBqZ7wmQeG9DP9za/2ctXQ5Z/ESjYIkgIYb6hzXDUCW9K2AWTZcCq+KGey
eefdZjc/NzXxZIVGEgG2QDl8VPSvoaNU2PxHmEYwx9XU8u3qhAcuKiuQaRzkj+3L
Cvzip9zL9Azay/v00ldNd41Y41SkU5mP0uRR5GsxG+lVcEy6a0kaaT2DTeEnV7wj
7mSQj3LtUFnaRMX+T55NsFVRlEVfLEHdPCVBo/3xwFh4MQlTB3DE5/Do1/qZsbP7
HGB6tOtsckqaVRyYTVhNpUrm4Dbyuanwi98Y+OEEbK9ylhQAwDv4/LVMZunypNb0
6Aipvx77Ak51JCkb8hrvhCZ8PQ7WZrJYowtR9u9/9jhgqyFoP75zxPDZYRRXHvZV
jCWC6siLGs11ox136+XPntgNr+xInt2HX4DxDdHucdsbfBCNPC7WIeQCaKTLiwp4
8vjDbGREKd+AT9raR4/lWV5rzZHhwSy0iHAGHnBdey3JWxoHo+ULXYhOO1mmaGZ3
sdMeM4XSOIYltFjzKp6MeCUqqAo35tEP0s25W3Eb4CrGuYFmTG1Tw+2uWA8Vnzsv
5uUPDeC2xYYTP9iCNNjqJ9KOQZw1sXlrQXDS4ApZoRAP/Rh3gUT6hB/lROYUYkwv
NM0rCBoq8qb08yuXcgjCFh0e5jpXaZPxvWDiRpsV/axW1CXr6Y8ywLILg3mfFR4J
gFsOvDKswENIEUi/r2wklqyOBh/vJJfwx6B0rcoowHK/X3DjSmE+egiKx6/lLkFQ
77WRWX8pQGf6omzrUfS3JT83FaZjRuONne5BNSfsF6J4oiqMTlRT9lpob3/9a+YP
6jyou2OTNxA5Zjp5fyTUs55QLnD4c/8MZl12Y0RO20XlZKyzjQW/YRpOJh8lNrNW
7q+KGAxcvN4DWr1TVI9KouOa4U1z4BX9LBMgTLkVuI2K/nWmoIumoxBgTJtrosAz
mYmGycdIKeCs74JbhXEj0HG7NDki+/wjZYImCjDE1rhfLbOTHBEqczBK89pmYLtA
Y+2t1Fw9qYhehExc0rzLx2Cl/VwDfMm1MPs/gWzZTUEelo+WvpiI+r6SrNB4CvzK
3stg9uXQUpHxu/OjN37axS8CRDqfhBBH0iwiHuArin0A0KUNz2nfrF0EZUn3dHE2
tvcG3X4hVKcUtRc7AZ4x+uZ3upzbIlxY1dN9sWLsJAMFcSlHKFjHVpdh5HcPamaf
UQF+ewdgBfyWEFdFvLxOwkr5Vt7Fu5xjIAYFZr8ao6fJB6XTe2ehIw4PPka1PVe5
3N35TR9eSL1iS9E84iwmjhCAihvVqWlJwSleXrMNFlMopojnpS5wjZMq3h4Q8qCw
dyRbgfCGRF6250mM+2a4ThaHifFIj3WI7JLQLIrQdjDmxVtESfiL/n3at6ky8g4/
rYTRQOzut6v5YzFHLWNfcGKJ6MpMtSeTxl4RSaJA6xceDMsivDJvUW4sWJBIGa0K
fz6lWs1inq08BHt/7+7001KTt6zVaLQzMww27srSMsEK9qP3ctt+fPRSGE4vxo5M
Ht7oq5OYOBu++ggdyjvVkYj4uQ3uTu/x8pPSOs46Rk/YVUUEIOAcIjcOBDu+voJ8
rBhFG3xSuupc8YEhUxEAjE6HT9RoFVSyJSCLDR6nHlSuoCFZcXpBUmQSO4sMEbiW
bWO4SEsl+Vs8MTWCyBuO0qqa3ShVEQsoIc/0aTQnROp1vAJDWAUgH40eeu05gGH7
64pAka76ISK3vxerp9/V4ySmmyqJjyqHHkppCsCjjeFl3f8rNfS/XSXpjMWhv8vE
ezGK3u/EpKzQygXhWU+gchbS4vGlHeBNiN+U8qY5p8nH3QGDgH5dTurEFHydgb1k
DCOH/Pyrsgy+xDEX/aiGtTmc81mt3dBo5P765skGalwuuxIIcxOOg2r2uge+7axr
RMpXD2JeXjN9IfUI5xXFiR17BuxrGa21feqbasSek/pcfSDR40nrEVECg08XHGdq
5mxBY1MG1rm3QREndDU0beTmev7AoDQrT3N5aXcQFVn7cCv8MzXfyBUSfrgdvBNi
AMYRF6nDJZybhkv3RIGudmWJhDhXA5A8ogj7jX9putGvDEcGjCZ9xIDhPiXpCMZF
/JIrJ3tWeQr+izkWbaj+RVvPKiFjCQL6ulcnFT0iTzdYA8nULbaZmptIfCYFWXNG
WW7i7H58Mh+w5yQhys+uLedukk+8L05sn4bGSnVuVFcEVVX2UHmPKdkd0OkA4f26
WXkCGE2aSafDqfH7MwqYOEXDfPhofee9mRmMOCTLX/P6P3khbU/Soy3Bc2jVA7d/
RUXjJymy43grt/7TQ95SfEp9OVSAn5LcJwZv0D+ZfkAYrhLB5NJ9GFs+iejXXk2C
hR74hxZVfM5hDlKOXCoxQD8IcvbXAcmVkcVtQ69wMzTOeJQpuDruPEtgk6nR4r8p
KPa/WftNSpFcZlY+gSd6NeCf7Ys4VQWw4H+GvAR+dalrejIqkLSTF1XgNGnnhzzN
a33ge6qEhDczSdI/D1DMFuMoUq/whpwLMgvK9iznrz1EFFe2IRFR7K4ocZKoQmdy
B7kLnpxUiDULRjRiDZokzqh05JaPfpEV3XZBI5GnZVMbWUc72vKAL6+Rbeo65IiR
y1IXl1k418XxjVKKM23G2tIx6Bigwn99iLWJ4/MC07iJxaoDONPbkmJ1aIhYmHAZ
3T/FY/feOhT+KNBnshG7n4JTbAUkppzoi+FnNIaNgPyRHTCMd023vfD7j2hVNSMV
dJL040NOIbzBYWcDbUsyyWTaQIj+f2KjJDrYNvDlcwil1TBx2UvLzB3lHyy5oGab
Reee0Mtqu7Vn/K1Zd6fMkeGOaHtWju1JuLPmp2h6juanA24MCEE4kZFDYgQ36lOq
gL9QP53GnP6tPHp7Fsni7u5nDOd6j0Fuq5rCMQIT9gSXY+gHURKcLmzi7OOlJY1E
KjCns9o1fkvO0fYIV+5D+mxjDLyd4UbiyXKrSNMiXRx3mF5dxiwLWsin+H1I464I
McpKf5gSjVeNqsPtbmNd0gG3+H3SU0YimoHc5BXug2v2nRnjiwniOgmlRlQaKFrg
EB8rWJxrS8i38EOpAXzcbomVS/pbRkzZiTrv1Ogxnic3M+lJu1n9odyctiJqh2yT
6Heg+ZcZ/R20NJ3WjNG8nteRGqqWejnlP+cBnEtGdtDd/0Meh/EununzDx79HcJ7
OytWp3XBXWUC2GIx9R+98JjUJ1i1l+vmhRS4NUxnQB9PfqwRz9wCX9mFehATtmNA
aK5wlqIFwd2I1L6Z0Z9Jtkj4VuqSidnxJEZhs+X+wGqaKBI76wBGhSHK1rPiGMl9
Hj2pDA1KpxMzt0E9voH8WAjDBynLeKK96SvigFd//gGSSwGGfBEY8xUS8fZxojO2
OpD1+jVATKInvpTr3CGlIRt52dcJEVopOkoQdTTj2QiGZDx/KuFpyOwjz7x0kppU
Mp1Tg4T7bx8iWRR9rIqz693b3JPLhQCpXPSbeiBjxHl615rt2UqiIHsKFPv7Po+L
mSJz9mnmmNvOhSkatxPyzPFjif1rFy6cXp6fopjqgT3X1S8nMEkrNGzPnN2AKUPn
DQZmICGCi0lQb/nKQpWqQLRQRYwLxWtIUXVzPs8q+4RVVyRexqOAH2YqSxzRjKoI
CpaVwKV4sbK3rCI2rnCTaNrESqWLH3SJy63Mzh4o1BSyCc7w98NtW4MsuEtNRq5J
2slk1CW8ZRoc/Z34G5AfdfT41CrkeE3m45e4qFg/vce/bCl5kYJFmyMiIhpwtWkG
Xapl5jb46D6UWZj4ul6Ay58fQpHdIedbjatOC6se4vLg16vdmH1AaZjvQzKRi+0m
frDr+grsl8Vz6X74AyfeKaFfzt1tHGTj06mRC09QmhGaRJPcmFXuEfPB5o1sUvBh
oOutpG7Xhd4imeC1xZy2v5hpN5Lg9lddRqZBnJyz7AY9UOz/jZf9I7Z4N0Mwc0dj
7gVTm9I07H028I1xOkdSMUQupTMG2H8geYmpb7E27XUcxZUDN4BKl+yotBmzZ8D4
pQT27LLzN8Xss+NpVX1ulF2tJnoqgb9s57ltVM61YfilkolBV7tEpzC6ECnooV24
J6hqq9uF6hFTwapedu5A5mFvYPQUssE9pkLATK58TvoQ6EWq9IcBPyaUt2k+06xl
0NZ2ReKFkWDH0eap4y1DfumS2cLkDNnU4p3PerST037QN5j2dhFBmydf9w35puE9
+TwiLHh5RCFL9Gw5IR5AWdtlZrmvdyCrEI3FvxoL+HT6DK6GF/KxVeWCH0naBrUi
B3Rjc/JO68xShsrHFY4gqZ+GyA4ir+nFTtx5yuQW2bCFC3SZdmCFlBbjGbihDJ/3
cVCbRvy8lXWVnyqfyM3MjmyrZPtxrI2veSBuLN34dh43EcYgsXRzKeOYDCYltPNP
eQCp+/V/fOu3JBiIaZ8EdiHdD8uiV32p6YojcvGopGSLgRgs+BYtD8Cu0iBH7v67
jCHGK7ERNac6884zPT3ow9RIYrbm9oXOaIx3RTcEegSySs/vx02w4UexV2OGR9Zr
Dv6gxaOZiXXXwlNGEQ0JFP7Gjbfg9uXYJfvj6++UJRHnN3kSU9NpiD3OnxP/FLwT
EPxlpYzlsYhlP+ZKUI+Lt5GDm+mJg+hwLRIPIi7dbO4u5GXhq0Q8TE3HwBGfxzLz
CYhWZjIBBDqhU4CVlU7GPH8fBwo+cKHdRZrZpIft6B9FuzhSzKKv2BjJFkiNSiLJ
jlu6b7uNYvTLyQ9p1jn3UxHQCGT0b1grQ3N81C5hXID0oSvMJn3AQ3bxDLe27D5V
LaF8Ca/Vd2wEqT3lhAOA/al1dkoR/ZMWEKu7PQLX+zH9u1GSGhe3u1LrLv04NA5/
jRufMpEKUi+czEYw7DlkPnPABNGuuYzl7aSUaFi02Epq9EgnhokEd/MV0q31WMXd
8GP9r6UthD0MViQjaTos2P5A+Mm4ow96GXZcPKWqAcBqUai4JAfuOZrQFKGQFYwj
lCK2DKvIx1wygD94GryzRbWyOrJbc5xozc9nrqgI4FnaBMjpP9jeDx8Mdix7ev17
vXl28dq1KuWgWjiMoL/VOGJvc3oF087aq7L7VPBHTrajQcJljMPxqONm9RTZ/zXw
0OqZXuoPuVRIBJLvt4pkWb16SZi6/yocyTRr7ir7j9XBF8nRFzbuuNVlKHLTQrZ4
MGi9B+ET3VlTXOLyDhcJgsh30GBg6I8QXkUIUP3ptbvSHYsCVMdu06nuShOIB8Z+
X4YncdK6QURV/pRtl55d6gH8G17F3LazZjGcxZ4BYf4ZKNbnFfgIDBeBz3o1XLCg
JojDIJkV6ucY1Mt1UZsDvVf9pDrMZhxJAcMFR4jjT9p5Mz3rOy70dZ8hvvXe7Iy7
9PeuL41n/6xDWjC0eiz/dYIfhLYViOQl+w+8ENY4PSrVqiZYeTWUDPAibXKr2CW4
Yiyi5iFr7wDP4IcABrAWoQE7J1wDG4eSoIeRb6VS920eTCiL3jPX+u3IugYQuRtH
1yh2n9NRekKq1qLLBtpMox1NdZa6hLADNI/zdtwDyGb6vJHKfdvxtvJJVUDERKiF
faGAtl7BADOKHi5bRV889FvYufjSNyWHFL5K5sCf0fnDOjL+A8hdr9ucvsdxq9tw
8xqet71FnC54lT/dVKy8R9zFE7iPQjYiaxJhPwLXgB4JtOC6L/hyW4ePub0e1glp
aPrUYjs1QhIBh/HzoN/wM7zNN8dU+rC3HbmfSVxA7KVswJOCwcZUV8gnKc1NH6K3
x+IeBbIYHBPIBehJwXJh7Y1RbylqcdWxocn1JvFTrCzHtZV56Lz0zVOZ5QcJBxhI
8U+dSQEP67rtgKUqIuXqyf5HO8TmDR32Em/ydeoyxedRMr/6m6iNppUKKw9/qOU8
SPa8SVgRp53Ylfhxsk0WiBpldPIbGFz9C4uLSMvbJ9oEApMT18BTiSwJA8bxtw4+
Glo8Nny9LpYcdaZ6HRYW8c29zenChr5nWSKkAlbX62LQdP5QjNrFUNnf7pRnWOOj
qQagXvC5J2yCRW+4ywgPAq6Emv4a8xPb+mnqzrENin/jiuQ3Q7fNdGqsLk2WY2Pu
ZD48RR1eqW6J04afUqheZNb3Rz1b33Q27vaRAfAUfKl1SqH5E9w5cUKa2/ZXSb25
HyHUzMp0aLWCyFoRKKvSSs7iVdd+slcmr6Fz6ZGHQiDdL5KhJQwhMk1imoYtkmzo
FPUhwifRcUMRdAKHqNc4HndztP+LcS0iyCeMD/LvCAVZMjYFMQiB69VY+8rBv64b
h3Xg99zOE19iVx5sig0fv940eaqgmw2VZW863/PN1fEX8u+pah5ke+ANRn64TyrG
FX1FjmR8MbdqV17xdwLks3KZn12b/pkgx79qgtI02fdQLfVg6Z5oDSpTFc7Bi5n/
NJGpt2z6mhKGNKjtk0xO/e6LYcAX/cRM5yMqvLrlVymIz1QHhnnpRumNznwjW/nI
Ik81y/S4Hmhud3mEqu7tXOM84P9CaO9bTt8RjhVmP75JrrtTwhhEBVCqj8uRpeDr
I4YwAHglSaH1npjghkwaaQip0s1e9TO7G35S3LqIhubvq1H6yDwWEPUoTB+NXUg7
v/xYXGEjA/NatBj0gTcueRuYfqajuZSbOWs20pKOPuJ45kULNYb0/5OlRr2ADEWz
k3WbHUvdLi7tLeDWXrDTkyxWuIlPmOvPaiS8inEMOUzfODxzJbK5PHzXr2TeoOpi
O7AgrL9p3ZPKmuR1JYPWBGQZ30Usr9f/Zw+K2p8bG19NY5elOljYOaT6QCpfc3lL
SIC1CduX9/ERpm0ooVNc4jj98su21I7Xy0Gy4ow2kZ7p5wuslo8UyZkqbic1cqIA
xrN8qM1W7P+qLy70KRcquF0rKNogySrH/8p7+1ttwWC2PUJLs/5vFvNMAcgc0vz9
qnvdZi1m9S4Etr9L3uBZpMtNPGN7ZddVYgS7Z0faAmP4vPi7e7rjISQLQsejfp4s
Yu+DMk5XdGvrtky7g0wKPbXz1CNyXb4+cKS077cR2vUpU3NjI4eJttt4TlnN7qZr
3tBrvTvCoo/UZTPIE8pXUW1/Rq6p7vU5aIAoYaoO+y/d5aEBUuIt9W3aXgv+uV6Y
CzkvLm/dGR9Coj4tk9Q+hLK8SeOpgSSe5U+1AFiQjthJ84PgcvwMOZkbKARKqvcC
XrdrSDPfF8MUsNnLv6ZPUq2BqfrOrQG5HNokUCYqcmxn7VS7bRAPy9PiH18HZ20f
k9ZtFCAnnTd6upC97KCSZpNJ4izvRQ8zAigjYzdKfWxNRUqzZqCPrSasbbE8t/fy
0pvj5WnmCkwHbf5YJGcyKs+VzlzGIrvnHmsUzWHDdSJhPrfIr5eUHmSVDLPXb7+8
oV9XoHeR6FFbhBdnvxwfAIML+fGVOWsWaEothPdtGWZwWKQLmyn6Q+ON56Om16JE
+Cq0LqXKe9jRFTBuE7RHm0W3SPxgBv6pNP1lGHX/1+G5gYEdYXVGQ+wnXHH3wccv
LJo+lG7a02xMjLUBP1h9ATc/OJ8SPdI6eiQfVYHl+VNmO0Go+qziNC4Ao19QSz/g
sKB9T9k+3FFugeekpLKN8aQrViCvTKGNfGGuQTecclK0+YqSVW/JIO9vBgyI2Gjx
DaZDdcSwZ9PTWD2gTGaz9uFwWMVbqm7L8BdGVSKZBhNdTNmlwKJYSyT/7ePgOMg7
5965foU+tx7g1tNLv3rirVggrEFkyD67ZUsLw9NDwQQxYXc3+6D09eLU0yEuK4km
G2yw9gmRr9TaFakH++vZ6zQDiGBXdVJ6+dSfcDcq7jDkx3nVT7Yr6Hf16mX7g7nh
jJzqo7KsRRXStWim/nHN5iFZ44Xt31mzHQ7PGevXfOkpg0mANqEs0Vo1qB0dr4+n
+k1RrDaGJiohz1iMnFN8FLNOJogbgP/NxUFqqdb3MVcj/IxBkrKyBNUh35+GUnUr
RYq4eb2SwkCVPLSAvePJz7lE1o4WD21RsUA6MJW/xbzgWqfg6DOkBJDT2HULJoJr
s6n3ZA0WuKy9b3/QOKSqqNjx80OpDa3tRMV0sojKdj2X5TwrgLHDeih1PbaXZreO
o7m7D8kFZeSGTOVNinMgvj3a+BlXVYN+zoKZfeD3jXJ0UXNCSa6PSHAdKuF3wEzQ
jnlYLEE8/IvgE6p21ZIOtAsj9sqHRiiNmISBmuHpHuBh/QAn5SsZM2jdqU91/Y36
hWveEXUfauInb7IevPo9IY+tGfHcRi7ZN+akq3Pf0OappGu2wX82DYp5bKbibPl8
fs8klerFGbx2EprnoaLsxI3ojvKK4stI9+JWJJlND+llPE0V9nlgcgB5ClaKh8g4
CSYkl4cjWMWdLnbHknqdNr/AKZLaMHFIictW5nSgKi0BCWD8rUMjtsLCXI2a0jbS
tEztbcLEuIF9F70/OPm59twH3BEhTSi1feD88cndC/5p9xUCTRBQAfpS1i01IxgB
AoxfeRwYcb4Kl1aecyvfCkfcdgSK1NDSRdAIgwpY45O2fdzm8O80oQxXxY0kdXZZ
1lzO5gJ8oihapY773cR69vQ2LZQ2v6dVTAhVKTcd03HCzfgxQdRcozzYmre8ohc8
edjC2D9RGBN5DDjC8EEHvf+vBiLfFhwfwA5aBqm4SukkI1dfo/r0FC/y+X47ubIM
TP4fB3WigRsgHjUxhe2SZirJQk1dhCjChtshlunZ5BHvKI0R1iErBAmKjwmphbdD
PT8MP5Zm0S4I3W2lHgPbhGUghxLiGkuNkruUQFL4Kz7tQ0UjEV1dZCAn9QcawYtZ
8ROD5ZShz+EJVAP26KgVKPDlNv23mNUH/F97CN/TJMfvfivTt4stOU93tc25C6Xt
Zo3sJX/iVY1ZlMMegDmpFf6Idt62QuQrXDXC9/XtS/dZu3R2NWBvrdNcSbTZEoSW
ZAzUKBmaSrP54XF0iuEh+sIFiUPeSgoPvodzHZgUDu0sbuQoc8+L1Qz8gNXEjfg4
6i60e/I5cd7Nz+LZ7wRttLFHs04tBsIbyhk0+aI3mFJfKrbplPt/+Dg30GzJXUib
3GADiBqibS1rAhzaP1riBMaT0rLxmFNaYAdftoS4ZXzARiZZLr+HfB7SUuxveM4u
lUswSdMcryovbCTkUUFHQSQhWGXWlRvC8TD238b/ZBFkc3oprCljbM3Upp3b1RE+
5MCa36W9CBkVbA2j9fdgcB/r1hmmA7rDvtCA9UqBUts9kg7G2GnQKIkOcNPjwmR5
WlY6ygF/D6a6IwfBbl6SYyGxYgQHDm4rzFpJfPbtbV9dkMHcUKJK2b1uOEGlYfE+
vAgjK3XyapzJdi3DfiMFtM02Ti16dbm81mzsIFOZPyVY27G/Zcz5VP6e7uc38jVl
ODp4E3n0kEujKeaEmAayZ32RvyqePclUB22qhzblViH0KOYmugYOm1oqNXRQGRkW
O/mIG7jJsbxlXgPzMZ/qU6eIGx2/TSDUiOAvLkDrilkjzNODOKcrSeC6dn/pOBnz
j00pUD5ARdtdi8UoBzL3bLvzcDyznbcsadxMIbFwT5Y6FdDhtHJuND2CBBH645Xu
E5gKEuagG3riJ5QDhrmhn7v9t61h8PEX4GHkQfg+QTLJxVIdZdaxGS/QpOgFwe7I
ohrtOr4bFI02Q9gJAxqhJD+8YeEHaB0z9ueN+5nfp+Npgn/yMbZ5huOJ4rmB5JK1
QJidHaARXXT9JmkInUZdPdumCUYMucizUjDJvLlY5EcYUZC5ED9NwwjwnlV7BrgT
4NJHPlzK4kD5pMIAqFv9m5W4xCULdNSppXqTPiG/mORQaUdm9lX3HFhkJYRr3jtv
S7sCYCeVHvVkzQnmEH2SczlUjNxuwZAB6OmcXoaUG9LQ75paWPMaZkjrpynEtf+X
m3LU2ewck8bffuGz3wwPPo9PLs71uGbKi+zqZoTZlqSYHGY6dg9qO9AI/9vCU9nt
ebtwY9MBGJD+dGRvVFwuWNUUWmHMRJyhUdQN+TIXX3F7cjlCtSn6aOwUtHYvU/sl
0Gf4nHvtZiuhPIwoHMrdjP2WQUR9iVWO6Ub26Oy5ZmsY6SXD43NYbTATKntRzyV4
eVuw2fYUgj0pralgPZyaHF9aPVktUsFr+4EUi8aiaJ2XakFi2mIak7mQqeoifzDU
P2Z1wueLKVesq3l9tiKet7zzCRSCbcQIeT1DNpBZDH5Fs//zmtAls63FBz3ycapT
idigFq2jEnWIxw8yScaxXtJ/tLG6u+xgTaOz5JQz+CSpFT4KU4KOKHIYdVO5TsgU
N2ZBYv9NdrUu8JTT+zX9k9TJKEe7Q1fbwV297rwaccjTaGbBOraY4jvZPjz0mx9o
t0spbnNnta9PXL0BtNr3Yx1DraoLjKJXe87/3sRSLStBAPvX2COBIw4AGeo5UDtZ
L6sWuEkdBs9XPUf5t9iqgLCqF+FIGR5Q1Et79tLMfYgHP4hHBXD6hsE2myBuvyLK
csvUdFiyj5Wg17DtcvAM2Hud1UX6ie0fUaDqJFK2IJpr8P3830/gl/pg9TEo4AkR
3MLvCiIJJFOXvUiGQqVoO5FRW+SoiuOni0/hMirxvlI7VoudaNfQWd6paIp3b8Pn
ViBtqb/t9S13fDtcFDwbxoshnzSqRHpS2CgvUfp4m7vkMT1Hh/xO80zrkUaK36j+
gvlz8CUM5Zvmq3SrPuWPqvwjsQkhu+mGvq7gEygEzna+1wGvXYEnPGyLnBO5Myvs
0bGmXOsVLzmLwPJeTTqIVbOsLGR+t/4btBigZM1TIEratJlKSgr6qDf/TRUulQMe
Xvn9Grf8JROD5aeqGz3tsJfThdFPRKP8Vrc4OyTw08F01kLIcuFpFvxt6uhvDqkG
X10dr5Fb2HQVHqvH2QtIj4PMZrdD3WMPiMV7/1vpPZuv7lXgY84KP4+8lZUkoF/8
2TjeforXn+4z3JxpdGgBoeowUxpYkh9+LTlvbGW8RDgZpyodFHsxwjLbRhrla7vQ
PPT+AoHr5/VUoa8/UKHeHQS8dVwbR6rG+alhYmIzfs7R28p7ruYLjSGHvhwX8DPj
mwpOwH1i+7rFcKjVg4+uTEuGnq907ooowBUGr4Za+DGKL9sumdDVH3UvcMC8obtr
lIz3jZxVIQeDOL0YdDcZTx4MeUPBEzWx7bZxa+Zg2GEmbI0jfq4S9bJnPwLMM2+B
3XOfB+0bdfxeV64LV40b7XYbQkO3CAylnsRJh6Tj6n6bt+xmhp9zCMwUsnzIrUof
mpVIaWhzwQaO0iO/KpgzRgbzTRfpVKYw5Qj7W/+NHv08dBlyt8LahN0uUDaVd4mc
txnOCx7rzTCH5pR/A4a9QStX0hypsWfH8JBqN6yPXePDcloUAg61iaIz5A8YkgAE
qfxF59U+3EZ0Mo/+PoyECSgEm9r8/xSiYm1ZPRHzvVuWamBjWdda617NkMDoQi5f
hHF6zkm8D3s02R32PTqa4krMnKUPk9lqHaU0r2ljq4Hmt68qriy3eLciG5Aegmlv
UFXlIYXjRHd/qbrnmcVbCgBA1VvgotpGrNadwWzQ6uAk7MJh3wwU9weui/tuqh+t
9kTUc/uoPhLdQZKAirsWCV5yKZ0nQ7IsUD9+2bDbe+SNvp1xzAGTo/OD4XUt4L73
5gj0FVjiMiWq8xp6knjayrDau9AvvwY0eh7jR3xbUrsDq2jxQQ6jIRih5ItoAUZK
9d61daC+Ndlq/bKvKqi09RpQJhIi8nUsz7pCys9XbcPc4xo3uCuvzFvWvyVKSOCr
lUi7EYTlG9iguVuXQyVsR1li8SqNnQ0LZyrozxX7I3RcLqwbaOxpPaprJB6f8Uqt
lHh3dO1Vw7YOlXXhX31bzvb79q8Knf8pXpJxO7J/T6cS36WV8E6+j/hea16JVVkx
0QQiDhQwx5nTaNADCv6jztOsILxpCs55rfYXUgwzMtYdX6loPfmpNT5Nrjff7mXl
2T7AqzPUgQjloHouYus9u0JR4StOcnsGkhZd0SkR2nPdmOayiBWuDo/eFju8M7da
Cntpf3oQYsJFJ7jy0BMx22qxwuDyzmb0LmV7s9Ds74pHmo8Ur3ojIyaSHV4zrxQL
95YEui1cBujDXy+yOQETV22cgyqNCjFrXyOqPC+EWM7C/GoNFayifU+NpVPaUv02
JtkhQ+5881jjvH5p6WTa9I9ANFuiLW1DZwVPyWE1HM5Exy5M4M5Qdr3aLlMgPRJD
fS/4677fWqOSebWlLqEoD+9nCgBDskNUroULDXr0JeLvarXoECC68YTHIHTizP34
3zS6V4iUzP775i/XGn+IFDp0zdzFOun/oSdGvf0IYn2ZHsY4Km5kaY+6NpaHKgmK
OFlmv4N2cRzmoM3ex5S2Mqp7w2iGo0xidYCoez4iQdP8L1kD12MmMjcULydhLza7
ICefl9XVCXxGbKTbjlBMe0FIyyubUjwLCcnEuGCb6AiSMQ/NHpbK5+E+9qUPq0qm
mUUwO80RmmL+79NVdDavf/W+mkmvQr5ZTjxpijopri4TqmB2IZv3hKtQRb4RRsRs
ZHCg0yt+ZrTDkxiLI2dgYB0O6hiz+zvje6mNsSP4mlpW84/+HIcMPl/GjoSoiEgQ
AY9HEbSfoYlBdtWKrdiXGlJlclZT3InIiP3aP5jRz4KRHXA2DdKLRK+FBFr2RnVS
lMbvgwrfVhMrHRxxg8fsouixmlgXa9zPnn5Av/n+Ic76VDGudBhIBm2dxKIVI4p9
lDib1Y64nTcC0H1KoQsZZlGU/Zoe2+EzU7HcK4LK7Ui4Ik78M42QCdHu8lpgsKr2
bc79FDprVILKduZvbbxl0y4mP0gWx3Wa8b98PeJ+7tVBjB0bxl3UQ5G4IirBLSTG
0LIuagiRAz1XAv8+eRw2yhJE8r+FjLcXXOSH1DbPkXHN5jMq2QPkmb2AnCXSDqNs
wQxx6wpSnRTKjfYkgu3Bb7w78hpxsKKhcTR08cUgt4voR+emI54UxAeESAc7Zk9o
07/8GrR6G+at+JqmhBPEK/M1oXwkqigPcN7nTg8G+tr0sT8wOzzGRGGbYvczqHCp
ehGMGjVed2nukhJME9yy5tzripFN8JkLjM/D3LPBCEpJpE35+Pz6WdgmvLx5ZqNo
FXs+LEGOiOV4cfnQ2Stlvz0nCZgC4XMJl1VV7rXGWSSoBIDRwnAS60K2N4gJyk+6
CclSOzBJ2lSohXFwuOvsgRJAp59jApgdNJfZlZHNHJs48zcMhl4Px3s/rU2yuIl4
9bkRKhrdrN7R3vd9U2d+8Y4K2vcfmWNRfq6sxr31ZsZUzT02DeefS8WF7aCEI9gF
5Pr5IJ854qITXPo7w78bJsssH03Ld4zwyPhODgKuR3Zy5aEwII3v9WfSip2SZ75F
i2wvUXqKiqSvh2V5qWTwZa9YsGVh4U/IDhWzNdPM/9QDDqK8xtGA/dyQdUwzmIou
UNAiyd4C0to6obX4P7LefqqCApiYpteGepnyMUyJGqjGeYbyxUPuSm9fRFFHehHw
a7LkUfxhbnaKF+v02knv124tZXhC6m1+76w1QWotWf2MjZl+kD4y59fMfwqeWzYk
SmhNwQEUPh68Wf+rNugovmeJXOO3dnx8zRubjPAah1jrspWvWagdBEiFr9ze5hL/
e6pC0pSU6NPqwajslpKnOKnNC12OiguaG29XzKzz+soAvC9vmhvMtDrptWHnSjwk
BTx1xUfFgGHlhiljN1pTT5Krcha4Yxt0DZc/JyS4jk89JsrpBWYKq+MgCdxP6Jk3
cpdRPFyd386338kp/zwQhDy82EjamgZFwq8nJnvqMeBRU76zcFAPylGOT5X6nv2y
fFjnr8gKkI4fn1axVeeWiIaAgcd58woOeoNuj70q2aT5KZxwcdmaoYIuvh2aPFaF
mL3YGs3aj/V0XQi2b7EeGzx8GpizXtMawT/LsQtjsm6GtBrX8Anv+GjY1/QSqDkn
Xr86YZtQF7wFmLyNs72wrwD/GOZZuMfZ8+TEWCc+nnDielC839rj+adMwTYw8UHa
tqmAT051iZI+t2MDjCZTuPltPp+OJfyLpsgtwq0H14ap9j0g6WGFG1NHUwjs7lbS
zNljPCSJS4A7hDLpUWvFGNYAZXejn9tLuZ1eDaoDM0sJu5MBtao5mUCsAFH7PTLK
cH4ur4eBZFPv/cA6SsiKD/MVcAHfSvmnRkQolKjx2sXDcMnMtXWMBPl7SgKdj5NJ
z967znp32SsG4w6IYw5EbFgcVSjXeIr7mfJIOBSZQfzyW8KZ8gC82CT0b+Qvk6Gc
dCBfRtoJg+n1NCJtDsdSw9vqwX95UPCQzLGOFP7LmravXsdQUpXMaEgouAkZ1QxI
NsBTTjxUCyCzMpPamEe+OdI5QRvqji2ftZK3AU0AWT+WYZMDPRwhzvnF49YZTPXy
EA5F9PEt1nk7f0epNOiGTmIF4XWJ6hulomcvyVns6IfR0ppWcF6nO6CIzePURpgi
EtFrM9ybh3xEEGSo0dQ8XSXDkGoOyTyLFdoH5SkP0FXtbW76d/Gjef1hfWQ8/SNU
HFlmUgASYOhdme+l3WvgG1EZWCW8S4o0cMSNko5qS9+u0H5vuQR80AHs59OGTZZU
EVWQS5GXd0x1JmSKqWVri3P6qHHC/uESePwYhWxpdvv89X1+Ch9vRWEq4euh+AbP
aIDxFjYCnPdh5FLcanWBJHn4x2JHFS6TNueEDiGjtCV6nq+mYAz4NGbIsmV6Mecx
d34l3PffBwzCeXeKm1rq5oxyr7h7RX4MKPHsbm7rWFcv3cHNU6Nplxz4JVs62+rj
Ul5DS9stDcsCERztRopHe+mYQMiF077kId/2xEKHU3m60Od+pXKCXhNTE/o3qi9X
diNlJl8XiaxJnhoX/UpI0PWUGZpB2/j5ctX2TDKl9ATnKyLJh5uuGahPu9Yvpk+s
QA+864Q0zDLg5pq0NfKo3phxtzCAkRI105FpvBtpoNuHcwglWanyRXA3rU/I08R4
oV8J7DK9DW2jt1/ThPzFocU5YNFYmPVImgLeuhqhMKZToUD1/82jlbE/c2tniJc9
+bqNfslKDeWydA54zn8ghl2LKbOjKJiIoyUmNZfZRfOTtqvR+8sVaLfxtaxqzVPA
V2qVpPPJzSVSkF1OzBY7HHInlKOqyNBmThsKE2h9qjNcfLcSVq0EDDdhCv+mVaxK
U5y/hA/jCE591Hw6w/7QGGQ/wgtyFL48sO7tks/4euFMjSLoo8gFyX1acGMsZf3c
aRJNP2o3B9WLl4qu9hXhq97t8II8E8gRzTeBv1tyHX3yDwibuJq976VO72gzwDF5
rKH0S2FO2CimXY9fQFBXpA7N991y3JR2VpvQS7YGeprB0Uh2m36MFzCzuUZT1uv0
Nsxc4wiEaJ2Bt3CpUy2ylcB9jVdTHHo6H0WVfXkX1guCppdgCK9QhQmOzb914T3L
7eRZrcjd4j4OaP6CL+cNkUwvw8eN2C7Q4x4NLxtMx2UVEiO4m4ayHX6nVf7pFUKc
oAsVN/9qqcjpNNwXZ/aRHMoIwhn3VhQQszjPc78ph0e9wbvQzfwUe1ZfJxInmvjz
SYm5bW++H/7iAPddJ/uBrHPggjSFgY8dNVznpzwypydcGWMr4DBTO1O2Y9I7dxPj
2EIXiL0aguysyA6m5CzK//GB8G/+dg9cgK6NQEehb/BYgzBprjrZCCsKjrDQJOnY
T76OuDG71xy+xLrJtyty/RSMiPiKrCSrYUM4rU9tVcflNayCMb5GlzSu19Lh5KTt
9dFlisuyifnmmB8rhff4yI8eiGraQ1LhOJMeK0e6/XZFbUCuUJtfrLRJagcN/yNt
4ctFpud3Sm7a4LnRy0uoszJf/Kulq51BuLMhmjguuNSRVlaqei+X46OiR5kVaKnS
gKRlJFyGlLJ4oSt9g2kKw7PNx7wBC3bECKrb843+1wQTQgqGgm8AIshAPcliEfty
4Gxkl1JX/o0aJ8OmfDqAItCGh7rKayo/3Vxud7uQE9Rcfseg/MzgiXTvnqczve4i
1CSIF5R4wo/miy3gpG8rRp7I0yMclRlRIkvCMOKcZ6Zga1p0yozlgZesSfT5/tyz
ZpVQaCbmfOUB44Ok2eBhyZCB3TN1Y55ODi6wO98r/pqLFow8QqgmlCPZkRvwurbV
3mJ/5+7BOtkcSpYJmMBZjbjOQDK/W9LmS2uZikAwzshEkdbd/JRZu/9pCWB0Xd8E
wxHTQ37n1w6wroukSy2+HIPDYexon5BaZaaLCOjKw29zGeaSgEZ62Lmhkp03NVQP
yNSwzXMMN349jSKtgeMKZHFbXg2nBkho4kPcOoPSZJGqk0cp+ti//m46Ii7KeqSm
NdAK7GoFKRjtMgJw0qt9t8qd+9onI361PmdIVLcRfOtSZ6gvGUwWtADC3Cw2gB6C
6HXmO835AKohJxC0+L4LzDNQdvEWgeX6HL/eIxjI16iscCpiRr8b0Gvl/US8hvDh
dGRhu/k/7yp+lWTdvTp9yzF7gE/j4JDxZd8xM7dbOJIGxI2yIUNz93G7Ixylwpol
arUJIdIqKfv9QP31Wg+2t8268KkTQvd/y5psky9FO19qh6LuSYhJFQz+WtkuHuJ4
IkraUvXqqrqcm8+PqDuNoNBvSuAa8CG1czbm+3tntF75ZinvSu7eBQv7QxS7sH1N
DbEdcT5jTxPQU/USTmn1df1tVJSsxv4vLuxV7ucSiwYij5159lIQal/LWjahrvuz
uy6Nnfkcvm/hp8sSLSqNAd61XRkmUSCdDtPJ7EHmAN7JAx8cUepTWn8dq0X+gPPq
ZdADVVL4BaPSCjxS5NlZlkgsEpri2rz+IbAm62Mb+fAj8C+mZuZhH9nfUxurb+o0
1wFzkg9HfYWBgTsd0v/Z/MWS5qkwBo++i5mrHDcKYzlpdlBTD6Ns4g0HSfUnQqIN
6AhIbYyIut4TKP4bqaNqBuxMn7QdjFhKQFWJAq6bi9s7Ohij0NJaUlMPe9SgxhyB
R6j0DAMQDRyHdPH8it5wQKvZQhpouHe680kHRYbNJ5VpfaatCPuqy4BYU9BbQ+cp
GL/He1PXGkPmKisOFvfBh6KcE8ZMkyVC8a+oq1ztOAm7qHQjpPJBAkgIL62oG/6m
nJitsFFqxWoUE/Neit0TDjUZHcT2punktbcdTpHK99dlmqJzYv0LmJKiWHP+qBNS
L5/XESmaSf7Tkicquw2Xn1IUc07gwesiaoLT4Y95VZKtKGERKNeyfPwF9gRdARL8
Sz7VqS3R/fZ58bIGscWNNgQU4fLJeqVBopmJ6SvBsplggJ4qy9qJI+pSF2D6YiOR
GClAsGYY4AvJHvxKrxycLBRTNqp6oXhxDdQbjW/qOtm9E4rNLDTo02LauyAbrHLh
ltOE1YuSgJkkoX1GtTg1VTTT1is0srQ+O1Ce3M4PvzguDfFuPXewl9m8ForiMldt
ed7oyFl1KblvlVS+QDQMWVwojS8zUQz08q00b1gse9LINgjOCyYzUfeD6u9Wbye5
rnaajoIdgm+tbALhVY+fE9L2sTK4EV8UjAyQfvlH98JzqcvrmiF4ZhK5t905F00L
HEOkDDxCouAIwQPe6+a+E1Z8/dxzBMrvcqwtauWc13rmPpK5cV9Iz+iI/wek/Hf/
x7zndO1mfal6fZmM1lgDRn9luPT0BFuA12R9nh/jTbURMjVjL0ITl0WlIdokHuiT
G+r/+UNkhGhokwIt00FaGhmONFj+XiBFuqUv7luQVzbYYduJXLDQIPP9n5Hwz5m2
ykiMN5XJJ52ZX1AlKXQYRE3MZxjZuerHUOOHiaXjVMCnx8XLfSvX1Ugt778V23xm
LVw7UT6XimfFQhyK9UNlYARGIzs6zhLzbULQkfDU/z8nVlgIZAZRug/AkD++r0y7
TwNsBGYWBcBL0vBN/UWkHVR91fEQTRokeD1X3oeWk0jfO0Pn3lhRqkgCrbBO1r5e
vywDIL88wZl9pBfcx2raGHuh3BfeAo6u3IuMn2ZIUUf42YwCTt9kbmY0e+AW903r
nJVV+L7JfuuUjZf4XbdtSSG5qHFslEJLocCNmmdnytFwXimcl/dsL+cU+PZMJRqZ
ApUoDegneRqJLG95Szm7iRTbHZBPsq6iboY9XwAsO97vFN0dH9sdoUEvyY/K6LYs
IiNNBoGoBYEBcImIlMOA9d5+cv1AMyfGqZdw8Y0aAqXb7BcZo9We3Nk4Y/fAIpCc
Sn112TZZIPr0IAYUswKjXAt6XVJOC6sHciwS36IDclq0gZP+3/lvDCk2ZILZJqhQ
pyuu7d74giZ6Ph7r+0s1eFKS2Vu6IJFHNF3hTCCtcKKYH6f5oUN+BAVaF7G6xhwK
qpEH74kqSTNuJGSVeFB4+HFPtyz/4MBKi5Ybrojlwne4La33xUxrSgKeY4vPL7UK
SWnrJ+iXGxr+aUPw1K2J9Ih7sjCquRu8S1Qn808lq2n4Pk1b0o41LrXwYbmTF8cU
254ZegLV75ffCmWm443eEtp5cUCwT2petEFwVKAiddDeUQ+11qJ6KHlJWeuuNOW3
QM9cZ/YFeR+GFvYZT3ekz8eEfGyDhDcd2mXOCLaufxvQbBcrRkuBWJO3YaqqIUXB
SOZ8mhOBRzbyYeKI2ELKquCdETAwDPktDvvleGvXaJUxa005Pok1jd0MLC+klysB
kK8x6B6w/5bIPqyCy31cSoD+nep48EL8MEJBOGd3L+SQ1LJRyRU1rahqSSN0DDEf
8VpAAyw2dGrka/fYK3FtgR0q59F9VZcZOfQpBSEphOKn7KlX+WZVx6pB0bxzamVo
yw6SFBIBSaU9XV9d3nbWTH/eHoTE43NvimhGhCOVnI8pi/t0AMKPCDmEFncjOKSu
B7WBKSD2gtDVRmYXnGtL8l+/RGiAblReHjy6UxUv/n94AexsFiSWaA863g3ZDwC4
o97UScaP/6PwR0wMwlO40PFTYdSeEw7mAANSQR/JlgD4m8AnwpX1qLh5ZbA4RYce
VjGKcz/L57cfwKHRb5LkBf5KAdnXr5CCzcuVLuNRCPRsb160BFKhtZdUY9YmK8Fd
MmxVrqCsx8FHH/q5o1nRmKcft9wLEYO0GQ6ZTYg3QX+fqDdKJc2XQdKgDrseohAY
NtDwTFeuS2fJGMIVkPfvyRLJLrUftCbJo6Hpp3jvOIgCO4Jzhv9CdX1wKS36nmvu
6lu3EweEUyhJjaPYE0NFaEFFkvXpuEV4RCbQlTpdFH+ZWPmuOs00dyhubwvruvbk
YHu7MbmvBz5HpusQs+fTI6DnzwGkiFxG1T0r/JvQ5wNRZWu5gW1KjGwIM3fsVLtV
sc3v+tFPXBHKJPiFQp07nowmtOv/7sWuZJqkauL0en6EMg9Syg0s8PjRLfszXXHJ
WlQtmXRRO7oHHsCPS+Y5CxTNq75Joc6xy9rLZA5qpuzf/G4AQkecgHG/KY+JoSmE
AjY23IA8j0FOGvdwHjUQqrzefSAMByFuH0/Ai8b4j9x2xnZa6Hau7t1X5pF76TFb
5L7nn2SCs1Nm2SRhT3H+PXjBh2ZGV91B8ehcvunVfvRp/52knh+8hgU8wf8qCYZ/
xE6DNtdipeEOXCJMslyL8ejwtTbDIQ/f53alQxVgDqC7bl1T6yXlr/G9J+HAi4Qp
sXMfY+KDmmUdjPBgTctK8eCGcVBum2DjKDB7cAoouxvVgd6ZLUKjTgFNdiRja/g8
kFquBREhjHZwpYjnbz543iOOE9fGi9v1+/Me+bit40vMofeSoRy0kgOL47p+qwWH
jtsIZPmANIQ2dmvOcT+ryoqAAaGNBVAb/6Sw+4lEg8UBuHGf8n41T6CmSbyoX9Pi
I3p/9/tfOyC+kbHcmQO0AAZ9aKYFmUcFG4JLXH3ghwNgOkWlCDOyhmiFYYPxpY3U
Civ7gamJpLL+JCjlo98H0Xv3XxI6MiwX3IfHYdwTX98LyRoHrZ/O8UfMXfhfDL3g
xpIKDBPKqeg/uQag30tCqwvnzt0+sZHheHPUoCG6VOMq9tNwvAs45roIhOkDsROF
e41L+T36ZZjY2GpyLRWDsEB46N+IpvxCdRWmvy1SaVSA7u9uQNLTNoPwESa5n5V7
X9a+oQP8wzr8GEZCXzI1zSa4d08erSnTLcPZEI1dT98oYumrCj9sg5MZCuHmM/4b
5V4pDE2woAt1OaNcUMR9khYxc3hbXuFA5tVwNjTN3kH+yLME65kYEbsi1s3fkeNc
CfH7pleUYrYr1hlxttT9QNbL5y5MlFsWqBYrLOme0Yptw2L4+7aIXXGZyEbco7Hj
8kOP5OAovar3yNQo5Semp+rF72ltuoLQiBMUdlZmHhKdGUnQO3KRJ+gDak564vU6
MZ4O2Vv8vU8mAgzG4UWDHjz3JtcrfJ1lOUplBE2EBO8MMUU3TMf3DA3JEf1M/wCF
8mZJ+9DKjZue485//bBESSLkGQOr4qwkX26NSUzLHn+0xOQ2mLJtanV1oYH+kp78
oa+/jWfMdCj/RiBhJxqUsSyq44/jfGegpjffFXqAlwOo02c0/e6l5l8Iyf2kGG7k
JORjcHjuzaZU/YdeudJD0rb9gjlUZzBKC5YmHpDoNXhD2bUfE/Q0uYSjzzxoUqlT
0M3Nx0VPbtatyq/6XZzwcINkcwNCM+yg6b6U36A/UnBUbOUECqVchOPNSyelu58u
QABxJDzU4R4DJl7c18ZibI13S3j002DAJLMYrxkNNVKZHb+IhxUZfUFsNfNeaSpW
UngjG7Iu7HuDQfeggTkK3g2u+KE9+L8Y/GPRO8S8Fqfc+UuR/vwlxBSAFGHJdxUe
LWM/u75e/s6WSuh0IYh+FFfDjmydRB4bR+CW8T61VR/G0YWU73WJFSqM0DzIJMi3
5diVVURrcErNdpgxY+eQLpzij5d+XQusTFf8QvufPonJUXKjPlcd9NRfyBFKY5/9
m4lzTxpb58UbboWgc2j+yoaxqGr3vyo5jhDh3zxXRmBli/S+LLwoCbBEt7Mbx5Db
hSzLPrQzGDGUrpp0+QrOA4lxwo0WBO7jN5c7WGd3Wpi2xsQABdsJs7wjCfioHDKw
7hDKW7e8xIYaqv+PmiKybCyJfyi8x05FORxvuitL12TacSVRfx7nbLXWId5ftQ9X
cyP9M7iQhQNZ5CHxUomIbVMVT6LhnabeJ529HQxoeSea68QiHl2pTscZCeiqWk83
vr7rF14Dvcbd9gnlQzFVrTzse/N401y9i4cW/dQ5BhpZY1VELvt7iFWwE/M3YVk0
KJVgHmdlvjioXnjdM0g7sgkXtt7ng1OKrXJVTq7GZ4Ui69QOLmuCOIrdCOguhsOj
3M8470l/Hy0sJvgiYTepnVWtMVLX0Lm2AB+7kudsLgALvfPFkt15S5dMnymIpOLQ
T6OvGBxLpl1KpS0VlLCoKampdqpLuZYEvbeWqRwmMiWn4nxbcyjfFrzTfCJA01zK
xJG8NeT8HCcv/OyQtRZKDR4e7wwz71ON0UaqFlF07wtwinP6tkDPXWlzI0G98GQa
ES0IeIejEjIL0OP6RfJIGrpDpvfduDynkL0nmsAq3rA0bHgzF7FRuAIqX89IxBIZ
8eMp38+nuKgFxZ9witi2mBaMmO+dqmclc5/dvQRQOCn/pqmo76GRWUnTlU7dTyU4
UWbzSHfwSWwRP8MiQiLBoeue432Y2lkMrbmpXXnBCUas3tCvXe3yMKOVuuOtPYfH
tknhFBf+2t4uK6BOItXjwONgUS9SA41qOoUqmJCV5BImdt0DSUxVCW6ivyYFDReB
sKlXC5evnVZwNq4jq7XlxuwvVpwJjdloTczGwsRnDpe9+BvIWb6HRqCuS/OJnGez
CstoBeXMLIqrRKqSLGcnvvQj/i/yjiy1gjolKqVQFXJUhj7pEN+RB7Ywe9c5+2YH
GwDJHGVwtkjSkDdXGRCx4f3LmcezAJojUCThtAqlQ7sRQYvdLs+MjQo9HW2zseAM
/OKqCAQ06+qVuKLm2zD5tO8f7ebMLGyMun+I3/OfykWD4542Os9BMZTnC657q+by
xe3aYY5xUaIQ3sta7daEA2Jqqj541yFFzO6BbH6bj9qK7Ic6cObti7VEDNeYpar2
Du0SU0wqbNo1ky/mlvnr9klj5tYzGdtjloOfbenr8RLX8USw746TPGjAr8qjNE9R
E49pxFH86TLo54MUwLQr3ru0sDrHUPk2xvCEEbmHY4tCbcUp+jza7SJai1jaN3ZY
71k1b710U+ct0vyi5FlIDcoKUOXgMQS5UKANE6Jpy5jQi4cIGovQT7QvNGcx7czG
ctYtVvr4QRrYbW4OE/Fq+xWCtoyvN41eisSssUJCbY1M0brUo+M/VofhVxfywJ3q
PWVomXUqoZmgTltm4yHWFw/1WfFvkQVJDaSSkNPFLrkJkE5GY5XuduSUZY7VdmMA
+n+jIvsWo3PHy22KkDlvM78EcopohvSzK4t25GgO6db1NI2OtZpKGmjhVzad81BX
dJ8c45t4Vt+huol4sdlktlzzFXM/PRoGmILg3RClpvfx5hHUSm4yJaqB3MWwz3ad
vqvHhlnlvqlWlL+ukN9JFxLLqXcmNx3QxAPxMvtbhbjDUMfWEZgvZDceAD9obZWQ
GDV5LDBBzidINkFdANul+jCuLbVB3fvZHjpZmPss5G64g/id2RaktY5cpo38ijfA
6gMc8mro0SjILSgIVrSgf/yMuOR8o7OE+DEA69yTEo/QeIiTJB4gSlb+O/KNV++z
TFrkNSbYX6DSgeVdT4z6oTR8uNIITXqmgfJ3zbQEjx1KY7KC01OdUaoPqG13Pa5n
i0fZr3TssAn6uXv1n4CbMURLBj2M7mpL5F15TKl0Et+iVvYa0hSYZcxuBi34O8K0
vujIQhfigzj/JOc/XcSEtZ+4d0Ei3E2MF2X907jyImF8NcXTbFEM21vRV26mhSB6
HjOvx3GhAMqzKr22NPZS1vYMIPFZbfyW43UNHz8FAP1qyzmMNVnuNTeif0f8wzDm
cnLKxjPy1ttrwrDAfNbJtcTf9Tf+9eSwf5OBT3lHhqtmxfn4GilKA51pg0OA2GEA
oKh+HNAtc+dwcN4/aYQaPh7FLHg7LCeXPVqDDyEmxm7QcUos6qR9uDjV9Ugy0KBC
xff1r8fJ8emJMorqswJ4CcxIas1aYROOG1Lw0vKabuy1LBKMwl5oBGlrfKv/xLqC
i5C5tnmPGTbYqs0qH0SjCAeYnrRvDBkniRS8ccBTqiW2LzZ+uGK4i559nHZiFben
C4OEbuMAxJrIYKD2q5D/aJ+e5dkrz6cw8xy466darw5TZYWyw+WRG+LWcYxcMTEV
zQyffNLzPcp6WJ+toem/ZjZ/s6liR7zV5eqlif8s39mcn73qTo3g5J180AqaXYmj
j8NSJwENgBt+nrk7uHNnVw7QNgqtZRkGb+k4R+yzaVnO5e55zWLmk0JmaYqAMfxS
J15Aijt7JcEzAsifngvJyEMMByp/RvUJe2BHkzqcgRLa1T0si/dL3HaEtWAcC4SW
4NVMmC9MfMZOuF9dftsabxsG4Zct0R+4+627XAZr7vY8D6gh+MiKzbRAFoywMihy
NhcVfGCutZGbQmDqlnyD6ofodGEV7GFkFu0xHQsfdRZCbx6MQ0DY7F89f+Qm9KeU
yRak0dx0O3t12VfSAekXVZWmdxlq/BOTfO1gudFZR0/zFcQckIv5ZBiUtlpxIAHq
1ezbE6yTCPxRf3FQSKtv0xxe48l5XZWyLN9sUfjwt0ySrIYg9IOmWKWjf1vTLgrh
MBP1l2U2NGVFCkU68IXX6QiXmKOcvE3eDUmPZN8W8zCAD46kyQ6LSEV2fJPPuveY
qfe5W+e29TlQf37Ne+oV+KpRdMvTd3kZtgP3XKEYIvS9roiKmS8ClwNkAakTyE5n
KFH8Q62NS5G4ym5MI37soFFR9uqE6F6PNXp8rJ3A1RunnOuyfhkTE8qauSvHSTSs
HDqXKCXb4A1+SnWjXZhoYGPIIl6bjcW6NkfgSNaxy7uo7UxAwQlYApwCBO+BYgsx
FdUpFcYB716QmKptS2zk2wTmOYV5rs2aN4IlBu4KfGeW1+L59AZ7Q2FAtBN8PoXx
fzLqoLkCdVEgKCMMcIwpM8vJLGvW0g8qvHMvwsgOAHA3o56pqTYhbB6MsgzJlAB0
2vXuKpu6cbKIzkdwhMGiTMxrqC92BolcJfydw17nE4TLtBTfT0uyTkdkiqCboDlk
DY99XPLwlKj55h13zx7oWUwi6EZz/PvdwjnBqmA/UcUvsc3q1WErwvJJ15JMn+S1
GQDhaLA9WIVq/e61SWY+6bPFBvjI2fwp6nSiT0Pt/oYTCaT9PeDDiGaOgeW9zQrT
U5MlE0kENvkcC00w5FPoPonDjt3KUOlEriYi+AINq8UTdqueUghxh9/yta8KpObk
IeS5GHDjh7mL2VV0ZZK3eWXTZM4RV90r2bGjzswQsdCkENYzl9scrNQiwqBQBIiD
SjKybW8XZbCqSFtDc5/HJHXrsgai6cCFNjAkoadeyAjY97aRXTex9fNCxUcuzeiD
lIRVcSRkRCnh3oewaBxNAW75Rvbt13d1PpxEhgRJQoYY40iNMpmhXPF5SSu5Fhm+
diCa+K6EFoUi2e6ml8Ialk9KLvgYyS8UAVpOLHi//JHj95le9uv8z03S+fWZ0TBY
06Z3LVw3N+s42jMi76R01bMT0CdKnGlmeF4TbK6c/xYjSBYE5wze/jJB1TQuiFix
oPkxiNbdfbnuqKJcXX3Teeleiltri9KAI/z8xqXP7gr6gQQJgjib9YkFD63t+NCN
ENhiVB1PfMbPNiku8EmQWxt1ZccVNoqYFqR3fS31yw7YvZtWrdVg+1p9bR2jhHbB
xX6O6OE2N4ChifSa1guPvtdveALWKEziXGqJA4VBAyAdELHfAJZ/yJdO4OQEqtNN
8wUS5DqT2Q15NK/YgdimVZBQoV89ii+2OGzVRDjFX4AWnouqcoGHBcUezAKj7r/P
f3qRoTZgtSQSCwkbcrWeiwPat0Xq731NNFSJ09HsUkAF60BZuEnBASUqJogDdjiN
XGNlvFKIpQ06JUyrj7KLN57nhueP5uflUHGpkyCC9Z0LfHK4L/yX1C0B0u23+9EU
XdbcGTQ1YrMD82FscSbDPDBMrd1zS1s3CT59SvI71UqxgTJpbff/pTdkWxil5Nrp
opnNs7QVbxEcc9Z3k3j6uFHYXwRCkdZ3A8loaLxu04+j6ZOfhXep5hp9K2+VxlpA
I489rc4AW+Pli3EKYUHnwPr0JK5hyfqzRY2QiXUgQSGDUF9elfIzDBmfE445pmQv
V2maQNIrFun7M5oPgJ5YiQFcBuJ6Iw66ZC0q3vuzukuu3RUIHwdecZQxQs2WFGg6
f5HjmnJdafaL7vN27hsgTgnigSaAWnqutTW6YuNOVAodGFfSsAFFx1vbLuUfHzEE
zgtxyZsNCsfTNszzbwvC6T94j/AlItklRE1tyLTVZdhmsm1N8nfs65uzBabPMpNI
qqjeBr7PmTo0pebwXiVgEXPxhXjiULSYFx6zvoXnn6JfrQgay12OihaRvS6wzg5V
WO8oI3/9g9+MUOGwitBKx534OxpZG1IbpE1LBxSLRTaHV34PGmaLSTLGAXZbtDcK
l4mH/UtT5ZISWRVlSdU9Vx0rRRQ8/4Qezt6B+gs9ABo3/izRSHc8aD1nXxpADWrr
HnAaqmObM/OZa9/RwGlpJot0IvplD1Vm8Kq+t04aQVy5cUwjqPuHXmHc1FKaIE/v
uyWLe2vaJ/lgfOSjC24fuAnk7VBzJJkn4FZmLCSCL07TQiJzTNj+vxIv2D+17RAj
rRF5Pys+AXDgAq3yviw2YScKhmXDAo+IwU4MJkrv8+MLRrPVKspMe8jUyWIOnk9y
Qcz7XYI5hCx1gUzmmus+9htM64nIaVdbUlgbvGRB8rZdJP4ajLGM5wzMGyYTuVrh
OfWa3YEEGftCVZ8EOtmyFlpgVX1zibbgz9+w0VeFG6mcO+VmP7aMCmhq1H8UjZmZ
/5TBa1/+8pqbXhm+oRK4KaR2EFb3QqJQ9ozFYf3oJUyz5b4uGYWvrToZ7fuNGM97
23FQmw3VBrZ0lR1hnE4KUGhm/3ciE5sHfhZE4uR8rGaeUE5OIVLTNPIhBrnErV/7
5n7VJCITtN6ZK6ZN1bgxDau71AaNu5B6EmGBnv6wqFLkmpk0qOWoXFvVMkkpoBq2
4B1psWaIUPI7S42aeDqARZ/C+R0N5KZIMjFmi2NyUZN7defdxW/9WajRwb3xwA1Q
fz25t70SvlDoM5bTePYjbLSOMpOtF6BBCEe2MUkju55o0gfxzMEFEP7KZFDHip95
2+2rSFfhaJ7YulClD46J4DIwnMlBU9b5my+DaEkRsINVdy9zspuVrh+dFD8Sqf+9
hLXZspTs5YlASA1d8ogDbZbhDHOBJQLQJwmIExnQGDk05XusXVGqev3kA/zFcHwC
KB6zYxaaWndqZPSpbN56bIYIlsCoHhWaeP/5MJhXukFJNZoXgkXjHkfVQnE1ooyn
0ytZ1eDR9yCD9OsJZrsI4i8Bt63jzQciUVTx41KM1OKNNPYfknLyF6ghQtJnlqjT
Kze/eXPJD6cpyJ4CYN4nOl55+4HDLwEScGrv0zfCsz6qwl8OcuZvF/7JwMbw/HDT
RJpX3tp7NYo+hkdxOC8mSB1BSOGgmtuhS2wcDryV/J9MGFaqXnkiZUZXLajklmGA
B3nPBfoBPGjCwDWPvm6vQUTzjRi1a6TueQ1B4VpzyS5LpHtiwCfklXpcbTq4Ed9u
Su7jvpv8YuQm1kagjf0cn7+vFfBaonU8b4dTQj+vnYigtGLNcpLC9gS/+609W2ts
r/ho/Jd2hBYPWYHSlxnIA3lY5WfGqza+F6CsKaHA8k4xY3Cwy2ZO3S7cqaL5bAmE
1zSN/9eRix0bTerXxjH2Vocis0AYovPjb9yFtnzO+obKP3AMfjThW3raX55TFqgb
/YV/AtdJ4wYCsUSuE9xHTPc8/7UO38nulRP07XWgsfOl/wXACDq4sr2aDnijwC3U
7RobWgNm3uwUliuoHDpsJE6heoGfNgY34Zlz4OjTkVSCqH23x/e2CGDjHN7r1VMB
832bZmpwV3+Iy7iWftjN2vqhakgG/+MzRuvH2t0jJH4fIMWDXHRcD0IaG8Enpy8S
uFGaR3NBE62ckebbNZts1+pQ0ZfNzekaObuki7S84e96uuUCUsGeRUrH2Xc1cYbQ
S+zVigziZHIB6e8Djp7p/DGGiWYLM/OclXJ7qr0KMl/Jwx82Ybnn2R9IddDlyoIo
w1FrMxOvDBGmK1zzAeO/6+mr8t0+xnLwqdCxYOCELGKiuWFDC7V3Fd6GV97dKtZO
+QKvose4r1zWIyT+em1xPn/9zrf29TZ5dRZqDIGxa2arUgvOEvCS0qnjnHlSEQWm
bdFOGAOes4cSBll64r4OmVDBiDbiX6i78ysn2KYiy6AZ0O1SGHxP4QAiYBLMKhzH
hBUzzIst3VVA2+F0w1WIUO3cAQoq5wuN9S87/dL+hxAedlIh39PYrh4yvOAC7ZWK
mFxbqfKeKyWgmkR74vldILpNWUlR3Ptf3t966qzu7i59KZyzps0hDX60rtaeQJ8g
7U8MXCOclFJqQw6FJ4KyxWfvKIQNtARpAAtiLvCpdgbMMmhLrjfgHdSI15wKUY4S
qn7aja6kax+j0Qp2KUQ/ZzmTcvp7YywNzFM4sf+5WDoVnVtvF9VGa9fLmaDffgov
1PrtnmXE3eVt58i0Z3kuPPxM/ttT4MeWQywTFaKzQ4IhPeJ8LQp2h4ZWk/AikETK
Foy8GUGEmJVzHmtlncuFwmsZ8VLTilRMQuhozGTockZnYxIOe0uQUUiKtDuN4rfv
8EzynlsY8iS49BzV+LuiUgaIUUH1VMMnHA2W1ElnDai7ZKmgyKSk/AW6EUzGT2NO
EXzyVH/hY0C7PtbawJU2lscs8bqAwcsXldOWz3Kso6uzwt3VSay1H5+7nX0d+b0m
cRVK9W3r+DoSRveUFqtD/g5l0lg5FuAaB+5oXPTZlW/uf9CC2s69womWVmfiVD0j
CkbplDm0G2ndSjIa5a93pruuCcz0ny1NSdDzj+sba2qQ6A12qBQV7kynQAHPnvAe
qoI8vo+H5gtqUWZ5wX+MMov3CG2xSL/ap1vFVIzjBUd1khiRe3H9foPDyBmykJTh
8otC1a39zusAR6j6JXqWBIqT89xT0xR8a4rMr6JLbbIl8bAUf5WKCZHtlIjVLVuf
CdKSAb1N2Rmifqkn2R3+Rgaj++miGc71HJIdt2fmd731haCxhmolLVqs1rALx5ZX
PeJTXKxBW335wOF57j7QljzS5ct1xSpOTcXObvMJRkOxRQthwxtGcOSzbTvBUHtN
wPscTmzMHu3uF7paU3hXJQY+DENjx+yZ383AI5Ey4K0HQMUv/oiZtmyXJ3rmPRWN
QT7YJqLtF64ncuEGGa+oJb+do6XMDull4wGkLOjpFpBCl1d5QH8WNjsiOC6kdZf9
j7d7LmVP8pjaJEEfd/iUJ6s6oqBFg2SYA4YUnhIgIt3AB3pWzX1P3eot8HxcfIDV
BLXm1YHw847J/n4fT61f7juj064D5feZ4OsP8PoKeu/e9KSTqGs2UnazmO0hkbUW
hPBOp6MId7FdmGVrLA5QR4knhK6OUUKfiOyUERCDZ7a4hz8ph3bCEF6MMt1okqzo
Hi+vih72hguR4oYUWqATmc/M3S0XAqOwAhQoRQVFs2zlHm9VkklVKR+R8zFja4HE
/cTS43tEwY3r1Sna9rUEPWU/dQpqTig6wtofcmHUYzMsatFeXrQGqnI/hJ7EMN1i
W0d6f4vXi1QlTv+Y9trPXB7gtdyl5ZCI9rkf8KTJhtoKdGXehiEdR39mPpmM5wuj
FC9NiZ0V4UWh1UG99F/DKr1fmXcBGpwU62NHBryl+l3dGadfHdQGhS+c5LXdRHuc
F+81Bu2cYYFdwN0A1w+onleB1Nj3nMGVlhTa0+WSQo+qKhWehzIss5hP6nFtJXLo
MzLLb1dMqa1t6L5Oe6LqE/HNs38heMPVpe70oshQApzb18J7cc526JxxoFW9yAez
ZHBUkBnP80FANobiB9HD7+9rBPm87ormtxcLCZ3CKw08hFo8aOruPaASXpFDDiTH
GQ0C+50jEQgbo9wefFsPAcmvgkm7n3NMJrKjTQyxunb3+827CFNMiMMXWj/EqWES
FL9SzLyKTVTFwRmgRyGCf+iKwIFg7nzHeLMRytsJ005WHRTBHoyzVo91a0rwgupm
KR+W23MLlHfy2jCTWX9970wmw6KFLZLeTlWm18uaWg3z3KFXc7PAM0vmxrq1f9Ps
eBFtHc48aI983saufTj8DqaFfLUdI4THbIhdtVuwa1qPNdVCiTwvhg/b5Vzr/fw2
tCfw4x+/f+c7m+gkqbFCHTyxbHDRsqtXyoK8ZXteeIXdEigjX+HgIPgi186FTZmn
CdaldPTjIGc/d8sLBdpOeYz09wgxVxCvlfbUVO/k8/k7kyt6RjaRgVST+Fg56fg1
WcfY2Mj3wjx1caPcrD8w0WRP3NHFGs2nwW41OA0rfcZkIO8eSE/0hy+lRmF3YT5V
kbBaBxdCF9DiJEeT4zQqaCWmQ8xY+hrhn6JcCD5gYCbfch50OkkHRd4Js2d03ekH
e//J3JKAqYFsaDjK+/iznFoO141Qc1spm3UaErdtkzfLm1Hl2cmqD5trOKA3Bdg1
oyrMYKyHVc9VvRLBq6qyX7aW148c3849KLoS9UwRRGLpu/Sh7CAoJsAX+9RmDXZV
A+ZuJ++PDMnicG7MDnWoDKlT3u3CWEe2y8o1O5FZB+5zE6T7y3LrsGDW82XjxTkw
gippi+ua/YSw1ZmlK3NwN58YaoS1oRCJrsVB9siLxpQ4nvMoT7O2QretTru+HoMA
zqgys1tioFDStBpklVqpzVG2IrQSf+g+8cZWQqJyOxl8FMfJ80SUSUNqsc2CTIMt
BKODe+8h5tXyB19TYz2L5Ew3b9iuNIOEulgUIyZwmWb7065m8O9l+PKN8Wi69UZT
rTHLH4asSViUB3scUP/L8CrnsQ0rfe8jwthn120IBHxX6CGh4ZNm+UfW/TEGPKti
o09BSMBI+xxXnVPR/fBRgw2cIIbBkO90QMSl1ykoFqSihRQEyrlYeg1g9k6LUmUU
yewACnPEGa/tkN4lU5pypUBX786laC4Mxx5FAu1UvhCyp6OVpQ/CdOLir2zmFTb3
0WkwIZLyuTaiaUSpoaBJ1fpmE9pbb66gj63ITVpHgMsl6FRKkzvp6nG9OjBcNDIk
Kv216aJbRuXxk/z3tklXykxf9wGxZJfRnYezioJZfjnol+eae0u7ufEf48GTFkSy
CMH+9seXEShJgouY24AtBc3pR1SJfsKLtK6GSa1P+5vrm/0p1D58m/dDkZQUg/N6
Rw0dueVsHGYvelT/7UnkbwYrusSv0ompKp3Y1l4cpFA8MBzsv2gncCajBhwKOQGC
YO8H7BCta5GsTdmVZ8z5mBxoig9Y+fSLeA6eHPDBxRkhjnd89T6jhno8BI8rYjf9
YWBYF3w2Octv55yu6jVWHzeICE9rGkhRM7J8FQNscuTnFA+04//lh0xbmCeCP/D8
YE3tJ1tNbZaWGu0YLW2z+Uvw5WtH2hMsecljSGdwLrGwCnCJo0Vb2HnXREPfvyXS
aNmiDIxT9J32IitRx0NR+CsMtENtB9T938tYSixZUxdARSEWYguve2Yc/877L0wF
AeolrD0dtRi0E/wUEV96FCigaJMm+4nu+QrSLKUD3GBDNpbcgCZUhuQPIR7QD+JF
sNOgQ8LaqYzJbtcaGDmPwjJRXWzkW9AK9VU+CLetIsFFKb2+ed1fhRi7mWGpYYZe
KzMn/5dXjufUQkIUvti8tesM5X9dluI4v9WFJyfpGBKsyRcA+pmJCRvqpLMVRw4L
dc/6k3/Y+7Xz8WeZhOUERIs14md9KIpJWNM4oPlUhZbpDaLNC9mrex7zMno7CZKp
Hc9jIAoOBZtoqaMNZEOGGsFPEMgnIg7gTmlOXU5H5KxadKhxR3CFohS+MhMoVmhR
Jlk4i+siM+QPoU1N2lYJ902dKBxT6GEuuw9SSme9xkhmcxcLv5JR/Y35VgO09x1U
yI0rM7Tl+V+MLks+m0N1X3Sv/F5K5zdTjcCOd5C8OWAWtk1Kru6DBl5ZyuDQmL0I
u7psLf+bTJyuXdQ3A18qgma+5oXGRfbVrfY1wZPrMNlW3du6/SxudVnARPNQepFM
XGnLUE5n09xHkh0O0xYbmrU9lJvli9xhfeSM3voMnVcR5ETkYYx8M+7snoi0vSjf
pzkK8GgMoL+kT8QtNKhMqEJ0DCVQtGx//90vURBtvZvedSjq1jX2XGXfngfdiAny
iWhWgXnJukO7MiLqKrCMp2FxzlK2PB+dP1HEeak2cMg/2Z8gjMu4tNBrJgRwAeYW
qGuqC+umbNBHqodSJCnaYyzYRnrZiL8/lrB/e91kAPhs33sqdiEd0wGBUTzpslgi
XcxApa+bfyXYT/mvB8fmjmpGKw1M23FJqL1ikMzhZaQaY/oYAEeeKaBpmydmClDL
0VZ8nCrqNIxCVjJ8RzrrnZa25NfHmFuBzzdAWIySd80mFyGrhTn8ECBlw4nRK/I8
k3L2jAsKrQ8jdMfS42n9pyXr3x2rUkal7Py2GciwXzYbtNk0r1SnWjP4DWTWfgB9
TbvXcHZhFM6l9FsNh9siPY1WPlfd2Tj2pdaaVFBi9dxfRTZiDFej9Fh9R/CdH+Xh
b567lLzf2HTl11YemXgwAoFr8lLUkrhRI/nsNNcblBOqq71UxQrSP3GmkMP4kDc8
9YxdUDVydeBkLgOJnpEmB31gHYshsUbGxV5W5g//sj5Uj2dYwBygJz48yJy929am
m5ToA6Sk60eNDOabjd2MHEnyvvq0s46fav7QXG2aO+wOlZBRPVUc7bOdSbPd4yMT
uYAyUJ8jKsh4QcM2frGwXD8dgJnGvwMMbVelKNVDLaUYF/j/62UzDWi0EgeOo60a
tcU568uN1y2/LQshe5x47ly4lRiMLCUmFS/kMZttfejhq49C/iEvwZHRDSxZri7m
s8Vog7kRIxYJYCLiebeqBuMhFlzamWbqwFsZV91/VAyMwQl1tlL+TS06Gagh7MTf
HGHFOuYyVuiIiccKbF2tib42jp9nAPL/egP0mv/U/AVfS2iN7x6+Rxa2Jhm3pGQd
f9HwpkkVrl+6O+gsj0vP/24u04PjRgugs9XYyGJvlvOXxrE6SOJqZG1M7yB6UMoF
f/w2idYfwjEPyI69L0eGgLgueQkzaUtkHadHPmVvojVVvD1QUm33raqR3vNXnHLo
etyBoNiMwORqT3NcLgp4kyMfVdYN7O5Ur+/Ckdn9hMPYirsolPrlDINZgNtCY3qT
BuI0R9nqhqfinQL7BXOn59QHSzKDuPxYevgCArZzGYF0U+ZSLNCEPnirGFQS8Jtz
BsEFAx8iu6/y+TaRgXmdL9li09YYMyxOATDcur83zCaHQBFDyuYqQgJ8KUMgdVkL
gGCaJccli7ItHbBnR3ntbLR0+6BjEpAX7AwRFsmr7/VlqtPjYxTcKqi0ppiB5vId
GeD0nIs+va3QV8B+gyA4OUu5IzI1uemxY8GKEBLnwm54eurIut5kCDpG0f2InyXa
GVKgxO+Z2aMngLjk2U7zIKqqMjMEZeeMUzwZhO9qlfOK3tPtg9c3Wv+XMtDyKLuZ
8viMHY5T2R23Mc0WfHvSu43eRssQj922CkrJe9TyQtQGeYLadHR3yXXWpVLBp31Y
+1cXpfFCcNlvdN9zIlU7f2iHIhF2y7aV6WjmUOVqIvWoy2oDYkgJ5FerOuitPs/O
B/xrDqYNDrQWADLFMIrm+XSirk4rtnW8BMHkbxVkAvuST7dd4BRfDaBszsuIwuzw
rYhRI7nx7CkirBEeft5SoPlyma++FqfMFO5TLnYm+HPUOOXgCQCwE4i4O1LJlko8
3VCWAKKxJXdCY4LbgUT3l3E0yQ41XtaWKsG0V0WRGTpmRpIdGTIPpjl+ttZvVOuB
O8w+ty3ASAWs0LTc7JYmeq0KKha5qEgSpwAKr5KOi2/BncOlBxplyxQxtmXnLnjR
6y0/tjl+T7fXEGWNibH3JKo6UeMys/p35oYnD5Ep1IJB9AGqMTcX7fgRP6TfhNxK
hm/xVeNwIfp4kl05ATFHi2E+wKG5i0JoLDpMZarxGWLJbVfYT0S51ZTg3rlGzGiz
Kl5Ch9aq7N4OcBaT/TM21cG9OntEjxmt49LqXH6j1JAPtC/8IFdVKDMoOkMbjD1n
XZrwGUsCEHijOsLbDLjTLKbZuAayjaqbb+ndFQMss6MxeNGa4PitLBaV+yXZsfOx
Q9CV5DRO5vdiZgpHq4KTcg9VXASvvOxC8mZDKrtCeWOreFkna03qB0Ig+1NPcqru
y/8+EeUYoUQplVt6K+Ml/KrUxMeKE/MQLaVLwfcvivoRZyG8qCsVIbbRk1UtfKBm
g8RMXXXnkIFCAiESRHGFM06/vh9h+TYUreReA3SZPRwdAyjP0oucPOePQ74niJYj
iPEKgDm3EKkEwRvAOiws5q4qoPNsP/svQfWvfeT/bKJTdI65UPoum+OZnQ/Tj9Ga
dsePFY1VkjPwJrKaTxlSz0wrJc9mA/7DJb59SO+TdOBZi5NwLiiscKUOIJxaq7ML
xj11da93veW5PYyB2keUlFlKcgRyzoOtYZEDp/3CjnvkphfdKyR8s3WevBDpXCvc
qNJwti5Y+KYIEOJwgaHuXK8ZRQhDdb/n6KH0vANi0DETgN27gBsoSKbJUKfo02JG
/HcDwGdHz/2yb2prhqRwWM9si/7ixBUkrWzVzUwTb1A8BD29QJ15Yi3i4OIimpkj
TD1cH0KRDL5P4+ctVdX2YHiEnpYqrr7JZ7GBrEdjI3YMUSfFS+Q30mi4eqNOuvdZ
707IHCoDg1/VRLhRqFJGqViuXZo52At5Q6MobikK4h5A8jpdb+eRpn92fOUUIM7p
7y5r/keLpaNgtgFEm4sJYujjuptEOOiT2IBDsC32ri19pr9eRxr9ic271ZtoQ71w
SsUre40b0vLdAwjz6fOFwl0bb4Yx3QlHfJS0l4RMu4qK4CiIAy+IeCAcX1v13xNJ
Pw3Rk15TMzcnhdhUs6z/ajyFmd+kWFMwaNgZ42t31IhmSEgIDS2Mubq9WgPq5Lk2
vfCFsFWbIJkA/zhfILfZ5jGMQN/5x+uqiuNyyS3rQdIZvfuZpaF0RhNd7MfwhpsH
Sg+X498Rr/qeWkeA0nH44S59EkPLb84r36tSkIpDxUpWh7n7CHhbM4wSZq9pISfV
84NYLsOzIl+eOoXVI+KKI77VrQlVFxNHuA9aKoYyq6wzS7eswfXc+Sp6Ln88B0yc
PShG1BC8ct4hKVQt1OWBLIQ8k+HSGig0moCMfBCne8tAXeSNWTWFraaL/KatDRpa
i0zqkN0nMeCvsYup580YWX47E/JhcUs8eALT7x/gVY/sdgiR2CWFA86F7Ttwn7YX
YMslFepYI3XJeHWnwziIt+HWVHAExSf8O8hh3cFNcHBlClUGyLAndKjmuCTLlN87
WLFgBT8pGkWhkx2tF1Ofd0gCUxWqbhF27yHh1k4Ej8SzVDf7Fx94OzfSoHr680bL
CjKah0hBExWz5juhL0mhh4xiIKlcWSlLH24fpBUnJ33vUjioxmH98dpvNtfQ5oAD
l6NVi98Ngb6SWMp+6ZoJns4frrhp3BLN+hoANSZEiRcO5ANP2JpsIB01J16WSZQ2
bkKBB6D88vQrGpjkcbUiYnw/qc4me8Hj9Q4QX7kpnQrSwZHt4rmYLkYIflHVZOLm
DWfAy6c8+AJeDdpCWNeSWxCAhbHCQgjC3twq+BJNmaRuql7MQOfwn/+OVKkU6j15
VDRKmGLdfdF6A4ZHtzS5CQMmMOlSC2tLpl3pkACFtAF0i3L8zhEkNcRc3gSLUtSU
pVDIhjXJxsfEVwnjXq6JVe8TZUGoDwZv6/E4QFBDFqru+yjGpc9MWMLlZmNYumF5
/A7WtAD0P12r5lGYjiK39nd54z33akNhXWezTlCIVU1vdveEIdGSLKSfdtkJ3KIQ
0nh0BLlEFM97k17vGhACCHdzGkxwND6Tp++8eD5T86y8qcsSkeX7u3Jyy3YSksN4
TYvzznVwptprVe1cXn741GsFai8BbWhXe/92aooB/+SdI4NZStKOikb2GXD61sL1
6jEKiKuneSWVxCW4Kox6Xt/E1V+092AJ1XD1Y28xOnELVDK/g2cQwBCGBDNFrCEz
yiwyX8voev6ZPkCwKrvtprhBkKxRNeZn1L0USg5TZszKHQE514Am0vxiZUHfANhJ
Yz2HN2R5A3JUbaDoMJsYZUHhUepDEVC3w+QnyIQgIr3npY8shuYncRwdKLjag/fm
tm3g7caBVBH2WW/sqIdBqm0hOYoDe8xExkTgO3rUkZWOhlo+zkskL0r61Gas4E9z
6CDJImBI9rwwhrnuLfL6yq6aHa6isMPJ0HY6GKtwywZWFy74LObzGxcgRFvgqiNJ
xY1/T6xhbR+U7WWT9wK4bqmMTWPivvxyJNgaubqU5rtfh65VfCHHryn2ldoXoJ0N
NWKsp+s+tZdzr5GV6KPteEiNU831l0qWENx2nCrH9mLoLxjN9/LZUkTaORpkbuDb
QY8lq/OhVE2v5M4etUpaF8rNZOK5Z3UjbCkuJciWN1nux4p7AWSKukg7lk/kacIl
YTzua/ppRWllciss2/JhIUq/G73Z9EEAfEf23sa7C1TG89i9WB9BdtTtlA/Vf8mv
rHoEx31IZkB0LsAe9ZdD/Rqhcf1bz2CgxaVTuMY8jN/fPBQzu/dnjsBMvUQmXgYE
3dzETs5+6N24ishBShKWn3qLz6tOwkmMHTQ5y/em6LGptBuDwx5f/z8gT+z44iR+
p8T+gps6leLHbxM22kz17hPgZ+n/YFWvQ93i8o52We4o5ieQCBaRZqXr9PJZCoWQ
hsSB8ePbBKpqFFdxvcnMl9/+Fdu6OppQgb/0vx8lyM5nkpkKRlq61QrbWUDZtLMz
BotEsSuzK+obHVHCcwTzKOpHROojY8LJlSSZlYQL+ObxxP9qQgiNZMCw+ioAzh0i
xc8Wjt8DViDN2ACRR0aaSvfs0j6+XcckvX5uqWpIiL93nf0oGbrf180yVXpxfsd/
qUeMGQao+PAsQ3/Es/Bn6TIHVHD3S5DqzMP2u+J78jopuejVtS/2CNldgGBa1pDL
OEhfVU10Bc0JvwYAeOVYwKkrMSKDmyjgc4ccs/Ysu9ZtAbN1UynuDkoQljOJGUoF
uq/iUWTXNPitqQxnxw0JyZuAt6ayorOPmychUd6t+NaYlIWV+GgF3Etpt7XCF1sY
YA6QAs4QPBaznGfCS4aCjav/m7l6qWviwGRNkaPNXylUGURqtE1ALJzl1gy0JUhU
thB6Q6pVajoS9vU/38tHodvBRE2CbqC8lNd9S1zHKrGq3dXemDLOhaYQHUBzscYh
kdQApps9wv0oINS8nBxusRlcHG0KTfXUEuHNps5ro83x30h8TwERvBMnNJ7eeVtZ
XBwWLhXCi0qqEVFHGTjkAIYCMbwS2QqkVYgRdPvvgC8FlxkBTnekSaKZJCioPYO0
04jYJw5Lc+5St9N71hqnPtCyc5BKrFcBY5nuVSO6xeP9edfmBSvM22gvzTTBBL91
em0bKLGJIN6VeTizUTgEXZ3KsH6FCgjAA6mWwkg0HiqDKj4migeyXgWKBM9zWXAX
z0fVpqw1fhJBUqukMcv1cDHwX5QaFrqENa3EIXh76neVTJvkumEMq2DjFTd3Tp+d
RboDoxjqpTF0BQu0ZzDfOffuQG2UkO81PQ4H6a5VSW4rWq64qn/3cOr73oVfDQIF
luCg6NSn+WW+CTD7h6B/GTjC9wPJuYWIfXAgoeM3wyrkd3Vonszg4BqSevVRvGjL
ELQTO9/WXqpmO+enm8FbvoyRk9OGxB6UbrsfQJFr9FzHlMT1zexfN/W01ILXnfwl
jG2k3cd8Jqh9pMlcjXtdpBRNsGHxUs1bwDuBVfhfiVWQ8i/93uBTevqOPb95rI8v
35n1nhGg/zDWfj3OzkM2XZlwkFnpUlSs2Mf064mErUMOIm0lrDH+5i3a0FMPox+a
CNaSZxe6sHXp4hX7hzL5EmO4kaSCRDeW/1qmj55OMfvJic3DpfsRRBliy18hkI/X
zaRaw0wEwl37CtB9Ne3Hqe62c4PfI020m0+3L7rc8vtnHyp/UKYhIn/QLnQnrMhe
zJO6Jb0gqqBveikUZBhlMkqg0yyG0I2IN/iyvSic2OHJYxYRD50l2D+NGaIUvHkY
B5jiwemHaBp2ny7KcHkEWcOGRZhYPcqND5h+hDmGlTd5gVhTiSVGpG5Pd69/Qa4i
v6AYU6YUehCz6ACkMdRSM1SL8g4UOurZzwfJX2TJlR+CGTHvWw2Aid1DJ/uCwJec
W3A5CFPEs0monmnvUl/B9CMSjEC7Xx/TEep1qzUGnikKEBHITFmd9YLNJmwLLvGR
DxSLhofA1UnCIQnS9ZSMUhlCK9z5en2pmtvlGDrAZfmnh8Z3hthJyke3CoJ+m2tT
Jcd5kH7GLmWUVcHqBIYpjF7L4rRFQyC8CbL4wr7Wpuwq9dyHEgSlpWd5igbDW++a
+y9DAkffT53rlLlJuU07Jjx1RCG30Zt3ZJ/x8BVeCxBzr1VY8xtZPQ95ymifTWsa
Ngr/C0JnQm2uCqmQ4dgc4/0TalJShsxcWtsH2OhlLKKt8MEu7Kz+Cprc6XSixb+/
aCfIiuA5NPP/yc0WGiX34zkuMjLKedTgBXTdZ/yPzwtgR8WW7kM5QUaezmYO+DpX
sCV9aBzW7iMNOlYbV3ijYB1drrwj0zLQlrg588rKG8gDKR80u+9FmzvqSgR4SGIx
6BddbHS6O6/5OhKksHtGgJE09xv6OgPp11flXuOer6GJwjq0TUdfrkHNV7JoFR6B
XeGymqDRlCp2cQAK6Jqf7BSm/1aYnAShPxGZ9sypfIA2roiNM4qbTAgTJvTcF3cE
/OJpvPoIphLpG2L29l2v3wpIbaKUSaDL8IvpjwtxMnSvDs1tjcHUMSc4grqhQwiX
4GLfzDVPb3UKCXNJriGjqQ4dyOv2+wMUAX0Ju7RL1GA/62flKh5/dNcgTm2JnZcJ
bVM8mzJ0t4NpYZnxYB1xNEp0hgGHadXMDa6flWTe+W3FS0nea+IrjaCriOQlYpTP
y032LESNxNr3QljBYYKy9sDdGvz4WEruYf+LEYtTeOCaVnBtG3EjP0r+8zxg5Asg
rYvq6uqYJLFC3vQZgV+DuikRBi/6HbN0w40H24TUdSQ0dpmaqFNivlvLwZ3Pma/b
aWa/VmtSViMPCiYZWZjoUDb9Z4m3yd82aAFDh0hTpYSE7F/m29ANClltLQqgYq72
o3KgFz9vIHlhOZ9s1bEESkiAcwTbyaKOdg9N/M2z2K7V41QNgiu9JBMER1SYGcTp
EtaL2/AKMdESyKBRJsj0QNVKhtSRRdn6tzgUS7zIwqbXuHc4D22Hkq8bpQUHX3JD
Gsz0iiWm8tcEt4Z3HBUm29G06orHJAnVQk39XA2fXfKMZoU4hERPFyUktRIwYdWK
dVGC7eC4Mru5LiOo6Ggf7ykwNRR6qIPWUF+0XPSspwssVaOe6UqKRTFnhrsxs1fj
HeR5uHxOfADxn+cOUsmADgegR9/NG0SoqXSlPgzmqKY/AV43+49GJQO0iUeCw4ch
GjMMHjSya5DnhhpA+uWh393Pto+EIXrLnni3r6L0JNw+ZngLd2kbCADYR/zoHhGx
Mgz/4aliPEkXyj2UvgdLYUkKjyj8JmMIR1DyyZyfUHos7JxPuBo1DXO3g9G0ST2R
wE7tNPDMwi4hkwOq3iQ3X+NssXPlqzpGxdlg2CrbYCLpoGPy9rarQ+f/7kOdtBPc
j4fPFLZl5KkbTyy7dVq0yRnoJKrzkKz0/oM1gvVUJtflOA81az3GJKewGz35mu5/
5dWsgr1SIASyKMTMUi7MiKOVZXF5T+7m6USVUQZgjkn5w7sk+LqNxz1K5FrAM12Y
FmSiBB4WLb3oF104Et5VnCzAVvwamChmWUW1JaEBD8ANnOp1/VtdeKrPgJ3NjCUJ
+/bdlV4PoWHRdtNLH6/y8+Gm66H5PEQW2NVMTlyzk9rr68bx6QlmDJYSJZfxUAti
GapY9fA484M8ZfIxO+yQDWIpcJBVYIAIPC6I8Li5DfV0g041bekVEd0sgxpkVFFN
Yr4WOhypTR0KT6Uuv5uo1I8BXJXLf11AJDCTxHOguZvQZ1QGZ8FhRj8qjtkwIAbh
o619b4FOspT8l7NMlmPTxjbtfb648P4aStb8xzMiBkJ4TuIL+Ou2gmLRxgmWY0Xt
R1/PpriVtLzZBOLt8ZZaM4Ot3z4hK3+FX6HVyj1wfsftdJO7Cdt267LWZpuEPUVj
RAELHGtNxMs6U6rMwpgA2x64Syibp+a3liPKGkmf6vtEY/MDqYJQUxxNpQ+J37C5
brNekUYobNvFpFjvLnMNqLr6ZxP/MjHM0MNt31S5vdiMEG4nET2Yb69F9RC9++O6
aCDNyCcrTKAOUS4TuDKfvdmt19xn0GWtaC9RMdwRtGeM4XmJOFR1D9ufhxtg6Gry
8MZzSCaXzrsPOhTUuaLEvVsMAOpivRfoW6DZzic2+S/LTAojVBUGQRI74exg1Sjo
o4egs5FUD5Js/E560Pi/P0fE6Nxq3raJ1Zg6jD1zXBlv6WxoY7g47FHet3ob7yjb
MDgNO6dUgMmYOfPvkMDKq2dkPTzSXMKl8B5cOezWHsuV5+6tMfxuimbzAhM2zHAH
bV7+HWDjt/dJWRK4KfP3e0WyLbw8AUD4kFVMdgULXPPGkRQ0A4W5LDxOmJnga6tq
f3Yu6WOVzHyEagcePxD5KA9LnDrE64DCwsLnyySeoniKAGY+hA8FZmjosL8woUec
4PY0WYoBuqezDi5KsfI1cAHXt6yBd8qZNm3gXme8RtlMHem8edn+9VCiS1g3cOUB
IkV4DHwDleV0fha1p+RoLv+Ic7LDz7XCddkBt5s4tqBD5o4/MBkUFI6u9Rimzy6N
tkCUDuy1kiXiATLdoS7TYB+uloBGcxvEoXILzTvAnxTtK+V4/1GneH/1YyYNNwWA
2dR5njmdOp8pirZMAI91/GiWi4CovLpAe/B0EdHMdfRyiF0B/OqTsyztTj0ux1zF
OO4yNB0boVO98kX1+4nxN7HEzZtyCPl4nRCmdD2EjPBHoPrJYNub7oxnXVV5Ygyg
Bxjx8D2WPmshB0K/VPMbwVvHM/9H6rLNifpT0rh089/qq/4ZobkJQI/+XwrJCnA2
/HXrwFBj5ptP7fft0cTN8oTmcYeZ6BCB5xYtEs/+12HTW7w5VyGfWX5r+UiROK3F
158kpRJBjkZ5qO0Ba4lh7dHZtlSIehyOUmYwM8PsvYBV2OlUFHBVuwb4GGyWoGap
Yfs7krq5xZUo88YvezHtG7k8VDOFDoyrjcMTjtHMADjNYCsd4Sbb3LJsiTytXuzA
RjdgcZGuTnMOrgDZ9w9ag8kGqyuEwsCggWpCaQ1LhgaKm0/nGsSFZY2YeSXxXDob
5GuQ8qHHuPCx1ckvqsIgR2zrz5fLybvHwNm8JXnKqOHeYoqpgpDXSWmWgcAxCEwe
SMmEmlchL58iP8pqKlDqRVLMp9vog0pTqs2VgP0IumCl3GVGLDg+9KHSB4jycJw3
H1m7ELmUkgs6LFGc1rIrmWWI5sREn5xvAXZhOKK53rXEwnC9MhQ2jGHZsy4nWW0N
6Vj/fKkg/2vVoDlPesTDe25xIEOD2qzLJcrGQ/Q/lL4+uF722L/8YM7HCUvDjBPG
F5h5lObw078CegMMcPL9l6Sc0yu6wENGI/qVSZ+74q+VY9iaW9XChqfr3GVDi2F9
IsgXhWzsz2Hyki3pXzylngloKZmDexkjv+rwbUJW39wgXepJ8XisQ6gpG8vaPs1h
Umt+QLW526SrNQRn/Ch8KQiyn+VTPeZ7fRXcsbiy+FIefJqeUC8RlbQV5laI3nYP
Zks8AVplXuALPUbwStueQztSDnjdWYO+9vbHowQay/8f98hT1LEXraPg4fEVZJKb
+4cwOpsUu+pYSDr/Fpgtm55SIEPwmoJKA16qlDRr2f9aZL2bnTrSDf0LWlgOmXn6
N/nKHCvYVIzik3DuQFtULQUl5zCmH83gSake1MgW05hytEEC8D+cpjxdNxBWQcTS
3ep0+QhwumMqxwWufHuJnEUwMdGNA9ZBpol6A7OH7pdRuhJ1yZgsPb/2fn9+flHb
OaW5W2SHcKdQzuFcJnPWG7yb88AzI5GAU3Zp0Nj4lIuT5dAbGT1K1CI2u/0HC7FR
M0yr/KEYK0fwwfzYnQEvmeJ1CBik3rBb6Bz4F49B2p901D+DekadKT4DQd0PZFCC
ytov2DgvzNk7qUAGHGgFqMgvT5Wpfr0wLO2d60GNFoWRB8dFWhoFcxWbvLKe8KmA
OfssUJQtKDTZ9RtdDQNTQplrR9DGkgBGO8ye6rbPT5ooXm80KCmUpzYgXhyAgYBF
JcxWtsLUzP7tFNdbN3PVQv7k43+Lw6BZecjjBYRnspWEkUWO5w/WY+UdfKo5uaW6
X0QuWfTelB7LFdlYupTWG5aHGgZwrCWeV4jOK0mSIriGcR1NBmwlFOgGdAGFv6gE
Y/7CDAzdILry53vkIYkvU/DjaxnI3sX0YxeB18mKHwXquwvqLee4Nq4h3gI4Dymo
T6Sko/TyWkHsBWdPAusDPuwCnryBUU1DfpEkgqJhPhlG2sSTCxsMPKqNBWq6lCdS
Dm6itaucWO9mwJf181o6rIRjDSnFuEe/qwTNBxJ1KNEqPV5l4vZJdV+LuFfzMaAr
OPJXdaukZ7DjWbj/mrXdckPDFFNBEeGY9bkOyCWYOZDzawBmZfgCrs2S5+aTEkw4
UDBd/BufWHZ+5yMiKsViEf+v4BNYvrIgIiY11xB9b4HGwHRG1hkmewUa2uMtfVT8
RON6DmbO05Xib99evMIIezdgqq3r1SmaOatD/NCZIqUNoYrdR5lF1BH8+58wG155
rrfyimQve7aIFbTH+Ecy9mrVjTiBy5I01UopqZYu98bDi8ajRXfqrtY26DFewF9v
deG06CW3KK0HTDSm7jl88wVghMKP7ARQUCi6d42jOBP+8mnWFUwSL6Mg2h56FR2Y
5cum9xPjJrpqX5Lga2s6bibNb3fzpbcct+jCl+dIvxu4mHtTcqwSdhD3/Hx3iA4T
9Sft3vV1fv3rWH+h4Z9GpYmG166ArNJgD6/OiAfy1NYsatZdJBKuzlQKwAg8UHXG
fnP70enPpyauWD+R5ACPmuKaml7G40O/t7cPbb5h7TlbOzTu6K5dmX+E0kWlkahr
IL3WbwVQsJvA2iHvef61QLDRxwnBn3Gh7Ie3pk5rQZjX8BuHHWOSt9q4Xe3vEpLa
aXppHRIP6pcbsXf7a8UIf9hDbSFO3UFq+RtSQ5MDIcf3cG1Cf+/6i3FUm/ti1x46
e2XIMJB0v/ViIASuHDk013hnk5Yn2SnWX1DyRA9j3+VzUZZlasTXFoNTA7xbwcVi
W6qFYojDw7nh+vibCUIMR/+xuCWRDe/GHvs/uDy9PLoKho0MIlexjNnHR8U8ScIW
WWJD8hZFO9nFZEdhP2UhoIhmq5ewZv1BaMeynlNqxz/CovGRrNQTBB1mJgwReIjH
igwH5kBKlHeLLvNix/Nc8sIGKiADAdxB0oToSo/z1t0ajK9Emji7oGDlhz+oRgVW
BKhPhplkEa/y8wy6cBgZwdpQ+qOeAlhi2hTeYIsxcNOPAlp7mv/vqHlgzwb7j2Zo
EXxPI2++xbDkozTOWNNuevyiGtBR5aCb6xb5Go/PzGUzpw4eZZ3FOH0C40BPKvg8
PtYOJgZBMoI2grLyaefTR5vn80Wi7FS2j5OkyNWkYEUJa91YmDErxgQBhXEQCJ/J
RIotNz0PHASwtQh+dlMYfWHtLj9SFiyW4WDOR9ED9U3cEH6geNGIhBSjU/9Kea0j
dpCbKVTa8VJfvSIkRWj/TzG5ON+V6AgluGCLaHI/XvKKJiQt5KXzwhINnBQ9bOpj
1cc+oRyPeVmWI7KjT4gCHsl9Kb0L3izalCg9FJyDL+D2IBG/VaZVvnZ9sU3e+bsk
wQqk2wh5nMLKKtdlVN5+9LLVfHYvHzFbS47RggzqJHmC1tNJpWOTs01kUiHa/Vx4
SQuDPh7/Kzkn7hY1/6CbvsNRT1sW+eDAQM/Q4gm0eZgQJe/eP2dUKaLaXXtVktMq
VRlLF+CC/UkqVly17JFF7cvog9sTVrQsA7R3G0L92vBpj6M+F3QxZedjpflnvCtJ
4Sz+20qL1lKiZj8GYzKc71lDRVuQvYaL5FP098Oxo5FpWsSdd+FxeymANeto4kSI
lfTgjb0R4EU1oQF1QTCQMAcXnmNCIfn/1LWXAg3W0lx4X1Fhblqo6ELYk2rDxNnK
Yq+DHPv8xWfbsQX9h/HwsK5n4K5olopJnN9K66GRlWDNQpPf8vWww2Ov1o7t63bF
PQL4n9dN0zmuWIQ4pwdrCJCWvMoCRk2d01FrtKaReurXrxkVfZ27zC8QearVFDhf
thOjj2A9MFRVO1GcGsaHxjr1D8egRxZF302+W5QrUR2UVnEn0y4y+WPVEprrgGNI
xpWSCrazP6+jLvFt8+Ghxv0y9/FjdN1EHb4QetmJ8kGp+xXisWsdGow7YLkxEBOY
/5EK13L8rAuaVYdMA5Rp5uIgxy9ah+dQJLyhQcHOgIAd9tp3KlKPy96O795V8mOB
2cAdOzKIXKJdBH2U6UNwyrQ/s6RQ4mI+n/s2UzQ5O+OY1zbNR1CaGtNUncKCzr1g
mn15T1Idozwd66OpPenywMrdkHXjKyCFVutgem735vkSWPm+ZJKYcxwze8Zv4uF4
1Ay5RjMynvds3Pk4EOGtb+3EqULs8IJjpOzFzUH5UODA+8AeG+kP7tvdzXpyhJNn
XKGcTpyYYJHcAxLKWBDqXMhPhz99PPqX7yIhVSvq1OJAgX4YmR7YpN9qedcGfH1p
NlNrOt+FAHj1k1V8xTWXo94ZmCzEGVAZAlIpPAdPIckH5IuypBISGJ3ItdsGUF92
ZI0EAFZ70tUtdmwwVZIbBNuZxKl0HKY8NAZcz0h1tzv0JQHpQ+wLg0giuaQZOcJo
I6MMfUU+v54DBeGjKLkbd1ZQhyAJAKEqbVG8w6gTm0kKufJQD2fjguATvWgqEULC
q1lA9eBLdNM3l0iLkaKllgK51nLyB7MlZC6BvJ9q2MzpbxdejrcyEc+o7zdLVcf8
bFgZsLyqW4ledhF89mLDc8ncSSvF/3J20geBa16so9eXbP9K5QVpT9BbNLGmtdYk
IUv8K4aJhn8vt81Nqs5rC2g42nru/nFM11HZKa82xIVV+TU08Am3eNz9OaHNwmAr
sKoHH2dacu67Bhnmu8LLkXeqKt9OeCC2jVId//nOT8iHZQyJbHYayk1I1tawP6Z8
EpDTZUe5O2yWVjle4eISUiquLxPDIQaAKuGihZcuzTjk1MV3kPe0j5iGl/rGHbSV
Gv/oPMlbgO/YZk9Hkc0BonIjLsiDh1K+JiNj7ldApAR61aKHS9cJfaLFy5xNsi8b
zGj7xnWdEHWOkW4BBU/4AaiO8MryXqwIgwGvgotuLAyAlv8M4dwI3hWspnUs/0iX
M/eiooHDdv5kNoRUHIUiNUgbwHI0jpYwPLcMzT1qJtJq7h0cDniHQa6Mu5FyNGNc
FYRLq2I0O5Lo7YeyymiavtoZWPIcR8ikMhNeDq0IlifZgI0oy2mkpNDmZ0q4mEHf
nO1f5YmbE7zTwn8o3+X8Y8Kbgb94wehTzPpDTx7vmhhrYrVL0rmQCAcxW2ce6lyr
jbAC88S2Oodx6jwlCpORgXAjj6tI+Rg2kDj87hEVxMWGiN6f0mP2U3900/Mh7I35
3irl153aYGysENBgogy8Y4wMh5/DV3a/HMygFmCmpRyKlXkRyrAle0EfkMzYF5ZB
u/VFInTgy6cVvWuSwwGmBf+SEThsdQQFiVkyfrnfAPw2YOMkBWNIkl/LCp9dLY5l
MZ9mUiDdw4RuJk4jYnuGasaYQ3fMSnIumD03YGuuUT93rh2S3pYjw+Tt1SnXDnpd
11KKdKbl3Y3NTypmcMzIN1ZvuyKaBzWOR/NM2xSnln25a4U93hMVTs7alv+do7lG
GLeNkSyvK+eQAiWKcyHtyi3C5bp+F4DtzsiCkOEqHqqeNv8vSwgdx8uncy9Evyjs
YcvH53tLwIAY5VcreKqehfVxuAp9gy3jIsdZX0ksAzlqW7kGqiOLM6BRQDxc//GZ
aWTELjg4B6NuQ8TUZA4FbPVBxKy8/QQykatLf5PCqCAET62n2GCFpcX5HE7EWfwV
xjM00lbgAUGm/Aj9NbVjGQcG3WAtPd0FiMhO28ci+dbV7sHM+Ju0DnEEOra3ijou
rVrw4SZ7TXCw25MFQpTEFMfEvCartjn/n0haWlwfCXnrI94hcrsSubZtlBlPuTja
br7DUgb8B1CKMjN4r/4bsmy8PTEu/0B/uhhgoxPKb5NSXU02s0IB40DKWM0CuUjA
784DesOjG5o8zXSw4JppwjqUC8cHvgd+92AuTkR54cTShwoWTpddPnt6okd6Qq/9
kpFN+ifY+M0NHDpDZJLQUr8BF5rhfQBZpQOlfBrK+nLhBD+Y8LyOstLDaMUCJqM2
Zko4jXZBI4NPvFVp88y7Mes2bVZ0tC4W4t6DqMCTnnsEgpad0SN4BuldF3XDfnY0
wNHP09egTyIIPAvAC1yAFi9RW/vZJSfhyDS58DNTieultG8WP3HOlAlC5ps8dst8
uqqKGEyd9K7MbLsIJRYZ0KqQFuw4ZPBbdut+BrmzlPFbx4/Y2azHuUh6vuz0oq1B
zBDgoPm64SGz1dOV7PES/7zVK9gaSvY9Rclcwkbmm2hGk5pJSgW9VJhvQO3m9cOj
qWGYnT2LmFSJE3YdpAoCX5DLPPXyc0jarOl/TohjImMRHMtpNZ5cWA29/KVn86pG
NtqsdR2p9poyjIfnnLh+59bVYZCIYzOPEm2CmC0/PI5JtBDT3mZYimpw/hlLku0z
egfQfcQn0RXF6zSICkg50pMnRLLXzn030jDXM/DtlhU/5w/qAjecsrjFaBQRJ6Lx
P2tA8iDJstUZsH/9cquSmkuwWLvsMBf7frVoQG5zLbj3hOu0Z62BnIaEOo9GXpVq
5Hpzn7zCu/WaInYE+siKy79HUFIytLPtPkNnz5ChhbLT/9Fa/T6fqDgHAgBr7GC7
UDwDnj2aXm03hK21N4vLtaT56pFmxe8YifQeJEXF+m+xec1Q7sf398g1egYYk2ZB
cK0TETqFACm26O2hP04gNptev29cfxpWhsxxgV9hR7VShIUPxksSg5UYQTIDtXHb
3OfWoAxkpLN9CJHQdZbnPCzUqp5O8LK0uPRSWssJ3oRtSTKFXYLN5iHLlFf7zLU5
21l640/Awly2Pd9jzpMGACZIQv7J6YNaCkyYLNC/I6F3DaxEYvkEfc5Q/A+4NeZL
2O40sKWNkzv93jMx+sCc96y2GPILfroxb6vIdrvWwdNOkOHI1l+F6mqK2tChVopo
g0vMwPBvaCWI8h28Bkecw3OgU7rAhGjNNCL+Eke/k2/M3z0FX1yGFKR2mxNvy585
TWT1FcFP/G3luDovaucPe2Smrj2tY5TeHOWIl+Wd/+JwXpDv1Zmg7XSV4SsxJp16
gvSPsAFJgBUkSu13gp0+k9Lt4sLlITC5oxszljtme4QtPz/Gm6MZpyTyvQH+yTIr
7CkW+gp8spZxR6POqUAKcBjRlbAOFMUqKfEfJ7164HFh4AVtDhlT/bZ+p4br4GaO
ao4kLeGypYMVl+gZKKo/uAqhWyCibOhxigWRPbnzhvWEBAOS3+48aPtKjrtwr0WM
ZsH2in/Rle+pTcQCNu7RYOxdrpVdJvj6oOLGY+a5MQijoHb1IJbMZtpfo5q2z5gw
fGPF89UZbv0Ad1HDk/15zGWbtTA7FnFUTc0HJbU5c/BHoVMeLBBvGMgUf42NNPc7
kSHk2iTLWs9ItxL33CyA8soGySuX7KhZ/kY1LGWMyITI3Az/kzNY+IHzgxjGlaXq
wa/dVk96/ICzFr+4f+Re011vUStkm9fKMmOGRRqwEw51avTi7RUMt8MSao8iYvhh
sAg9s5r22OxPa9NdiQXbFyIyV8UAOQYYRCro7s3j4cAHKARThTtbjNeKbKLGYTt9
GMIdtJR0lHhS5kmLNx48f5Bt8CCVUtfp+oWo8wwhXxMomuCXFPldPpAYt0ER96jP
+s9+oir7mz5EXjr/bCS+LkfLCn2FGXa0L/PQtoKF71xDSC9HfxGjlsAo0uCDHFHZ
ObtOlZWKIXj4wHGOX6IQLLQgC0p4b8BytZlHv+M6yYzIVxwi8bT7EfZJNtRjrJCe
M5EfWgGNxYGM5JMj15arPNLxcLvSgL08LzcaIAXwY6NE/RFdQfHawje3E+egY9sG
47FMjUJvJMVwFtQcQcHOj+GhZK/LQj6NSPqbI/eeDu1kZL2212BglcimCvoaEPsA
pxAem88m1vx5wMkNB+pCdEp5U2Dlaw5pbrw9oUwn7qkh30dW1kmIiZQhGPwQlEIh
Y1nBh4vGH2AbttwJf3OH/ZWwjqfCPhf7PpgJePZp2s28bc6q47HumduBxRXEtneL
Jv9a7s+SZ7B/uA+Aj2KBd972vtBQO8wHo5jhkXQWPYVbA5mM/CBKYZUxr2Px7EIw
d2hSQqf34AS4g3AMcCTjwOQaTn6OX2oZFsINsKhub8H0qa0y1161zBto5VChEnCR
qhP3wdcBYgxvUQWdbwA3R/WhUottddc8O8dSFitgB883Zw0eVkIhcxWwseBk+FcZ
sw8PIg0XlbK+I3E6KUZI/VvCq7ZjP/Ng/SF7hFapVRvb7A5aFa9FiLtrCurbyrBQ
TgZkOppAqCUiEbFR9k3ScF2kDXxHYrrOt0qZopv22xdFVxVCK55bZif3yIhmVrKB
elFmQSJ0whaH8X/z0IUrays6feiFYf/PGfnJITFoHPKzfpOrOjC7hWOdlTBa2eI9
K2NHyC/4g3/YliIfBOBWulXpt/giMTJ7ki4gYpKkHZIoilgWhf9vqGr8t+7/CKe4
BFZzt9XMDCXzTgs7qgASqDfSXy4jFpUo2DyVF+eqIzrwqGgWUwbcFpm+cLr0+EcL
zA6mUym7ai0C7hTIEA3JnQIFHrdSmXvtq9KLlE0SQ7z5DWYLt5Cm/Whi+z/lSUFb
XXsMYY4lFe7DMpEvzlabZUzy76CL6OpkxVE6GMv9sFCG3qvK4px+pvC3rNs4OStp
YujCFywMn3r455+k+mCmt/zLX14WRRhcDZWaumvVaDzSegTfKc0N10IuRAYoVxLd
xs9/ZCs0QDC4TZl+OWjqEuMMbeYLdrzdtProhf0Epsoovx+NwL1vBTJs6/voakcR
kntpz4mcbNn3ET1unbRX8UzVTlpAyPlHvpfdqS/VoYR9SRqvn2Iyre/oCNnlpR9W
VgvXsEG3mxpa5Ioxh3pf26Vgur3WRDeWguXDYNAGiTHJrjYiY+ihvaN5f2IA8T7m
PA4A8nitIn8Hf+mPqp3QIYrtzO9rRXcWARMEbL5183EDxIq/Iqy4NWhswTMPCVsa
AZBvQKKzONP7VeAeHxprkp7MJQQiB3owXMvDixKyyq4gxS87I1xsPRHTo0rHdeYY
8r06GHLejxpBnuPiB4leT9CT68jepA8TW2umzlvN19PDHDsMq65PIOmT64FOnlSl
7u2EQirQEExY1RWbbYf8pDYaafG4Qy/+tCU7Mh85qyf4cdzPiSjZqf49ihaWI+/U
2Ak7jPrjBqpTPefIWV2r7t22oed1tK567hh5IQBMCfvcTE03sReHhXbxyAWDXkff
5mfv6pzS3U7Qs4Sks+DsK1r4+YU/UqRrqPENgewyMClBXkR87YoozUbo1uxHbS4g
CSD8q1hAN7yh1DDLzgzuiwtEvfRQb8V6d5np/0T+apJZhOaP8xIgRPOxw3XwUOW9
0l/4W/6iExUfG+5hmCtgvtrmHGAtQ06q47eidpaiJFqLOJNs/1lyvjOfX7DX+jDO
xbS+VxAG+gzcEUwsYAI3apeQgjhAwioZY7gHPyqg4XTcnO2pi7OuH2wmfc4SB1Bk
uvDsYIfbMTI1I6N8xccNSWchCSojvXW96wbIGDHButQl0DT77LUQxVwpR8xQvoiN
injo1dHz/qk2sTnqz8TsDS833TxJL5NcJ25P1zJXES8tdefG5Y9ZSq1CWLP261nv
3VqEyutUtSBiJFnY+dToN9ymyMPsRXqSzO01o3Y1818XSSKXlU8supgb16crdRhx
wvm7HgHZ1fLAg+XuKxWchMAhzXH5JWqs/VUxwSmbs0eg/ZqsKFVBZw03uzSjGPDl
Ou4+8nrk/SlWWJwIQE5WPNz44swqhLbj6vUHy4RAZNvCPPw4OmV3htnDJXx/GsmM
++AzBi7jJtH3+rcfAKe5EJyn5I7jLSAaYitwoHOrrwP/vVHeaJ5C/xGBtqAttYQv
rOf+SyiYlARqPckBUsESfPwVEMwwBB/7iKFpp6CIKlISMcpoj1vBMlda6NIvCCuq
mdhkFRAFTKiLyEBxHbL0ks+k3co+vcsZDxx2+jpiDG2YhdKt9hD13qPxB/tPaGur
/8MsdqGhbbSBfuNsF6LIam4rDpMp0clz8T8NtdjfR/M3x9xTY9y5HAv8Wnn1x0oi
WBJUZghyY3k6xq2OICBxiWS4zzvRnGf3YKh+lFeb3dee8S+7w4Xixe4ATcGVx5xt
1/0KKIEIzYR+XHaZ70QUpALlwPSjKM0RM6P1ctjezbiL3GwLcYu41Fq+6lES5sHF
CSbpNsTXJDFjILhXorIt30tnHMdSXgxc3EW18zce3foPeZV071dWYtAeXutK6chS
6+OEzmYBIpXbCMl1nSd7mgrbTzFIAAKpRTobcDT0MTnoCPz0AcVVf3kMU/S7ncf2
TF/lWPog71EhtO0QF5lk5Jn0FOCRSzXLZoBRpmkEGUHbRG7EH7Pv6I7CuFjxAUar
oL4+QcNZoEdon1v+xKctG2dUsCExdN6FLAaSwmhNmBomrwfZpRcqAXeBwRm9BgFl
lavSfypTUcKRJbuqRBsqNp4cuWsZUfRhgToNZXivF5YIL21gbU3+qB7h1lie0E8T
Hm5gKgr5dSU3//AxLSlir1BOBgX7P2oWFh7sUBGnlmOYHSjdhUhP0f0KJ4FO2Vfg
jzlD+GcSiK5a2LQ2jvQH854CQWly8tCFeseTx/tDEjKbw2vXbWwRyJeTBaEtBAM8
ghdeDraPtfCJjkpg32y48wFu6Am7qVIF1EWCIvVq1GvwmD8pYpHW3G+6tvsrR4PW
+QpqMT0JSQyvyp8I3FC8wZ5lug344zuHKQ8z5qfpO/+f7tQk28wFCpD4jE0piSxI
mk+hHvZlUgmfsyakpNoNwvOBHpdxwrTqyHq6dpbQb4cnNyEuLvb7snFu4+P+hLrJ
uivQZU8jecI1kEmgFL/55M4ojJuQF78AhuAsmzlCrZqyXv+gbEIq4o52Zjr3boN4
Wm/7Mm2Y3GDev6c8uykah/XZbq9Sp9bjgsin9DDtP8nX6VlwPuxOBfwfsLrT5XGB
g3lgz1zZBFfyok+TS+NF87Y780Y6grmnUqnF+LG7/FQDyxA0ldq96fd5VIHIgV45
4Q8otf5JhEqi8cFffZcZcULMDMTUq67I7adYwd2pWONgRAO2aZ28Lusk6soJvbKE
JQ4S2vmfQOx9VtUoCVLyKlmluWZPoXd8g38M+qflDHvVgYKYQ47K0HgObJtdobXO
ID4O2u+nqsYrusxUblqqv/FhM6qa6CPkISJ3GV401X1xi0Xfx2j9OsfM5hOI3Xdy
aX+b0UxT0POoPVclBK/2gaFrmPSDyvTZ7xU3Mbi/juIR6MTxiZf1kCj4kWTVcRth
8EyJa9pBpi3tjuAxVQgAyJuhdEg8LjsMWwmuIoIPuw9j3CiwZVngt9HVj0yhj4sr
IDVOgT47S7LQMGwmAtsQ+EjmxtOfxk5qkzOneWAOqUzc//I7b/ShRV1nT20nfXPy
rIEan9dOwUm/x0odQhVmrzUURzvgXdLFKGXrbSO+46NnY4jaahuE3f/U16SjbH5u
Ypg4e3fDwN9sksSxZHtIvA7+Vz8XRkM+LBUTAL9ahUBNJJ+PjcXzowgA1wHAskCJ
xm4ed8NCPoZCsTvc/iTKzNOJv0DMLLoP1FDmQuIMB0F07BQu7oR02DVyiE6JQdgh
UgIEqk9Hexd2IwoBq9WP9TEuX5kmSFUgL9REV4AcvWV/8/76xRiAeOpQyWJUgTJi
8HvoNwVRts+JhZ+/mZgNjca5crkadlxkzmPwbCA1ULkigrRi2i2PKOs6emddflGh
Aupq4hfyBXiGLe0L9mxVaqFZnScCi9iGaDUmjdrkUZvvMx5NZKUSNMVIkEzY0Rmg
jvwpMzz0Agekw8HaVaDAvpPqvUqCjBhqzaXw441ig2MPGTEESTxNIC+nH6QmHzfc
LPNuYntE24QPThcJVSEfVsk19MVClJxn3sTxfsmWdOiDgu25spfOraaXmNMiRAJX
JtxYPpQjyEmmqV7AbMS7FREqxpvz6nea0N6CqfpWs4ACxYM4Wy5ux1qj56zYAQqT
oqPLHcjLRf8zRQuscbe9MPcMxPQZ2xqsJG/S7OC22p02hqyPU+3N35YT+ShldOtx
9sICRAf8aqr4ZlXRA3uEDgrzFkCL6DMf+9X6vhzW2YzR9WdDCIQkSDb4dHUx94tT
jzOVEJ9leFsuv2mwF786zdEZBh7H62xFhaORouFTLZz3nSxQg60TxgncdXP19WRO
eFaty/55TvGbUEMGX7UepT1anJx5C43orwZ/t2Fyh7LzDMA1K3lcOk2bz1ffCWPU
Ts666w+bFZAMOH1oHMhrr09UF1xtKKdM1spU/VHBd7I5QlD56UBcVgf13YK3SdD8
pqbv2uEH8MDCiLAf0RBX0Cxh8CDj69nCd4IxGqjsoPg5JwT+PbcfQThGJ3DAXJm6
uLTAZtFXDdhzktIwm6tYalyH+75IbQU73h464aGEMrS0sEcXcAJbywYJkV7ETS2L
iH1WtwaD8Hy7vp0um3ln9vvy8LszCKSEzvOwzanhKb30P1wsQql/8dsKhqM27ZzV
lWfxRVXr+rOqJsrCEOb7wVqenTv+3osRLhhPVE/FkDnVQIwqoIdFHrFi6y7At6vC
a6fSLso0Gfen0qk65Ufv1QNORqmUxtL1RG77Cl0SG3CXzKhuftRdt5UYBTj/7zM2
VqdnWhzHIlAxI4m4xiRQPBmFt9ceqRQdVEBL9w9Rsm4ecR4ULRh8Y2IJSUnp4KV9
3uRiI2Aj1rc6rzQIsKs9aYD5osKEw9ksttBf5A144xHJCGzdlL7kCkjq/OuiTmVE
OLWZ9sT9qB0aPcjoIxACRVoXEElMtJB+jbNIH66q90P3SYskJQwL2hXnITmHdGMo
ywle42LgwVjnUM1rnS9JRcTEc6usDxu2n66D7zsCDMBL5jpwWu3mKsYHShiFgPfB
JpUOfRV+mnAL98xRrvNvWrfcJMAxKrJRJ/cmg8Zd+70qZvXLzRjQLrTlIOKYB316
gCIdAOWJezDpogv9hyvJfipvCQ6Ijkq+75WoCNJeD4FAeBcTsMzHNRVN1Mh+JSQu
xLiZCrl9shLg7tQjXw7HwCJpbCqJOSqJPuYtg/zwjX3K9BsVUN+rXVTrPTLylrqH
GNvtLN7RPOY2PRc0sEBEp9BFRlf4MOxCL1VH07KKcMnWiQdVR3vGSSwwTnEZcPEO
tQqP1QiQXKmB53FzcS/6XVsjfCW0xWvg03qrLFnOqFuSQs6NDoOaZivnFbL0ZG4Y
8CI09uimG6DnU8Fzt2mymAWXEdSh3TnBBOazUFWqEYye3o3ykGD0AswlP4HbKTa+
T5WZ0m0T7d0tsXvsSB0jHZYnM9HHGyTxpc45gsQdUNqTrP2L89vJrrlgYjTy+stU
hJKVhF3lr2ursaew0ybSDHh9l6gHEJTb1x6KETUt+dPiiGwbMGFOk7nSQXh0nyqI
gY8OgNPyGSZ37+ff39xM1EhTJ9Wij2aX2lAAUftScvaZXff+k9h2uwdcww6xPn1K
W4ija4zwbTaLanASucC4NIIBQ0YYaje03rXRhOadz6ltAcPOnfQtciJB7DAYw+bO
3wCb1qqTKbM0/dN3GgDplI0drsfZZEj5elRfvCEPu/ntf9mjJJuZUsxyqeJKt2Hl
U+HAbxvVObbjd/8m+BPMs/DIgGrODTlutsicsdA7/HZl5qCxWr4ejCpba/3P5juO
hTP4rp0jQUDZ8Ht5jHpeRRtMVB6l0skMl7oe+tvN1W9Up9crKF0N0UCK0i18w8k5
Hzg+aOR7fReWxRFx0xb15J8dbO0qh48x8cn8l6KgCgjEh0UdPPL1VpAUM53xnJ+o
2BwULoeF+Fvj4bSqTqaTi78ILb3Buzm7VnNVw7N9p3+kxKnp8R8XE3XmebNOEKMh
BdwnClj4s9bPtM6xnwP4eVjm02iS6hHxo7lGZ/48gQtke7Dd74qJTD/18xTmj+sU
K+x28Evrzauc4TbGSEH0PQ+xSi5bx8Ox/dQTCAz7V4a5ePSSNQclvXhcWXsn1UUC
QjC+k7AJVZN8H9TnsInU/aVrkwjuRdTmwYnwd3kDl9TKRJIJMp6RHkQNC7STHYHu
G+3mfrda2kaPBgkaBcei3gVydaLX9qUshXq27ZbAnJJsgtZT4JZ7K4V37pRpxThV
ofaeoRcRzk7OGHFy7t20F4gQoBJMEJl1ZLhnDCIzqv2nYbIjSrwt0DQ8poa7GL3N
jl+4v4Wtw7Hyohi5x15wGCnnEgUJfCvsathnzmw5PlfLXWWZdIqVGzzzSEOe4qYO
N4vuJBNkgqLaeYfdwp5n2xCXDLhMpNDrEH+ibrN9/LrUEkmRB8kBVX6sF1d0uHLe
JYmXikscwXxEpYhfXIpQjaCH2MaguORGraSaJk5debXrzq46o1iaTi385c/iEFm1
DFIU810zsCXF1hI1Dlkkf/cTO1WjRdio37tMb880jZPSujf/miNDbxcQ1gAatCGK
CIJf6c9yOvKtl1o1dKG59R1cM4AIXMew7TdziuhY8YCpkBHqNVf3vXSN6qjH0qNt
+Hzfm2y75fSfWWuQ1Z4GCtVufhIR+XWnTKuy0zJgL/qGfOOyUfmqUIelCIYYwd0g
zRhLKnHHHk4t8mmsnJol7aPP7xBNOhjHNOorJdtYCnJkojDYKHgb3SY99Hw22Esg
125oqb7DjuxuQGbS+yKojP2n6dLWF5N2FmfmwypClIN3HM3xQnfS4HDAvDxxw5cS
ZcR4vaqnpMMsmaBdlbn7TUWV4xxfFlxwiyA25RweaNl7ybR0CQChI/R3MNgHWA9H
r6M4ImhUTcz61zvwy+kUofmAGvFHPStEbl6saYUyRI2FUwccRTVPdlUQTncVXOEH
NJrPNX6srkNJigZienmh5Uy5DwcxZqIOSvwvDxKuZKqjKsT5+tKdSWQKpIFbgN5g
MExiUz0/tNoy2D3UMOBSESDf4sZBytiU/PoFJqdNn4mqcVeqIX9F9AGBb1cmc9p8
6FQIcVqxE3NBHss+/WRA7Y1FH40ptFuCPTiWc9zyriXW958RtCXXZozGCZOLcyzv
MRuD+NfOWQIRCpQVkyW3t7qSn1PdUdqqMLmAHbbK/EGYapX7xqan2rhbFB6CSV4i
vyi2uS3QOm+gnsn87dUZq0DdM1KrtTO+U6HNW2bpk1t+YnA2eFRnAUqN+enV4srx
cL7b6TXelI+riYCDzUPu5CsFCFcGn1oJBU1PzaESLZsbes0St8caELvPnFZdtERA
/tMoT4G/ur2sBv/nXYJM3t6XabkcDJYTXu2jEvqs6o8+Lgm0Crefb6YHtuz6aX9Q
QVqhcqaiPvYzartkMhJoBaLW2Hie7U0MEZekAU0PKWSfodA3AXRy6dI3IRbQoHrD
cCvPX/3Gnf51L/GNNkmStLOlZNbw5fRWBJ9wNt8cXj6v4Fhp12D+O0dpXbKXdt3k
zUqtg3JX3iUamsd//2tXWV2dtAKmnc+uxKFgxFbwa0xqppE8lrJkYViTYlQOHeoh
ogDSN6Y/ierQcUiGyCiQ3Xq9zEBsLHPxbbbLP8qnkWvystJOOESQh7V1dZNp5rqI
aqkauYCl/OEQsMl+xmcsB9F2m13/hirJ9GqrhRlbR8H1wsbwrw+P9WvCtCl4DrjT
cmW0NtYuSg8khSpb/OFSW3i4nVzXABwFOrB2lD9YQi1jSpsfA77ouIVDwHMUhF4G
m72eCkiWSMUNq2fqvSlL85o77B4sKTtyMxPWar9LMaV18S69YBpw7mJ/aiv/o2ta
MZyrpyMyfxkJa+GR3dd7G7t48WynqpeF4cYJ2IWuM+5Ui8/J22HaBF0pmh2Jy3Db
Hi5WcyO/3BRd5S8QKNGXp7s0N4oyT7mAu4cU0tFosD5bXXGAMi7OaV83XL+4vPc9
1h8unT985cap7xA6JfSSVNFvFKJ92f7ebQ0sum6T+jXLU0IR9c0NnY+CU3T6KwaC
RlcnQBjjo+GMyPAN2yzfhLXs2vykiQe3PgQZl57lLKrlzIdXKqxo9B8FgAyjvyjp
fQrMChN41ShpmO5wMoxqsnxxk92JmMDdo5DQZknxFp2AeBLYkUbDKYdwOgpCkwUQ
kFeErCMdSUJLFtWFanQ1Y1HZUg5n8hRPdFWhG1Dqg7oRxnCnoJpq6hGpTbF8AlTu
/0Rt7rcrTuyUX/vs50MLAqCPRZsRen9gEM2ZdpKLb8mi+Jz3SffJh8oD644nNdlI
/LYSDPicehT6tN0AWvj4+decGmfNX70zKk6oJ9l24GIeMcrPJVkFnNuQAce1bkBt
RqdFsS6Ok15hE8yQH01EaF5wICTahCN+WG6mECghuwDUN2iqceC3B2OQUm2YXLYE
JC3oM1wMpkCwyN2u814Oknleqylk9AECV/r41hwSGT6GFEXCFoT7oMwVIZaY149L
znKGeqUerw3TPK1DXiEUkTbWevL0Q1UgtBFZH71FjBiByTwfpmpjqZUYhrZRWC5i
Hry29EoHm4uvGTU8tHSvrRaTxzPpyATFC/3Llr2NL/8ahDzajPgHg4tkd5KsfU+b
rTtM2WLx6+iah714LIOSRDMftGqn396Gkwy+jK0XVk7vHCsdtILMg1Xr542Ta7Qe
VaDNmLjl/rNPR6bZ9QB2hnScBPZeRO4f85PLAAeojqWQbsib2exIYlYL0PfQK2Vi
4qOJ7louVxrHf1S/lnOIZ7lvYQ8PqmoZ+iMP+jSfvz4O0uOkVX0uJYlOaHnPdWpN
+RIRIDMQLOsWZsHidIipuqtq6RB7fES65FdTmJAqMq+J+BNRRmhf52v86/vF0FOQ
Em23VySSp4YoAlJeKAxS5nozxkeWNV68TD4+8beTgKWH2HyA8vLOAA3rWBGfMFjK
rT1qbjNv7O5kqLngyEMXy9X8EN6JJckz8Qp2mC52EWoNXkUnzAySKcFsZcVCiFaA
n/ES4cPwEgdcpONKMeKrC4xG7GGhLSvCoVaAXaZiFMwnH1891O1EtF5gzBCIhR6+
YQVUF7JXBY4DkfQx36BWnD6CWmcPdsIxDg7ggomOuXSrhjroCs9P9PU7LsqbEq/i
TxAGpNQo0MXFclDwgTt69QdE7AGTqV4tWjVPR/wYIhbozUAFkwHIODEHricGMUAb
KzQi4Ic/AHd9EpWKS+UcMilbYU9vaHshmcIxC9q7NH3bHFOmnO3zqOkXt7cmRrq7
UDr0EIn7XiU4hjk7rAWo7nvc4kYb2rm3aP+grmRYV8NI3UNvOCeVtBbNJr9F0p48
7wSbKM88h3bam6w9KtDiSou1sfZTtJe4lnsPIAUVdErhSgDabQAY8OqWNCe98S6K
TPoWEssAQ/5F/VkXA1yQl5n9jNYfmI2VDvnTjSNeN5R+hAaTXgaGkCQADQ4n62A9
ZCgTO1oQq7rxhJcdIxscUvYK4i/WUaWIWdEnAYjgYKmqRJIzjmPbWeddDLlpkq9P
xqcpt/Rfxzh0VGUBHxr53tzsK2CoqGg8Npbv9+OIhLSd0vpuPbrxKH/pCM7Bl103
p5xLmID2xDPsIIdFV2yOUELtlwKvixaRuV1IpDvrxy5I3d2Z9fhokqNCuB2NaZik
w91GWlbQO8m3NOKkIwjK61t+D6dhEVhz9OI1g/J5mCIkCpP1NJ7MpT9gHeAFhV1w
uzw06XiNJ+Sae/9NO/MZEZx6cfpLp+wYh1fIhAPL9n9GaOtT2aOtnZwHbRR2zL3Y
hArPIMTVaSNTuZUAIi3Etao7aMkC4nDJ3PE5fOwcsMDBUWjSe/ei44GRXtAZlzDy
stdDR2x0vq+hG0pQ5hxLffg6XeaqeYJZ0oCHq2dSvdG7ehtwexpidablM8hg4tJq
F8ReCWcRZoYKGwnSWBQ/YFgwj0IvHoZoZDKZ9fGA/27M+Hz6h67aijbZjgiaBUxV
3i2xXw/doKrWh0m6/A8ZWPeJ10oOZFss6NCbSOgJN5+Qqju8kdNbmOKBDv+HmTe+
7LQblomRxTb/pUgtcVy2toPUPqWPtK0PY0VPOGj4UHvriBXuIAmn0eGVSY9pAv6x
5joMAmtw4bvnJg514694wRqW9j78Et2iAoXX1LgeMF9P3uRhQtLgkrrPsUZhfJxH
1I68hslT6hFBiwH8Ls5VfXItTwUmnOXL7CmAlohgsl+A2CF6End2sgvkPL2pQ/rd
7MwTcXwsQOVOYh77Vk0Jz0cB9IZRFfYThmJs76kvDCi3nq0ulc5C6xWFW092moho
p0Y9akLKQe9R8O+KH6xiNPFTX6q233vK0+/erLtsxMtwjlogp+1ClY9yWjAbMXFv
WRXJ7Sd217Elnx+O5J6Sr+GhH2HyoXCPVMBzhXrXpsKKxr61OJMlSuLQ56s9yEjJ
E0Z8ipju58BKrqyIU0j6zp/CTzpO7hlPWe7nktWv3Jufe+kjFZ8EZmhYqqvIlI7a
1AMzxz+sGyIavAA5Kqh/aTQaCcp+u6gJvKjr9cWpyXQrKu4NwiiX/f8u1TpCjkpv
67297YZ75Jcv3VaF+5bGPTRcWxBiewXMRLjo6Lns6v7xGAzI1CoGQ4Mgj1ftOEkv
f7SlVS1ecCfehpZmoe5+2+8FJKtQLo76IIGJkcBYuJH90/9VwtfJRjnhpo7GdeYW
NX1NZ6tmsiyt7xhSWJGQTIoXIOC88xSTYLD5kqhX3yOrLY/aiWyKwUVSSDnd7qOJ
Hf8BlgMCB8IsX0I04XPbAAMl6pSGpqykiQo31GzxTLtmG7LeKJ9w5Ga/pn8JSARS
Rhc3FJNzICimS/DM0z90b7taPMF016tG+ruS7IG8Ta4akOmohRP37Dy8tNbgjQ6x
pWHE98ee4HhLtUJM0xEcHJAzEJtk4C292v47+hCViDdKrgC56w2wTy8Cb9Fniq23
sTXNq2glutS8HV0EVuAMEsLwQbWAxp82A+/URkQdgG35ZpE8aNcz98wHTX7tMwaw
OB0qtSF9lZVZiu96L+h1v9WYFbykmRlbPEZA3mE41QbN397vaNrM8/jdeCotEk0G
ikdpeTVc1GvGvmkSXOX9NjLnQyXwJWUQA+GP1TaKLZnVwwf3b4dD8loN+cgjb+KE
oSQUOnTR/6qnRZnAZjAuF77jQ1B5zpjEIN/aobxksFxer9jvn7gRQb7bM550EApi
hWg3eQmNU3TVcaGOWL38G/0C6P5JLEKw/WzdBBXKsEJYBnWhsRpyfCL6ZfRLESq8
gCcWCiLBYkiLT/PTlB4Z1c9IMc/EJZdOPKex1gk4ZyXIfTAc6qtcmrAyLaVvm8bg
VWe4hQqpWTsJLH2n1+BeGXEyCTBg0MglIlYQiXTWVgpT9x7OJUZyp5hbOIAolSeG
5UlhIjWye/K798UtahqRA2/vhuEKj32a5OYfChpzNNXAaU3dN7+ZkYK+F08Wyg40
fjNYgoJWl8NYwnYNUGj3OvPK0mfUHDUclWOKiHymOeiPVfyJkh83G2S8AEx0qxJK
GeSq9NU2l6jY0SEdyL/XomJTSqCaHSzUdnXt7oL3qqv1QjVG4Iv9o6xoyOI/bFLE
4LgheMW+adFkzS1Cg3j9D5awGU5PIE6Sp1v1WI5PqFcuHz9P71ZyoXRZ85eMzDum
MIiyR3tMlYYqSsWtWG39DHIkZuMXHvR9sl1t32IrGCBk3/ZZgsW68Bkd4wswAmux
svQqF93+6j4sFG94sdVpkEjH04Ka0RWkKGaVkBtHYnNfgzZtbyjtf9VRM1mLydBB
CAQJaWQyE9uN9qMaLkrcWiB+V06iI4zOfZ/zi9it0E7fl17wLXlcV6Axdds7D/AM
PZGO/nIKbi685M5JeQEmymTeN3ld1Z2bFQEq4F6uCArfo3vR0+ETON+7x5iyNUER
0hJF1IlpfU/NSYnBKDEMogp/0xcce4jnkgFxjKA2ZLvqqxAQAy/5jbOvunIMdNE6
zi4JGo7GTdfkpTb5+5ZlawFPlpIr5SRdvyNDlvWSnzPBCK4uBtIeshkXIr80evwP
SkGZMjWjGcsueIp+gEi55UTGrT6TzRIS3Iv+guvxaD9KKcKB7pUJnQOJiUSF8NN2
XZSu0rzuR6f48u8MGMm13vud5aLyuM05giBYGASX1gHXv7db6Sbl+4IjCfMrptjG
0aP94agED+izlh5k5mTEIL60UC36O19gC3fke4KLHHY7DcWtLt0efMGzPIbY85R1
qqefRkJcVQGw+sDk6h8CCLVhbmZHKwDuHAjrgbObqhqs5IkXBImb4M1CXUDel3st
IBl7c5nT2CtfXahVNq1nGhQGnIxeWuD9K/ZR8oCI+zBrVVHgH55sk0LmowU5DfGu
T9opp1iTLfSawdTogsEORDOgZNkseBQtAUAiWogFQnt/9yz7r+57Twmeuxh5e3aV
cT+h2bn/R6PSbE8Xh+cKRqebe8Mv4iZnCIrRloAQwLi965jTP9Mp3GqpxEfQgnlT
jdRjJSUatz2lRxptaiP3qU6FnQwyhq262wbmCF68tCLuSeHkBlDJ96vMDp7d+pKn
M9SX69IyIy0Q7kPlLxpFi5fwDP+k+5u+nAUrDekxDbUH29m4rDDDNGkoRtOS4073
qioHv7gDy7WHoICP+7v+/prLvoS/ehnj5GkXudy5zyMkemSo6s1XUg8zlVBfjUUH
VYGAZmVvcA2D3fX8sfiKunrUsFGbG0x/JjmotOvhiEpv4X8YTXtSQVFzmlhic0Q6
0hkKtGcGCP0MkzxBV8E3FhqdbeUPgtdeutdSNPO+STjl+LhF6Bsiv4RJjrMm0QAY
sw6btd24b9tZtIRad930VzIf/vqiDhx/tEAV+4osgvEB4WsIR+ZOcfoQdV18Jj2U
Scbo8WwYytiwdngozz5DVMA5PYQorBga2kK8COeFkuGMS9fzF860CPGeFZgTXAao
atXRveakFmAI9KRhI+F/QZIYNji/sqLkBGFZiOMEEYcBxbKzP6Ic4K73SMlKv0bZ
OaHQOJFOZbNF1cmN+75+P0nYxAJTtvPrLPEIqCyauTB/2Zu8P/3I5YNb5WuNYbgE
wKgFWzz7f2a0reTl/mygZauJnU39Gn4X+hT4jZkQD8qQj/P4+5sXHYY5smBK4/l2
AZhLLPFB9ZfVrp1L6Q9b1HCuTRd/pIbPbHe96GL8J1zfDNBcEnaawI41f7/2Mpl0
CL+Sd0ZqpAuac9zdc/Z/n6PRqyTf9dV1asq9qoDMKX+wJ0+OxW6VKSX7XlDWf+NO
QTz/92b1N3pepXPgWMCltix2WTKE+6z5paj0OAPlhDzTnQyYfzDCWQOshWnrvbL5
V+GuGfTtzN6I3xUMnbXzKknt2d65der3GqEpz5KffqwHvrpdtzD0/VShfmnIU+5v
/M6lAYHViG2wJmUEXttNpTNkgF5i0gHuQp9udS4L5iEQuhejqjA+GMucwTUHt8XH
Vnmc8h1Hev1PVnX3M8f3ldhbXD4SXXDw055fOoW/7qujGxsMJiUqqFR2sSo463/Q
mFsad5GzbNLvQdWB002JEVc3bpEhGyedzbWtEvhvOyWVlK7lxpHaZvNztEqWYFVm
CbgSBSItrSm/MReQUvWbZcfU/ImgnGdRqLl8253m2u8cF/wyHDalYKfeZNauLBye
mLD7buvmC8eJSEcVqCQkEPqPo5lguJ9SBPLdHtYjnpkTJMli9UXJd4BYGb3WWpRZ
WLBOYOhCrSWZo21lxTX4sqb3MRqCvFFpaMT6FLRTTDRk+SiFqSSNuNEkf6pk0IKI
fW5nnAwgQKUPWHYVq0Pv9ghYX2IIJ+EpxfYMVfYwEYlMrSmla09T3VH634vHa/Vw
Lsk7KiGIv1Ot+2WXVbdiaQScHMl9rnKfNnxoQzcv0nC8WYjom3W4nr43CBFfzTeo
b2LM/eacTKgJOHB62NKquJo86OasPHQ3QkH+4ndnAc0oAVo2RfilTNV2oizVxFDc
iHQDlBuDj8nMselwTmeeRbdYMeUfah/WHXiChiqbUEWlNJHl6OhN0VRW08gSQhPh
OS3veO74F3K6Ndy/HpuAJv6Tdy9vUR9TWHMrwUFuuzNGHNhi1+P1xba+awY+Vx6n
oEIuJDzigqD7XaS+UkvLE/eAGOEzH5JCKJc0sK5VSvkPW8HbaJ000/how6UdiuKD
DDS3z3kjYGSakrcGSlqteFK9Kwk6W60jbit8i3qRWX8wQTZ7MrWx67MPmNH6OxEh
b46iy4ZpHBrT5a+ClvVgpJmWtxZ9MqwjyGR4tv0poWeP6uhr4BhpO5jas+xRTz5+
ztQx5n3fmh67UdtEmy6/6gGG/Ug3E2LmS1BYqmLF/WxJ51hYY/KqrGpKHHIk8ugS
69IX7XoxZqtr1T+P7QrgLuIH8ekqjBGEBgX/59SydkAoIQ4T0yeGeDAQtXgfPZOP
0xSe/tvLUDwAeusCyI5qrdxWl0oJP+qN3ywtm1PVEJ3HqKl/Cb9LaNEBgt6p5yzX
aDEkjk000hhwtTvJA95T3jRAUJhADAz2EIq3QCwrLhK/B91JPfTWgce8/mrEnpEp
SoHIB/5mD4E+GZ+vbN1iAzFjP39MNTd7UFKfQieNnVDS1aBSvRnUVlQASJhT8hLT
DrbEno3u5keEPQ6Q3eSvc1aZy+kvjGllAST2Il+eLkfpQ2i3+2T7xOE3P915+wKw
4Ovb/Faxz6V/XyG1I9k1ks+8FPfuUm16/llJLpriOY1qkEI+owFf9kE9InVV9xwU
lDrEchzexm32IcufSorZk03vKh4jFmsM5f2zyq6IF1vCEZLsOv1n+3PZy3ZSUkeD
+KVInR/j+LaNnB7zM8dNm3AiX1E592nqSWNslF1/V7AMi+ILFDvVp+pKjEYXOuu5
e0BJmdkmHNRmB+5BQ5YHscUatM1VPdP78k1TScATgqPfP7bDsSlNsysOlhFdlfuE
TqxTuif9jvY1M0JySepdnR72lwBL2U8i+baRzhZfbywoAXqelMOq0kvd2eb4YPrK
U7DvGIRcpNCPkWhG2/BTvd7EEGrkwVd6zzQDDqLAqUyWVILLSzOk6WquDmI56jmQ
A2lWW2dcFktLVegJ97Px9zY4UuYcLxifTCaI81IAxd+cIxZTp7WuCEUFvydCF+I7
TrjtxFoXB83vKzO0CDnwvbJNts7DDv5bBiQPZPAzj8Roveu9uxCVxguGbdAU7gF/
8xffnosOZDyxTWpikNDetnQdFVnIGch9pIY+nohMHLlMPaClpijz1maaIQ2VBIuD
Bf3pXSLPbL2AjpbHnVHd6GJBL3g5LjNXQsP4C9q1r/J3LbHbojGWgSMaeqWV1zcj
AfwvIl6XD+w0Kk2XnCVwKSLSxxcYOh4Aq57dThYCLXz1MPeToouREfZpd8QaQihA
11h0KmmUxuvgFAqSfuo2u7pLbKoxvBL8tJba1E/nAZ1tN21qwvw+uH/wl4TjeOTc
P/mTJ7lgsEbHbQNOKDkgEmJ6bgPnpYhiUUSHM6F24cs0oQfuOt6bAJROXBogoum9
9PUCoTunPW31+bV9bjB/XnYUUFUgyszeHWfCFdJwGfWLfhki5AyXzh5WzuBXc2CA
cwExMNFK15jqXJqPb7zGL1ShTaXQr1mSrBiod+YEwPrscJpCBSxeyaAimq9cU4W9
V1D7cE8PbK4cClnD3PBkRQMUxodIEvc5r3DIXW19dELhgVocFEoXuJg10euFigNk
pWr147OlkzuHA3T7Y1cxCyzmCxRDQTKAsB5wf8jcyklKZYl+zwjb/OuaAiM5Z2Qc
Wprf1G7xcNPAtEL4V3sCaGyNhuY6M12Zr9ALglhpZMqcVhDK7RBdH1rQ6uaMNB4C
A05H4NvREYTtmIx2UYMEpFxh2eAZTrO+oCf8vl0L0JdG97pOWyOzfrqchPzi3ai0
hBn9qpWxdLpXzgCeXgmluFo+rv6ZFf1s05lBVeVwcs7QiFBVHAa+h8HYiG/JEySZ
vR4AKTQ2BlT8+8ozgeXC0uWCsQKIfJnOscKvwiWjD5oTl7agp+S4QS1rnFUA4cdm
KCsMLvh3bkBEFHN0KenHnf+xp3omuVd9CsARxRvEkz+BaOgjSqZuoibuTPokwuRK
X85Jrx9uwXZB8mf5v0V5aPimYn2ZW8VZXSR/qE5SrAO58XE3kJiajz1Wpew2s+nH
/5rR7NQD0SEWbCTsWrmZ01nXr+nWPxm3G4RnVTfYJZiOaLv99pafWu80K6D9I044
H/K89SapKGh4FW1xVwTToA+gz8qim3zkboPc1S8HwJTfVQh6k0+t72NEIflJjZtU
CCG4BuRRstCI+7rnLXtNldw+PSpRcz0Ls6IWbmnCr5meh1WJNTh+n/BbEUG/WJF2
X32TqJrapUpq71rlfuUzSh8zqB/nQne3ro4kXPVuYZCit3RdzP8q3omaIYwqhtgQ
m9u60lj66Un20JK/6WR1RKq/FGlSSJDdnQIrN+a7d75RRD3pAKTJTc968U6TVBCx
L4fjvbhrju+cuXzF2KQkeoiEDxfHEYS0EVEfQDAHDWXfue8dQgj1hm/mQvYYAiZk
kQJiyNm8V8sycDJn3KBIw6pjs9Dxn2vR9u+Mvi4NQS/LGNLJXE/AvK+g2oeQHszl
awyHp7lAz9rOmwmW80S1Idm5Fo8bUK3bkMMZf+qjHN0TXrFbmNjWcUHi+4KBO9qm
EqvFdrf9JEcOi75PZoEb5/aNMhFvP/Ndow+3wu9ljO46wV3vIIIAxSDNR309NBn2
IMIDevObeYEHE3sBS7BfXF9l6eUJZSecO/83oivfOsMm1g3urHAykFJbIwqsYm+X
IEBUquKjDcVKaFScW0AZwjzadkzS3RkYP9oJ9asrWn2KIY4YQJlOBRkJ4ABiOH2D
zDvJQO3mmu6FZneDKWEL4TzZVtpAEtzpxW8gUZVL6wXR0JoL64eowBhMQMAya/O0
+LvX0Cj1Hu7xhAkVqR0i7WViQXVxyLn6w3gtGzwR0txEpAWpV9AAu/IJhfv9Nbu6
vU9UguNSaJSGcD9MfNP0ZBP1xezrnFnUwPYwVL9rqhlYQRcAZYUz49ouMqVtDsp+
4s3KwtHcEOXODeyLWZhmqMX3UMYCm/vfbwLvNP4pLxEEKH44xns/kriMmk+FJJ8H
B6Reavda8r4lzLYY5AZcSLy9KihSNzMt/s3VYI6XZleppde8grRofCS7T12L4hgQ
CZ/flvPXyZM0MON2k7m3A8BiXwbAbfU9WxjYhGEkGtVcKYZdn9ruJu+7dPib2MTO
vgvMdzyJQnlsa0zQJzyzgp71qROSAx+kfIQC8CAP/PgLz1w6+xFQO4nematE4RoH
yGR0IyZZzbUdNuIGc9VCHxu7bgXVQz3RFjpBrcblD17hciOum60ZSzTZ1NhARBuQ
OsJHhZoJfGTctqxoyoCRwYPR5QLmwyaGHV6KpCB/QI6n3czDYxD7SKw72jcLcNRs
lLP+fY+Q/SbtPWOdTy2ttkVnHbzH0RI+ewJkwCOdMWajJj0TVgxEnNxy24a+tWZU
GjTCwGrMv2ET1zQUiLahZ0qGkU02naTfrXnxabghRbGmytT0gxNL+VMV9kHlsj6G
dy4khgzRizvMfNhbDLnxMAUvH5i6XKBLSUsImJajP97cZ6K/AWLy4y5L+KWFUOYd
FyHRPUN/Hq9/EQG0BHMDTkqP65CJVgsUbGulVAg2QcvCC/Ac9d3TCbP+0scvVX/4
5/Z7fVnboTWvS6eHmwcvN7Gf/NE6VjG1/Mluo8CPY8kgZc+bQmSUybiipCmuOrfK
LxvsHe69NTqUNNVLN3VR0HwcMV4JYi/Z3YDv0iDGDAOGaKe5l9R4wO3fUDy3R/J5
Pv1xmHtsRNkhGP0B2XYjWBRQgRP+wyJHuQvDJrkcpMHHC2JffBda7bFBhxqBhDvV
AUkenK/PRBzMQ3tDaBqmqUGT9PHnusMmCnoNp2hRdibhAmbnhvLFCYrH74Omat7i
jV1L9svD8NYvMXa9mNChWLGRjj61akYjtyyOzOd1yyiEaa3SxH1EouYKW5QSg9S5
wo9cOYagG4jPh0hOJxV2xp6/u2nqoWqjr5BA5MRCJPtKMBD2L3PGOeMAvhkH87PM
CgRwlf9Gppbi0iHwgBsW9OGRZeIXTL1dYe431+KDEuqq0LIKj20eXsqSFGQtcVXy
D48rVKlwDFtgQiWyhCMmjt0PbgoquQxadg5bfBwRmM3Q6C/VaTstYxrkMF5LCrJs
A602IGjbbTImYbTl8VeGeocTyb/pthSB+WWcKIK3kTTP+OddroFDxz4zlstXdqJh
YjcbK0KAP54Y7QAFbRE4ARanoqKS3tBPsZRc64wb8AgOfphfAgBhhv/IT+eSb8ie
+pOqh7ZOnUtYHRdAeMVW0kLhXVemAfH16uIIQrI7LGLW9Vdv+XL23caV43D/1eWc
35M7nGC3cAfHwxiECpL852SS02RnMRYbSTN9EZn4KQxfsllD+1BYf/y1vDNTmq8n
vgCwG1WBNW7tYe7HqUl4tshRMsb6rgJ4majWGCgei/97JpDVSy9LTSzJEqOKEtmV
pnKDz745A8Uvw+Jlz8ZiRCPPEN3qho8VtFHxMsmSGEPF/fdqqDfiNxG1wtS//t0q
PWTW5SFBIdc6KfK3NVEtM02A//e4+gepV8VwMSZH/oKEYyu+ravkTCeXVSMXCTsT
cj9MDFTsM6B+ZwCBDmmUvLOrapaMBl15EPemrr7EvIb/XGT+6D8yQadcGGknGlcn
zhUy5luYPWCGeJ5cAXML79A7B/UUJQvoPTauvllra0SwqAFZr/RE4YSwevNgIbSA
RNbjdt6zJCw61NOdEu4kJunEL+2hgAsYCXNlUGjeZPcK13z2fGTh0+Hh80YZNRHe
+dZtV869YTf7eS3Db4vTQZZsZLwO0eTGDseqbQqsQ7Oc+S2Kfg7bztbdiZVW2quh
YTAJRbvl9uT5rYK0b7NSK1c0uFxL5p2u65FkBJqcoPaZt6sXFW2gv8Lp7E4W65oK
TCe/tCCWD1AcvMsJi2js3e14B22jnVJRNEBNWFFoxQus5ke7oLLDGsip+qERkc1i
M5NB510V1/oX5n9YLePSniZy8hv1sXM4AojGozX2spimCqDY0h+haB/xCQUqxg4Q
PYBz+xjuLHE5Mmxqq3S50CbmXzQ01yh8AQBW1tUsrHoZd41BbT1U5gBNzfFD2mMH
yJafp/XN9D7f6bfMYleuIsvXnFZX9mDD16Z85XvgfAGXaCGZGZ+mDLwI8Cju8hrI
KP+56hqbRri1saVqQlZXBy4iIYRTMKJjb5uDET04nVuZxXlFyvT3QRpKhORemhzc
knIQLesfFV4aHbFGc8p5LK/chNtOKjJ57oEIBmLjff3bU8jbNIVIxb89v3/3hGrh
Q4hlaL6veUxbWzFyr33r033FEKpJlIgHJELr//b8kh4+LH3tS5PxqVjNs5eZslZ5
/kdTnyScsysZJ8eOgReizoAqD0VtBO2EMrux5+TQrbcyDtFsymoNrSqR9Bf8B042
OA7+XOaR8OnMAeG1WSe0dxdxl45PAKxJO+3dvejd1pTm1ukMKkmUZdBbigd67hsM
JojVp5bHCGT0u3NS3CnLFUqtIJDWIN6bZmsQTLQ+fX8HB6lNuZSBsP8jp76mcxaL
BVgc3+euojFNZV59xxoBz3+ZVAVYGNCG+S3MVm7q7b7InYjwtrggwOCrlc4UnaX3
XbSFglximbwdIuScD5CVfYUmmTGHlZjKmnu5GjELEAe1t5o/pbw5jEfMm1v/uUKE
H1VFZ3tcEWZmeJgH3PIWf1slDqGYFhCnSFIWlqFdmfPy/KBaJHBXeQ5kue6EJ5bX
lkilc30jZM6gas4KF/6lERReGs1JXqbTQszBXjLn5Zk15c2MVKuPbQyAJq87Y5oT
HkVjUUKJL8+EmKWcSg+l4TQgN15wq/j5U9FyVSB1jgH5JEM6bSasln8BRntvWdAZ
/R/sFpSY6kneVqhEBr0TW4qIhDPWZHiQdrSwOYAXbYA758IGpP+Sdv7C+roqT88O
mSQ77jFdhJsWbuyb6K7luN/XY2s/y/GEiu5DMmdj3igS9+Lu7hwXaNLY3i88ZB+c
N9bKEinnTUiAPO49Z8ke7STTHOGiQEwFaqI0P+poN9GydP6py8spjG9o9oFPXpXJ
szzv79HTeKeUse19NbYXvjjub0mvwnYpovutvzcvYoepDsgKmxnY1xNcJ/pWAf9A
JOYMJjlvP8nGW2fNGQ2McWJFq6F/9e6THhm+UkDUkQB/2HTGUAiEYHVQoAQz9Nor
8xKV/q6TLpsyQVBdbAERcemy5un2h1oModwHMg8m2W8jQ+/JUSVP3AEBpJHVS37r
clavrzU2uHtNaOLOfw3Wydsco0RISTfPP5AAL9zzMsLArztHkW3U0b4Uu99r/FPh
P+1QCFhc5vE2e3F04OkaxsdN/V7kng4URf93zVGZrkWJqaz6JBKuDXQTp8KV17Cf
saYf3SLTUnrwfnAh1tJ6VdvwAYMyCbxXEzS0BrSQJhsdI4u/1hfmkPbYz9IHrisr
1osjTVOGxk5EFZfQEOIqrpVZYgDrUSScXGPEWMlU6kV+3MckMWUjxQ/1AuvWznq9
PoOutuFFBEna5Mi8Ay/ZOvdQTzhVQYwaZs5a9PHjE7v888Ugc5YXiEH+8I+Y8VLb
VLR06dUKJJzNQE5InOYdWzLqm5wOXDKnAwvmWCoPieCyoF2GGwsXOSQTQAmmSNkv
NE4w1IrjTUd2a11UYt+tg9lyZkFgnZK/tNT3NILj7GxqXRd00Mh7OnX4GqoZS9WL
q8wV+pRESc3WKDTEGF2IPQioOHcS5SbcpNyUebvTCDCi1Ru+keXYgoQ24R96jbVR
9UVxaepdK4ypNxLepLCgEDRmFMpuSNk47aTTKK67zDqlnw0heNDwyoHQpun9DDwf
tSu7QAZJlCqz7jH/s6MGTSYQcvllyyVYH7WTm3pnptf709HlXxRV51NK66mdC2XM
gHEron70zWXoaU+k1L++QJtJGp8WuAy60ZL8Xp6OVwCLkZxvm8sQPO0FOdkgOMWU
eLsJm6fxQfgXqZpNVxe0Mp+oFVMuOjT20iCoVPVRVwYBhxaWkZeroqL/J9kB/qpZ
/bV02u20v5Llso4xRq0v5SR/sJq6Wt/bwJUKUeCJyj6V6VMiGyfACQQZTlzA3PLD
wm8CRd9TELZi6kwqFEKx7pDdu5/bjZijhxFGeIkzfNn+qo0F0sJ08BsBvxebFy4C
5lVdGuraAGv8nlgKzuWuLJaAKhh50X1OH7EJC4amQbv1JhMtLMZnU9e5QHb1RhmE
MHejVoLN3WTtIMuJxqk3ywTKrPwRnGS0gCrD948kvKSJJQDt6YdpK4Q4WkxGm3YB
1QLnh66lkEwN4PZOs3IqhApRS1etXO7C9yi4JS/G2kG0yoG1a3JDWfyTRkts6T+b
daYHfQHGlUNDIHNtVHID7+EXRXJwD+BKgRz/LlLhBSzEuUV+8HYNmLVLqQhNqfJC
3LnjP/DAh9adQ0fEOWS4P2R3CBB19z+aZaX9yTZxay/dScHEXe26SDhJNVCoUC8d
WLSbhfJ2hPkR3fkSzcc6Uc+sjqpC3FIxiqvTplKXTcS8RbyNAypoG8BXPdhS2jGM
yXw7xuuQDILIn63qb0j58Zv340Snv3kSpq8/hi9n8WogavjBYY9j8DHJuWAvg0Qm
e8UUSYqMGm0UcJ+vN4hNYENtSit8pQ4iUhQN37bw0KjCSAOkKbmcgAvUbh6aw3ZU
TqJMUMFjWVDGgzRgfAv6m72AIKas1zS1nB9CzS2+HSgWHJHK5h/R6NoclmxwmUpX
g0bZSuzUgiJEqoUyulJ2Anmn6jPC8wDj4ji9yo3ph7rW1CNzXSxJyY5w8LCq1FzE
CFfoK6c/57AjoEqwKMe5P6MIOBc5Vl+DvFV6nB+/B7Imt4C91u6oxH7JI/mhncdr
Mwr9QEF2GF+FZm/j+1qvjh1suquw24xfoL71fo3iSRrpm93sQ2k4oZ0Pg6eFPXyT
2CZXbQ7vYHlLe5v6+DkJo4Xn2MKetQAOupI/I04ZbR6ciF7NE+JhMvDPTvS2GmwG
90GRxh1RXw4dpUyXxat04r3XrzmH6aqpqs4jJLAASGxCno3Ah8gF46BurXlGZfxy
CxPdyUboYh76jCAjkUCHkw6NxB9s15aXhkojaA8SbsLHcbY0A6bIYlF8ahumUtM2
TAMzeYb9kbd6jZAIT424l4w1UAHChePMPmWy1TfQCqXP/l81wKJhK1ai8FTpTnHq
kRgsSDlPMiaFPhgB0OEsmOmoSj3tfR76vu6kOWmmKKkazzhVXP5wU9u8QPoSHu1i
Vt5GACBhbqs/jxU7Xu86CSBxWx+iScCr/lN+v1HcXKasXfacUQJ1o4kBN8QYZEam
GnPiTgXb7cseWOw4FBVdQ7NT/tyQP2VyT32eP1ztNo5zCjwe0/8pyfWSFBE2eVs0
ySTcYZ2Pq3KvGVKsP0Kj+7sdcXE8Hm0nPH234T59wHulcS8DKKUIhkOwkseIcotA
HgxDgf1sLdKE2fA8pX2uWpRzMYNwBddBwtfG175aNvLpbdc2sU1+ETxaTYgeoKwl
oAPhVzT3zZUXcQLfJs6pbQv3JP9STLd2fBYx0RjYMX3no0oX5Fl+TSm3D71PFm3u
f9Q6jUAMDellGrLpPkaBCgkCZyg4zoJ7i0T4n13fNyD04KFy9NTcyl5460tCGaMj
JlYP+AzIomNU/0hqMJlZ9KCpezLXMrbQ3+IcnanNI0zeOAKfT31C5YPwQKdJo//W
Kcgt1FSSxOCPjsqcWAYCt95m0BqnufXEKwU74cFzCOCuBvtbtXAIWK35X4DFn351
CXujsy1swANh74j8/KRa89wx13B6YTV4jiR3UpJKBymh1hP8Iume023usONHwvDW
EuFxrYaDD1+U0DxrefDExzXDC3H3kK0qYS809+PoKISfwxGbur8MFOplLVBSkePO
bQubkSC49U/2hFh0je8SXzG390ZnDIgRmvPysuavjdoG6tMtwQjx/NaB4XmMriew
ssxAYR8/u0pfO/27If7BsOTISWGL3AYrSfMPT2fYitpQc0H650kKCJElnhup+Xw1
DAdUDWM3WKnYTy/UW5vUXvAj2OE1vPDDxxd0e8Mt1NlvXhNNIbKSsZ1RqPgvZsWG
lxY9L6Z4UYsKJVg1IW6Y8epFG7dDEOK+zFRiWODh3Kd1rGTXAO98qX7AKqEq9xoy
6J7Esx5tgsgTGODNMURc0KohUAAkS9fLGRNCReAHT495Q7AMutOHLJZUVaVQ2UOp
w52+DEwpcSn8zZeMBZOVjtCSYLI1CKw3xzXhTlr1lK5A5wRw4qgYxe4PxaOtzya+
1cSPgx79asApawzxcpWqt44J7fVh8jm4fJOXXDR1h2J3Vxd/BvQQW1qFbmZsjd6S
07IbWN9IQUloCLbgfEJiU/8cCb5RnEbxAavTRuF8lr1lRRIxY74xzldb8zthdh3D
n+iIGiFaMhX6EVbg63a9V6oNY3hf7WfwNSpPxozspyhR1ZDANdtAGriwD7W9In6d
aAKkQY+KxXu71N3/jhrWgLVyBZzscyhq1PjIM9wi1CC6Xg7176rj598p5sdazK0T
1Uz7AsLwjE5zZRRa0vZwQgvNs4IEIjkIuxN5+FNuOd1htFxWn1yPRjUV1nrrlMkQ
0MwayVb7eznhMY/qm0spWzbHZJrsjyJsBlgGyB55ZtgXohT34Yk6W0QmBU0KpdW0
6w2b3f0XGC8sjKCy2qnuggDmU3bAw2xtjqZb0oXcIr78ewjZuPBDQi2yNn3gYCdq
bbtRQLlomfrxvDaB4vITKcJjuiGVga1QkdlPdDIzJ8hOjzlyrcSzdRin92D1kPLP
bmGahou0acOJw0XO45U06P2en9i5qipsOyoR8nyY/yRyLlBQMQ+qROo5PmyK1z1J
dIhfCPAuB+LppST88sPOssdRGybACaIR+gQb5pSuCXUmLN1Gq1g2BHX35722sFLC
ZLJANDgGlrbJ7UORcUvMvRvCA+I+Gs25KuPo97LYeP3EqmoN9HOY+7jedIm3r0eI
y02UG6ZTjTcvFBMuTqrTwIduTqmKUnMYaZnv1JB/YH47P7cOWaBSn1npALTnfqRa
y0RQDo4HwIig/L4fIZldHExbKDCP+wZhWHs3rI71N0yVnkXURz6JMV6b4KzimpQu
+Y7OSflAtAeefPDqIHYx93xWCa/Z61lKSSykho5qwIEMwAr32hGlQFKObCvyPwni
cqD5Qeas7IvNFhR/fZ0DEaRVq/5vGFu0Y85i+HqeSdWYjA/GzFlvKHDaCNir2jv0
FE9PG9oDxVqJzImJMKfA3AeNC3xWPKOaotZjcJ0Osa/QsVhg0GUgmFrdsRlcf5Ap
auslvcMgu4T8/XIverAmpGoyTg6kzSYfRuDsrzlmTUU7nZVaEMtRLlvDSc24swmJ
YHuhRcC3RUajRy3LYtCQxHXpw331xOFK15qiH6m+tJcjyapUNwrsgPWxZfr7Ur0Z
ehL4A+dcXXje5bCNH1UP5Mr8Dx6MzSe960bgpcjrMiybE89dNuWd8ILhyjH/Vlnn
fBXwwudOVTeNuUHaS7DiSWDjdNqx9QIVBcAHOLKn1lKdbwkIWnOKKbaME/b6nLf8
xsxhZ4AVbbIQpLjkqgLZgYNqgV7ltvRT9ecN78iLz4KmHuamBxYxtPf01RMgfolM
VHFewCJEaFnqnq9UmT0NEsg08TzzCCM25DpzCv6PAldnl/GcIb/R4imOI1lWDqwQ
8pZL+HwIhxYiB5FT7U92XNXVBv9ns54RuSV8//K/AODC7Auwc7S+jQdzCRGpBh0j
B6Y7KZAgaX7iKALLcni9HbL8BTqtd6HifIekPS9WO2GSbpguqrI+sk3wUl/fNz6r
z3TpyW9DO5g0oI13dzbvVxuied+VGGEdp5EGsIDvJ5NzU6Yr3zlSFOn90r04MjVH
e79xCMQib1LBtw69iYRDSVK4Ch/OGyEn6wspC9CTKTmOPT42xkNx+HgO3BHS9DbW
u27j83IzYq50lLF3azhZCvwXYmstVfIeCLGHlxAEmKp9ipBP81jVwDBNHay/tKGq
HoVes67IB5XwnE1HRjcW6OI1ivV/PZDXho6dNNeENpum0HR6JarRtLdOYRCdaKkE
tm82GFhLipjWhV2VIlvEJj8alYMdrZ4bhkWQsdDFEGd5VdYpxmnX7+V7CkWAz9Jj
zbNOQslBwOAsdhH2xnwbNZIAO0mxWemKSCDkZyDtbrNdoNNExsEfujYtINiyaSgv
0pr02jmUDcZa5NyYv3tf2a7DqU8LNRstOb+EyXtPdUR86o8c8FJ95gMBv+SeSUIe
bKVZlCc/8iQSn0zsZKTofug6x7vKaqTiCMa4FZIm+JZEAhw/nP5Kn7XqlwouJhRB
Vrb8ba6mxOrTBIYeqeBDe8GCF7+CpypeSpqZv0fdSfEYARfU2YHElMgTi0bP1RBk
bV1bTjnraDBcaA/M5OUrJ7KfVJDp6Jmy5Tp7RKHxHZL2ytwU/fWmTQtUvzpJks8G
KYoJNZc2fPxpOj7n0ufo4/Jy6iKfuSIVlQ4WHOu7XciYkXHyBII+NprMKxcSDZkH
nD8Emt6skHUs6iZAKGeN7gZ6Auho4NML1tlJj3eb7quOd+QxE1gy7WwZJ73nq7Fh
V8NTibmzwufNQ/G8VcWYUHYGkrj68JpIzowonxR+5+2XPU2pdfuDBz7xWqmLRECm
KmNyZ5B5TGIlyrFSe86dnAlpOIJ8NTWOMkxQVg3skLvk6bl7yusuPcCW/PM6T1rB
it/cETYcnhecudgvYTNqtg5idz/8CDWiyBdOg8M2l1rDZElh6aVYi/zeUi+xxDOc
xhd8JxRbnvwEu8xDN4rTqLrb2bJYrBlHa6g+QTQgQTNxVj3HIrgiaVYmZ5m9Q1Q3
6DPCu0v+eupe4sknTINM1i4LNLzCYeJSOg5sfIkVhl5bNzyz4RxDulJzPOh5DVo1
PIMu7m5vAzMpRnJjDoHAHC+dQXjm12rWMounlRZvPVydlgRZuaSd3hl7NgkcvkLM
ul/0X67V64rE9TwTxh5Veqq7zJw+3Rjhh9PPIf4KntjBp61x0qvceU+mOolvS6vX
dj/e+e3RCU3vn2elLVJdQ+UwrOIfh7kGNMn+py7WuCt1aFjZONEwQEIaEJta6I62
rKvGcEciH0MFfr6EICwSwNvHdtdYymLBiu4fDqBBrp6bIecyCFw2GQTN0dutIQUI
f7P1GMGE26ypHXkFhVNfk2ZDacjqyrUm0831dZ4EigLQ0LBMUE9chNCify2gK1Sq
nacOAvmpMyBoiJMyTECvAHEiHGgCPSK/2jqFRgV5Lop5NT2RyaGY+QfecmF9lSWX
1On9w3ITwkI6lml8JdBunq5Lu3TqN9AfgmlYw8bhbHLkiXoapHwnHxN/QUPuJwUj
jO8aa8y01ouBrurQG5O7dJoFojl7CVTXGo8LUHNhIoUGRc9LKpxX6UCLWvhreZLT
Vq4qEe7pwkKsHfc4YYxkCwC4RFsfjEqvXAc39szo0vy8IBniK/zp8NZx7Z9rdbgU
DgtpD6nu0y5gktm2Vmd70feR7EWlzkNmlaRIWqGtE4idMjl7dv/VGi02jjvFyImY
Sx3oVma5MFLtIrmD4+rZlxkC/Hj1TXyYmDy33HFgOBsnGFgog4YzBcQFp/womA9A
UMRWSgMytz+A1a8e+s4wjVHibFTKjvQI2X0YeNOfL0huMbTnEdqtUqRZbPOE+VbX
zmtGvq9vfimab7++t47raz2ZY/fVevWvQHjYqebKNAqlD+teapQmJL+Uf4AqSPaf
PIVZ/QzqLDeAerT3fzVlmYk/AaZ4/J1onsm1/kQZshDm+hABSPUPtw5bB8u+6Wl5
Zbpn2pXfpnb7oYCE8aFEvLpP3j3/lgtkNGTgDEilTXImZIJ7gV7DofwBae6Y4w/q
9e3JNHfYT2nBT1a7MCVxt9k0MZ4BgETbi5SKarfjz1izj7t1ffwSUHGfsIIF59m+
gf/1eR7ml7uI2UG+pxXu2kNDIlPZg8JTvpN212RDlqCi2pKPGhJNEFBMewuXGP+k
YKEu6LCQdSV1WkowdWoaq7RMbhl4Te/PND5peE5qrRWaB72ekQGcTrjRJYxw9CBU
ezMivUSlZ3CVvMypEdZaXVmauhAQe9meBQVPlj0bIeAO88xBZLrt9Y0giOHo0oYY
APZGBH+cVlWd10H5zvZengaY5Whk3+dTgeXeCIZrEGgPVuopx0cAVn8FkttSMIHh
tRRcz5N34r2Wgrc2GTNxBxL0n4uL/bhYa+qN7EgR2HhRr/X8k/UOH9CB2J37WmnO
Vzj/kEC8F8PT1kpWUGiMdKwWLx0VCB1HvR4pUzdXkj3Ar27GzNbekujRyq1NXR5c
zkbJXc95J1+80bR9Jq+mgxFIA0RgWUaZ5bgPzesBGdKqt6LFwYHqsBEfzOv3O133
bEQxKO1NSd+cbTdI8NGNXZE9sMUQLQUMN1VmFtf2ioECy3TGc1XAxZxN3YgGZz8J
W6+Oes9oIV3jGUODaPkh02opRBghaDYHyg1DsQxxJL1Uul5aOMxZXOmCCXj/lO1n
421iyYBUz4h2IplYnitI8d4pOoScT0+lxgCxvifarJjGe2nmxlVGEIs8Tipl2Swb
XKbGehEi2Ykf0D2G1ZNpZfzAVFAcjwWK/VYesjsfOc2uF5tvvAS+lK5OLwA1m0Op
z226H4JtBTvdls3ElZlcsxHtISRn4N2CdM07zIVj3ufaFIkd8mvGEC0PDT2Rz+Ee
yAppS2bVwzTSy6CRRj1sZRyucgvs9Ojk1Yh1cOEOkhk8kL8YD3ouJ2nsixvEkQhu
CwWSIlz1ngg8blLUyTK7GNdXN4a4dm+VYABwgOvsODXP5xxUH1y4ua110FWIj6b2
W/UI5FrqZnsfeV+Z0T3oNwgb9THWfQnUE3DdJbpRfhxady6zWJvQfJdyeY8bwf/l
5l69wwwcD+dVsjIyZfWDuwWKByYUx3hae9D6iG/hQ5mGzLdaJWnIC7ksBnlORon5
DbyVHJxIWXl+JMoy8fi1uIPrJeMfjKNw3GYQS9VZdulbXbCNk9YHo8F1qVQFYGAI
PBKsl+rSqCZ02s5q/q7w0xDcx1iDbO3RPmNjJVNyuT4P1Wp6uNWSRBwZaojJtmjW
FQA3hXOagg6luo4YYRBUPv6BMzVWrr4p6P7LYb4AoM0iKtoUXf8c5VeCNmBX2Don
TbEW46r1o/3h1wp1yba1pi+XYwHgWmhN93B1/B/fvHFU6zvb+NfaX/FM7ggRvq3N
SyzWeogsCz7TCYXwLb5xa+RsEoXjJ8G+X8SS7k4OtCb3Jv9+y2U3wbb2Wpyt3/ru
ed44W7HEpUESdXXRCoBfN7UGBuzGlTqUglMaYcfSX+9mKtEMoHmsW2vQJNgf3INN
DW/eDMu7snIyrkdFyukYFbSqtA250UuPvD/qXqwEWTGFEVbxBTQDbO90ScKh7fXK
yDYpVcSIqIlUdePoy7PrVJCULKKKOQXaL6RYFRWLWAQDxvsO42YffemINrBBPPgI
b9aDXKyLI22LmQ5W/ktyX4niRxPW/cotOoIpaU95+rkpDkXKCgQ3CeyBsPyYdy0+
cV4u2ONMV4QkonKr7MHA34/GRR0Ole/WNZSh4ZEa+1ngdzM1v5/nce5/nOa9vDMh
YcMzO8f65LpKRCsrQCzJWINJRzExMrH2Oky4tmDuGpJUtJLImj1y8uInWPPaDN4X
fC9bic4qzC1hRv5XTQUL6PdugnGJUdhAkMSOqczO1x+I3wmNiM5fM+P0LLKEHdcX
PBTOQEiTFOL4qBzuDMSz4StaMmB31/v6p6M4VWEsZkAU0tDlSeXqAZCJeghCor2z
4YbcrrEIt3xKfZH6SPr3LaVoG/2xxVTpnF4JNME5mb22FQ4HhYHMAi9MyQTXU8B9
pH36PUbiMR4mLU3sdiyCEhYa1OL3gvDrveg1IrdA4Mbw3pP2bw1qk0PNJSdyAls1
ASmler3L8w4uTliUkHgq8FFhKyJJTWLGSvxoF5gGpg+evFWl55NyHELwm74oGNIP
1NcFF0EPINDAvu8Qqxp9Vhhv8OahYFKQFuEVta1E7jMWphj012nhmKhbVQJUAvte
VckN/4GU00Mtrs+PzmFKCDf8W7IpJePaMUiR9566HyhM3irWFx8rQXKncERJw3mb
h0P5MlYb1xUIS1a0XNAr/PSHsGl9O1nJoy2izMW5SCQaF2hA2eVhi8IF+1UvbJOq
FwUkvqZs4xyTSZ3m4S/jvT97/kGZpVW700LDToyPRk4jkPJvM87RBaz2uMS1dp9C
bGGOXwwyIYcrAKVe7C3Vwj7w6wzV1y9imc+RTlqhW6aq0NJU6D8CGhXRATutve7d
/rU+SJ5/CLBrmLdQxRui55OORbZIq7ezX9BVosKfeTYY1UkNyeTe4y1vgS1Olaf6
rEGBHBnAX8tVagXZrvWU2iDFqtr7LbhivPCevNy4dI0BvaKFPpW9SFEpQ6Cq0FpA
21DUx0HpxhbkCBcMXCwfFvinV09zw+2pp4kbQK19Ien7ohz1Clg1dapxH+vjVaC3
RalMokduwqSOvul1XS3FcJjYus3/VqMygR0AtSQrVn/4thXfmTRxAeHDo97VAgTb
VvtqblMdfoHdNdQTitV/QXHtMNEDuNT1YDxDLhXGQWrNaDDkhJGjx+fdrMDK1VsY
Ukifxec6O6yuqnxZp7pu6u1U/bGIz+9/oNKI77C1J4aNgzAe715HaRwv/H0rG5/t
6/fBLqmn1WW+C/G4miASRksIbowPeLNmwF5oerWy2kjMd/ckAZLuW85iJaBij3y4
rv8wUCP9adIK1WyqdUzY90MbAwxc9/eNmA3fIVgJKqIYHa8FmBYSHNK9RdUbEVuv
sFdV2Pu/WnwBNDlXEv2afbZaKcb05nqVu1JeTEm7g1Jnhz5fwM1kqaVKbPUs/NYe
OgUaTkbN0bwDKKG6CYtwg1sJkTji7NBl2Ws8eN3vGvsJ1y/1MIM1Xs+0TYI4ND2W
+4RaZn7usR3eaULxjVOR5MQD0WrBFvyjhQJgYdg99uuemOlpq6ebwOyXg31ER/bi
yBfUHii5/zLabQsFLyNDPr+fhTzlkHr9eOIvwMJ50CiOqgYbsqmrW2qGpk04G5Ie
tbRNr0m4W1qwkScupFRlf74ICADJfEUKbxjDeB55brgzo4rXpvX5dpbYUQryrjvi
3YF4ecxeMdbau+bncVZrqv9m8DVB8a/aS5KxFVsvvAjhMgX2zw5fxGnKZhaB03HC
uonscq6CwTY296sbtAExOI4KbyzwqMenppcrUOpBBrUCvB/V5fo9QoCs8q7S2ZoH
SU7/N0bJdzVNoJwDsG7O+ZDf2NMLB+bo64C+DIkgBIjSAfRisDG6cpGyTGSC8nfw
dSPfGpD2EpsuhzDT6w1nlxcTxJ/X5jOsJxRbm3mwmSF1ny6Qkkbe3wqsaUcBedUw
JZuvuhjxYvxuvCWHpJEzz1gG+zu2lbkEatTTL1F5CqdMQYAuZ3vjL9s5tk8yYhLF
T+HRAn2Leu5/PIYp7q6Cy+AJUgCuaRPwnIFobCcTEvSE6dSleRDQpQ5yDHHRca1m
aaMvgYB40PkBGJiWUS9B7haMoCJs8Sss7VSLds+MvhXx1qz9OMzaQy6IpA/uiNZ6
hKEg48kcNIkL13QuHKGgUTaB1/kScNXrBY1o2kVBTz6r+oIfYDfqqLQ2dhXqIyRX
JW2z4FyMakslAuo9hJQehh6eNTi+XsfgmJWv5tu9V4RDWiC3o9Eqfl37frQvA0yp
nu3kn87WKyzXXyiySG0p7teOiOJdVAvpIxozx+kToTZQoIdNvx4PTEeraZMGQz6J
dGKSgQdsu3+jK+mYAZ5bUgYIaPSaK8d+mk3Lam7W9c3ngq/iwPlmFc7dseDBGUAR
QAelp4kqPHJA+VBouw8kCIpxPwqWVPIAF9s/FKUjT2hezUOfM3h54AaftgY+Lhvd
KGSDmxYYeVlZ+TpUYJKAFF/7I/c2z49o8XyuqRDp14CHSM7Kvp6dK+vu27+5H08+
9TLowZP3BVsFm6fNlmuIg2MJJa4XELEo/B2eiR9G3prGACZvIie6bkx9CsT96nWn
C3bDg/jFZIHgJD5YeFPCqk4fykeQ8RY5gxjIuOVqftn2eTGZt7RPCOgftA+YfGom
1SyxLg9fZTxnxHiSQRTpDQgyeKDNpg9xpNfvQj3FpL/zfdxQ4+elqCKczn+JvvWF
lkPYlSgybgOdKX4XlxXfQ9X8rLEh+H/0wcH6ZD+nzdcZ9391vsSufvIzQrCPz66W
F3bSepOUiiJEFtbxI8daZd8GzSw91tt3F4T6NuinLK2xozlVnzZVVRPU6TAi3fKz
5sWSa8Ql14qsrXqPQCFgeMjzVWE63ivpJklPFQW41zsw1s5J1z/pCLr49cZc19uH
4BigIZiTLvCBOaOQHoPIJPKStdghnRxnLCwPsBYH3MLv45smuQUr7wrJhrGpIjC5
LpqHk3k0fxPd+ABa6v6Ceg6xXaKdOZDbp18aMci/5XISsL5I2PdD17lFtWiMhbcP
M8NDy04OEOk/PluN7IVqY29pMPNOEptjrP3HrRdfRj13gJIfr5oVQGvxY6eqHxyH
GT0DehxdTKGJCF/0WBleUb5u5qa7TN95scjh0kui4qFsh5k6GunXnCoWL8+nvYtN
nQmS9Y0QK0ynPROFC+61tp9RxdOrXgn+vaI29hUcqOEtbWimhV7x26YBJ4sX/b4j
rUKlMQFZNMgBlFhqgXJ+9GtaJqVnNrMNwRAaZ9/cJh9uJ/ps7nfWKWF6aa/yFar8
HMZ1qzW5BzgpLXSHh8uc+UhYjm4HZVsSCYpb/94mbpJ95u/p1o9hIC7Slh3MKKro
L0+53ZJCkH/sK3+CyEpWGXjszbJV0SwuhkuoBYVzD4c2vn2dg2lkVJATPw4Yc4Rp
qxPRA+M3T/yMr5aWVe0Ng5QrxJENErOZVYZxC/uBgIHUt516jKVqz2wglMzjvkzK
3wdZp7exzANACrgqHyNwD7kNaJVXJ3cb63HkCpxN5hDVGtorNot1BJsCa0Xgjk3d
OoHswEgAbcq4akC3bTYdZN0oUFTJ7cdLzzuaXWImRBC0jd48m8QAAMZFRoR03aqC
9d1yo0/YGi7bghKvUwQ+5OjA34yl1py6WMZRyYmrHBod0KzPPLU72uBupJZRkEpm
N14c/ZFSFjEA1atHgQYbgk3vNxIPgAYkobgOS5m2PSoLshRlaQCG52OeX6y7YaC4
mZFvqHZpl/gbx2W/oRuXejVU4Of3Q/Q65UCA5Na0d3lgFLDGcDPm9UxKTrHds7ro
w5TRAkbRo8vKg3nZU9P4GlCgKS/7CzReq7WfOwAQVY27H+shObOX8BmeolT1NQPS
SM43pk5eMPTkPMswkvYhvJhqvpSfCMAAsds9/0tumeGNmpkZ2agFGbCyQFa6lZmF
4eNDerWu7LE/24EavRk/fGnNbFDL6vXaDZhYE1M+xpbct9J9xt/m41P4mjzbCOOO
kpD1JEjhkWjukKQMn8bZQOqIT8f2QilYKMkCFIAs59sZv0+AIlICU9+5umQlxfcU
M5o++Yd9nG5dKQVxZTXhnxjHbaf7uEEFPFA8nuSA/KSvH2glRAc3baGx6AVERm/z
zdux4sSdClAVXSVYMGMfnW5WjZiBhnX9kUYq2yojcRm7uEbD/rsXpA1ALSJ3YSkJ
bHPqloq9RWe0UOn1AZgESQXLjMt3qo76PAZa7aTQ4EyUz8IPH3TQvcLvlJwBidSg
K3Bbv9I9wz2+zx4X/CXWERh7WAauc+KEjJ4KlnDsjkZJeOX7IhAkuzLzwQDs5chV
KpS/i2/o28osQbg5p/XAWMPHniH7+lh6jigcZ3FALuCDDlKifHZPuXqpmU7NFv2h
po9Z/AfxjuFaB5ojqG7s9U5HUMxt0XviJVaOAIGgO7VNkxuKKUXVbj8WxJMaHmJV
gzJMUjG57fS6Fy43TCPlwHjdE8Wl8F85kV1EeBbuxSu8dV6TMh+DvpjVXEqmGLMa
LLgQb90Hlq8F0cACcxA/MjL5C3p9kWpWghTEQTCWcDYMKHto2s0gGm3lJaxZlfE/
dL05u5BkEY9xeE5SuhPSewlcjs7fck16qBUAkrSMpVrFdiwBnJxDtX2GIOAvFjun
Et3RQhUFmdgQF8Y6YKYrOZvRAl/hVeVbl4ke08+6UqzmkPer7VBcn56iq+Kt1Fs6
sluUhOl0EcOvlnUWhl3aLStZHvPQDEjPjIn8XF3WVrUk/xT++bHMks0YgianXKVn
BWgKfsRZ4IIuMTjYlTdJHR4/hLaOh4XxM0SfdJSHCtw3WxQSrb+4dFLvbfcS5ruz
GMYNqgJXC+nwHwstVACD2Bn+Qh+LJ68jzsdv37gLbZnP7Qo83PsJaNE5NN/FyECM
b6fgjTMVdYiVzqsPC/iJUNoEJiAoYeYYESn/tGVda31d7/7RbSAsxHsW/A7VcPN0
Xt3WBzjlC/YvZO0KSpF6HeH0j4QdraLkfzwp4ABIIW5cjrW6iMQ4Q6v0L4319r04
y1fMEySnnTm+qHbxfAiMWURCbNzw/Phx/0n8IQW6QBLQosqZsyAG/wlJya2JJjhy
yL9uVyee3/XdJGBJfU7d5JewfmM33GBWRj8a2QEm1XXjHfa1DmDbc9nCcLe1vlaQ
PdgjX+6PdVv2yZmAQDHBMvHsmol8FafIggAbvvwIJV1BNTnvVNMF2y2ZFokPj7lO
oHSH97rkhux0FUiidxeUfNvBOV9jVGAF2E27O79x2xrav7k/KF++wcq9D2ChBIp5
RCgW30UhXDFFvrPgCkDXvMy/rwjDX65PQDhbo7S4fVz/ZS0Ec+F544pg1sHk1gKX
5+BQwoQ5VXCDt6YC5k/t6qHXC13TqxWZoyB3arDaB3RFD9M3TVTvgKqyyGkhhbZe
wosdCyf938ZkbnunmouHay+P0mMbsuAkaTQ3j0JrV3a4r0VFJ1yCQpW9heS2qvXH
xCmxX9bTNW/87CSbgRD96qcrccvQ/mOiXrq0a7wCiRYPrx/tOh33s5NMV85RaI8X
X0xLR/7w2YZ8k+R863uhzB2eyy+1V8I0Dliu7RoNcmcJCiPwvhpdnQ5Yb2JqvEFt
GWu9ML/cgqX44ISjWF9ZJWeBhJR/1+70FGHu2qiX8d4zMlV+xxhOEOG7D9ZLGUW5
czndbPivt/7+0uxRmIyu3AHJA8lYeLlE6dsuHDkmoSmfzGhR4Yy4QHYBzUrRws6B
TqQV7A3/iuh1kKbw7M/aaAazFklMYrmUKx4vESHz8Z+CLAdi9rnNTKVUpOP54UCM
biiEihwV9TM20uT1sAiDYFnV307wjzwrN57/MjqRmr814OGv9yea2TiPpc8MXQIb
9ky9/VDRcN6d5JOAaiFTDUbaaY5j71nWO5sL5KSDg+XPownXDwDC/R1Y4305PClt
aWbiWiL9M8024+eRevqYvecVne3/y/UZHv0O9iyh/N7xZIx+nswJcRD3VOXzdEgd
9q1jPglEa/SUrZyD0A6U0nZ8aGP2v54MqkW8Uv3IAgnc64OTIRdqLj+Vn5Tu8OG4
nSYL/VeweyFS21VUw4Y8olobvzmNI89pwWeG2J6dRi1/gKkXR0LzmlECkgkMYydU
hANCTa1uYwxaKPg0mjtHHShUVIEXLsGvh6OZ9fWXQxtZe7K97654gd0XxzAC8HTH
axzKxnsmOaMuoFDeTEHLymn6zVEwOj5mA+Z6Ot1mNylVdB4WMsVW+RgQRAUJu4JF
74sxpmC6Rr2gScHAjH6ouAn2CbkTCCdSRB3lo+WS+Dc7bpo2WWeJk23mLvdx0PgU
uxVNslQC0I1hPWSdhbciKwKRFgtWK4jCvung5NkiITtMjW5135XFGo6ic2sH5eRO
OFBnnBFcdDdIgw7Dmp0HODLF012O1Azzf3MpmwHM4m3gMQCQl6m7P8S/szb+0fJ9
Evy7LtqxV/dSQF1/WpnFl9COQNEWra4yH7q3sh7n0+Wy0aqTgii3THwns5VVVJ0b
C70DOJPhxFk0GjIFSs0zVFqxls0jAzTULb82i0MTDvvlSC/1D/FESjy4J2C+cw/e
0r6Ud04X51IeFt8woN+h3cIDJ0GT/yuQuEtZEP36fihLzFmdjbcsN4pDxLsm5uI/
xMuBe0NLEcevX1qSZPLw7CDfsQ45JljrgR3W4jWPJIj16BmIB8tR87T1rX6pj7tc
+GVlWMANBdHcsCUuuEf08Anft6v9AD2S/yV0QmPtM+x3fMx2AZsXG7nnZr+gOl4f
6/CU144chcm6xAJl529mzV5leAD0yxOpmFZQs6P6f/A7dHOGzCdYvFZjDfPrvshK
DSZR4bOPFgow26qIAkwEssxHHe4Z9jqAmq49Dt6gdS9qz448XCxVQ+e72DzSkWZU
fvfggDmx5KEq/LkkbrYnR2vnzs9w0+h9L0o9yU3KDF/gVFvK0k8TNsk1RDsyGwaA
tg5K2JTKPsTjMeSnWnvVADLRrizasocwjJAA6jR9y7WTMglJXs7zbiNY7WIYx9S5
4aqZftnFPGYjOkCZgyYYWsIS9Nz4ihK4sQlDT91XIpUNAxALmNbyc70HJg7Yy4FX
azpqf7PoceIiOt/gPKt4BJ0a79NXZNotE+7MwgRWWXgwLuzKlN9nFjA9sTGGL2Rk
Js+C7wXHJ9wxEPLBeHe+LyMH3PwK93PQy9xERdm3VB03xKePwNW1UKBrPbl7tlY3
a/+xsoSkJqMBFbjB4Z0/89JczoN1KUe0tWcdtlNgHxGOg503upCwa4cEAhIwpGoj
TzAHVdhEd2JtuFChmoX9TUuQpqWcW+VxpEzQpN8FMoRSsoTgd4VI/7rncVT0RfGG
25euQxhesMuCxSQf8xe6GmT5Z5wcX/84t0j5d7j4vcE7UEKIg8Q+Vko4pQrRL+el
PqfvoDcZWNl1ZwAc2eVHfGiEF3gvuOD49yJzIXDZ4WHcI4ads7mMj7uj4Q/28SBn
FWtmn2tGMb6akUeW0XDnrq2vTuIi+sIspZ/IgRnZ3Rl3UWjk9P39RSIYUv5/ER7W
nd0fVwpu8vByQDRtQsst4TwDO8O/iN3TuAmggFBRaRDZgU23eIfuMS/jW77YYVSM
bSGzWly/+74gUbPAsENm/0uf40iayboNujKaUi/xY5v9g3AVbOUcvTD5vUGrmPY2
GOqXbbROuFY9sDFUP3VQ/Xib/0mOKSldVwVNEzQEJtg2ew2pXTCa6yC3OuNHWoVD
oJQP0lIW/wZMB/abOZpL6s2Y4p79p/vwb19e9gXHmaLkq1BCHR5hgwZFbJdCdXuz
Ti6yxO0af9qM4ElVY2QXF5yJjjIZM+uN0WXwNAX6IVFIKN77PWvW0nRWiDA8dVn3
fVi9CjzUbnOVNzAhzcR2cgVkJ46uGwvy7igEVsCSGPUHPp2XeUvZ/dzUWcYRAvYq
V78U9gKK7X6QznQBrh6HxzMU39LELUt8vPV/iczMqfBuN50gc1jWvokH3rIJV4wJ
zQ6SwLkrpBAOawdjoV5bMfJBRWkzzGmOFebu1GdW+UPjXCIBgdYr668amSiNqLVr
46IypRsqT+ppUuLtrzArrGQiQBZt1w/QupcjUuQBXTTPTnJyNNkyadY71F+gcw6D
KtGNqf4pDCO6Ezdf4oP6N3n9talUG7Rad7DO09VU2qmoE+077YclILm5Kuc6Exad
s0fswF16x+6YHOYatvzjOwlI/yJu4hW2FYo6lxyza1/0dGT3W15TytBfhAsbSJ91
8JVBCaz6qtb2X8Ytg2mcENFOoI1jZypRqJsxVRP+zqHQgMxLx/cFFQSLQ4qACUcP
EC1EGl6MBsrDFGoG+tOxuhoPFf6MplEnaAkYRyMyZ84KVpjuRSHLffBOMXH+uonz
uA//3hNzxQrepLXqcz7jVkMeJshkqOZh6PrzdD3HphB5vqi5Cyhj0wlJyb5VZYoo
r1kLQQLpRUXxjnSKkTDG9dRmzpmnsBTYqCZJsoXAPt3vHy2QykZGunT9Bl5jZmo2
lc1ko7JtdG6C221KYvc742s6H7Xkq+S9B6HYms60JijCH3OphQw2LGiwAJ9E61X6
GQW/gsqocAE1aQJ79dRCM0gu4Y1zjMbzsB5iaCt3VdWz64lHPqQYkIDGaIqwXBTi
UaA2ve8VqKB9InewFnqs3u2odhOIJb7t5QtXOIl6MEJKjUYl5mRvtFIIrkfEgbU4
ZQ7exVnkf3R1yTMw19cFH51Aur2tPhMQV9tKRUJ5I5+tc5WcLE4M35KQwA1y06Gk
nHYwkcg53He50FQG5AXkG6UE9Ih9l5dN+eB6LatYLImUKYFotOEXifK97RXFTKz4
y8xiUVS7RfQru+srjRUSYv5Q1OJvHKqVjfofdS5ZBgYHlGh63Gr+9qwjsPL3hNSl
fRKshmUrXa/9qci+Z5VqKo98aSAY1PtVUxCTx/FZ05k7b2e6SR5ewcealLbDc7Pe
nnkY28TTMaYEXpTZQosCccA3S0/fTxMijdVDrEE5d3uGRGdLsvg8fqBUFEIKQL04
0QY6ACEu8GKqbbXv6+D/YSQ+QBJBn55jFOU2J100YfMqqYZMJEVenDjPocK9kA3l
BJHERP+8U0ZnGoaR0BcPZvjBpVHvVvrr0tWnJ6nx2o7o6FbD7NT0R5vJcPS0W1u6
+Rp7sNMlboUn8EdTtjDvUj0H+a2N21ITwolJlH93w8C53wwLe7kvRExksEpYofnE
l89X1Uw8oRykRWSDC7lnAoVxQcz4t58Q+19Yglyg1TMbKr16SBc0DPDP34SwU59d
o/krOHbJpANf97ioGscIXtqChLA8uPm2BJFE2HOlavl3K65pEXZS1kggwifife5b
C8a4EDqssySD1xr3Qwjv2aGwdjD48IvCL5ia2vZBXNcUCDv/PwjlqoNSe/Pex3oz
4SVF70VlkDBXOjcrINAKoZX/9MyLAg6oL797ZLbIiEqQj0EroV6+0fd7kkPKyMm0
4IrF9oMBNNXPnsunosGMY+lVd4J+wNY9m2fVhloKapWI111YNgnLcVkcHP5LMr+r
8nnOn4+SBk8U5uMiS5HVqtjbTZv+5zK36PhnfCB+W/ei1Fnv6Ta5lrH3zA1QRxM8
3SioBLmjSdd2+K7HHqVDAlk78uc5uu8vR+0l0m0TuU5pJuOObYHKsNr6MqBkB2Ih
XKncqWc6mveTHXwSNHDaLgqjnlm7xf7OXoVpWTjzhBg0KGQmhB7mAO16TwgOeqSQ
ARBg0bNYLgHbhu6sRV40hXFkYKaKWRsjpsicHJKBA63AgGpF8o/Us4LRWuDy0QCp
EMD1s2qPpes3WbCNCAXSKgEjI/L5ZFJzUjUlpcUxcKbLsJFv0Z06d2fE+Tle4VVG
qmsRr33yPqUZBuu/dwDh8EpkK6iukKscabR/o094aaHdjwX/4uzJ+8O7MxZew5Zs
AUwNqeH//lrY/app2v0vYmx3/OhA+rEBN6n4vwbwGTiw+F74/NzQsSJrGwvA/o2n
ysx+ovF7unxX8u9AtsaCt/j7yZhQxL3BToUgV7u+GgegySdV/wAQTIM+dxtzmjNM
xxNRJcgw42bYPfsYAmEfvogmikmrgQe/FrFSoU7P9lU0i9kpMMnpmsH9gsX3KEl8
2ZsZxynIFTjXyNlbGl+Yde+joOngUj0n23Y2y77+351FxGReTOhL6fV2vJSMpP9I
V+g8Nv23TRZnQTf3pOfrd5wcWjN7wYdMcwWUUsVOh3Fd07JAOs9UWevDiaLh9x0C
YEUXtCj/XQhXtHZG4zWp5KR9gIYpDg8+PQXxj4gcOsav7xaeccBveDw4LuMpOV74
Hp4TqlXPV/uCWXlzYzT61oRCeomu90HZMJD4NZnRopFmtXFwY528tZMPBE99xOK2
z9qR/fRuiYiG+uXsivkA5LAVbX9j8Dfhb/VJ7FJMXF3//E0p45atfLH2F3G9wcSY
EEcXPiWDZvWnq/8h1B4AhxxkTzDcpKJBxt8DiG7HKQf/69g1jnZTZBbd+sNK7RPE
fXLZBafxxle3kXeBooAjjsaPg+SiZwl4VuYYlUt0yflwxmRE8xqZXA/8pZvJ8fMr
M1wSqZy/AyIE3+dxiSF5SpcHiNYuoNVnHsRoAmtGC5xuRsHYjocFJN4i8VfDnUPO
1CXQCd9M4AQTEsnU7/f95IfeHmUgTPV/v0xiDXA7E+ZPbFvPxG36WDQ0JYNUnmMT
1Qo7qI9rViHJ4FVukTEC5IAQ/1xeRreWtEyehHGj0Hprkuluftxegq+eSXwG5ZPg
uHQ3XMmEPqWFaWhHJ+qy4FxW4I0gkdFkIHyhnr0TWAdQ5Xf+0HMpiEhJDE6G7xXp
oLMGBF79gmiMSsYNZ20cX8yHzteGTOVi99Dd5qdE62N/M/h6uKQMMuFiLdYB5kVk
plq78GefnSE3NFNfxkvc7G6ajwWA2ESQcarkP9cuxL8xoKhip6QKzuzWM9l4YMaO
zMpy7WmR/dHlve8o2VRgobu9YyY0y0P+Ax0n9UWySmEXHtspefVzEBZfw2OnZOA9
MQtb3VofTxtdxIdlfMKtjnjahVJAg6WegnnPo81E71itItXDfzyAOMD/jnlkE4wD
JODGDQm4kV+gBj4C6PPIJgNs01+UqTBS6gyrjijDpSWTVffF5Hf8n90Z2NXZ9TSK
n9yiSTMvAuQyuwshWUGtosBUQ8l/gxJgJtlxzRYq/GAmgGoxpI+yzEtBsG5Tseby
sQpivlf5ObmhUkE3x8yyxB9Qltdi1qc9PDs9Bl1XDl82SB7/ueFfL8A3zPlSaF47
MZASCFthRJAYzFBdf2XXKL5Ymixlv4Cn24eZyjsB14uTdhWKywudVXeXUh4r/sCH
vzOLPEAcUauxovejIz9KsUEwOG28It5t/+z0YF9nzW9zl1W/aj+pCOO2IYxSSqCy
FFQVaf1uX8U8rFOHWQYSZtkpgy3kFznv8C7+7pvw3CYN6YDTjN2c+JWM6hLJY3Av
9Yv1NOBZIFf2/wTEdg8Xlja0QH8FUVG1X1j+kFbTh/pv8S8Qz78pbpGpen1EeqWO
dk6vmDKBQjQCbKRqiJP6LhCu2RVU7dQtYDMZAzsiiJ3X3eATbRZHwFrX4l7+pJin
nU6my2vnS1lU5S6DR1aE7Tul3XKKGjS9iwLTftVGAbLkDWFQxZceGXa3x3AbiU3U
m+E1f2Nzw3uan7wIIGKLfVsRDlAnkkwWjPGkOxCDTyOi7PM6jtnN51O+Cd228OLA
xh0WaaQ4oDEzhbBoA/gjqtUrbODArISJ4ZhqeQ0Xt3A2RLfFwc9ZvaTcW11tNTVO
Hbbv31y1AqwvpdIqyMMtB/++/yGg+ndZlxp8Mug7znhauVE18yHKlMv1suTE6osQ
QLY/6FkoQjNvxeNX4xKFRfA3nIbOr1IiP4pJVfP7gKEtAdT/ChXFvmcUCnde3JFc
aIHBhyRF81oN+yvkge747mPIx9ticOf+TQJki0a554C2YyFPpUcrQ/+MN7M5OK1Q
rKXDZE1G2hLyCreHJAc/NQt/pN6sL2KLTFsetDtENM5lNqz33p3L1V6xEUg1x4MK
9kdC1/dDkAwtf8Gpx1bY40KdlMAhX9zKqkgNHxhw0QyOpF9evcqQvaJli/JZ/Dos
hqTii9HgMwsmThNjmBFFVDCclIuo8Zaau3hwuYogF0Tb0MTUfvqOHXGRYdYtdgZS
CWLWJIbHKD28f8+D6oejCUdWmv1ihzSmCBNHNqUe9wcSSyKhDbU2JEbbVoDrGCSE
anV1d8YYqvUNIlI8eM8Xi7ksk/cSvXAt4eLv/XO1rKlKTBnsQHgQjZZm2a7y8nXi
LEhq/FgMqkXVwVk11wpDcEa0VgQYVYfeNMP55lK+yiQ1cyQS1uuYQpPbH7I8JeOv
EZPaopkmnJbDa16JmvwWvmX/UlZSePmmR/xGOB7H0DIZTDKmSm42TSEa5GXANCfY
ZexJ3PjxK1iwqhZmukvttVC6VtxznUY0vveTMIVLigN3K4URujwh+vkiCGaSytRE
vTgMA5Nnt4Uo/D30C4fNzsiYkAR+SYb+SCFlhLgV3ikjzw+1nsdCrw2N3FLxbOPT
7zH10JYlQxSdWJ4i6SFgxn6R2REl1rynqegV2FAW3XMppwKhsf/YMQ+OJNbSHLjR
q6n5vW3tmPBNXRsbsQMVp88StuVfkwlO8VvG4ENGN6VFsV9C0BWI1BCmQ9arxGQy
0Wlk564oxPaIbRj51q1XSX3aMwxckgCnPSuNdQ0aiPEF2go9wCLS5pfd1sgoZD3o
vtS2PcouMMbKgoD7u+2G3QzlwjdYHLrfi7LujTAsMKF+ezC//qe50cNN1wcoHGlJ
sqCzT70SEaMUtmshvWu2ScxTyeSWqWBHWGuD2WoxnoR47c5pKH8i+iqvCEKEfljt
SmFag0UXzLqEEVlEuWF+PeCyD+EnvvTUG8LBv3+UWobLjactk4W21/4yZNCpRxsN
muIQi6nUsqTw1zPkmiX7okEb032iKKw8ytVFTASMvok80ZqgKbZJGyAQH0dIF08c
Txhq5POEEfvgtxO9jJecRL2qhDSZo8pzR3+O4Gj1jDs6CsLzUJU2pFx4gMxlco+u
k+nbDnG9+9Y8dHsLObHX1mJD8PQQIfkRLKy9q/uYDhOiL1V561fwB96k3ac8fBSK
9Z6TDgbveOGtgoxlbQcifP61wAXsJO37DU1h0gbWN3bcJQoUDBoVnZB7Di9jLYNB
CVslKE1Y7xQJHt2j9kQGz458P6GDBAPaLnR8I8mZLMFhv2VmsUEsYoj3C7ItJNyw
w1W3f2KehWkFTuryWcHyTtU7TlYsOgeVKZeMvx0mrmtjz8AppfusRc14ELzCv6Vr
kcEARFCZOl2zmbDEUiTq94kpv6isK6G7j5FoA+3ovhyLPhNu/HlYu0LoaSW8K1TI
rG7ijQkqMmYjAdpIgID5dduh6o6d0vFTXiuiRQ1jZ4l48l3hMG8k7ePgxX91wTmI
iG7mGnSgdl+hO+8BTa/Q9n04DBZfSx7P7HSNfYUIHc9StRywDjjf4FLbHXgERIvU
I3kvkH0vQp0fvVzRTaQh/hlDC4WU/NvXzC3UKWmDSkEJSF7ymHkMJa/Wy8SdpDkz
V41JNq2vcMshQQN+vsN/p2iCC9u4cPvaZd9IPv0z4IiBElRQmRJKqUtI9CE1SXxF
Pn84VmoxjnIlmBJrhSpNKuYdXhy12tgLSeRjiMqKbE42y7IEk4BvNZ3gwyNcnzQN
8jqf/Pe8Wfg8ZRU4/BLKXof7cAbk+XTESbjU33kP0gj8PPm7PIFJRbertkzt07mo
wIUF6MmEbxs7Ds/G+jWtBM2SVpDbqehaDdLKJiTOC7CIfH4BAmZf8Tub8MyV3y27
nxrzGkzc7KloxWpCE5gV6rTXHiYaPZu7zMD9/ACBA5fE/8MuiIHekp2Jw22iDKUn
BN4h7I+ZfvyVWKV4pHGv6SOzad/q9oTs95O73sfJXDpr3HjsfyP6fGHTE92lGxa0
WGlEqW6oqPXF/1yFKbw3iWJ/FjVAXHJLoLslyZsigu0JhI5btgyk45l4C7doDkpl
nu+rZfkdGQ2UVvJt7e5BR+WY23XUpdA5QKL//IlZq+Uzunx+dNA7U4ILSsolLV8N
byB48F1rmt4735oH9Vh5aZQ4SozuxNh37u0j+z2uJ88jLDrfGfpFi7W8Agcu3VvH
+w//qKnheHtQZW2BBtZ/lOuUVKPJcoo8HxEtM2Gdn80P7ETIEPmyOX5LrGLj2jwJ
VKkdRPz36GQU+wc5juKa9DiHRRW1zwFT9y4jmUuolG+M9JJ/QPz/qg/h0twAPAZK
g7S1p23wWiT83bbSEDZ/k5oRDN5Aop3HDhOq2zWQ+lzschZ0HgTlyT/5M+WdBb5S
uOBSm+JF2mCac4BCUHtoE88EEKgch5yNL4J35X+6jcGcI0qN4s388xmD4JTQ2gYf
sUPq+tKgnPJXr5Rl6uxiMBtQFjqFB6stl/+t5ww3yX/8XQaKCmHG1lfS2xrlopMK
O6iic1xGld7y1BE7MoRU5NMSLz6d0X3fIQAMt+FujTDvB1G4waVt8QrpRuTTYSem
aXXYATRDAPdHQUfY1POVw4m9pQg6c1BqU1JxNAebPyksXfkKzM8nKs2kXU+MjPlv
nCpVWWTWdOPl8WYsW3k69MzkBbmyb9SriXftIFqx31PqMgW8lIM1mPzlJ8dBPCQf
KXokdDY9Qrh8MlXNC7YQaDp/4De44rZa/HOWkBmLR3vIL99Z859ENQFOXupz6K2B
OiZQOc6MO7rvTPlCaNVbywnwKcbymBjXqZ8+3rikG5/tR1iWHw4r8dFEECroWJV8
ogkWtJMHLvqGoEYB+4/8DdfM1Lfx937teT0tORMLx0actQLfDax3OXDOoyjHt8Vp
Q5Ms580Ow2uRdQxSLT8P0J7jMfBIddLFZZP+cEX9GaJH33Jm1dxviMl6Fe7vbVJj
Sm4DpunEomx5focyOMaJ4N0SwusEKf+orDVdA9sxpJpfO51YhuQVGaZIpSkDjUqU
lhOxOlwDJ8OwmYXTDDPX4z+Hq8vaaoJaThfkBZDX9O/05QPUqvxCQl0bcjfhnfJP
rTAevr6xiV/5BCQlzlksFciX7Zj37rXCdbtirRt8LKP3C41oNUEfrG5gTlMq+9Az
WxVkGhfzzbaFNj/2y71+AkJoSHb9ZvLc4c6lCyi9X2GuNLLCDjXpKf3iGotVcL4a
I05QX8B8byL2TBn7v7cMulWgmGwkrL7N8VLB150XhBFNatwXDxKyhARvyvGG3rBs
3U6sQSfrzKOw4h65eETjM7CE3qrdOTibM/rrYJhcWaUE8LvYbJ5PuHSM+GpC5Jyp
o+cc3gJuTLdthkPLWOW8ntcNYBW+TcoSb+/W71YRx1kK78J9H33kn9gkH9/DI+NU
sU/cuhGDV2dbqnBLaL0g2sZHzVzbLOjzzGfigyKuQCHAlkrra9zzpnV5YkVKsIA8
vkGcrKZLcdg9cgyrUSFfbBhS2drKyqdARrbkixQPijcuYZVFMTy6JLUL9t1BWYnJ
70HYTH2R8h6YB6TWZSTdnaV+KaXxjzzC5KaRw+wWsyzCTw337C7TYvaZGPOW95qU
InsVXwstWf0w7b51aSpheAw03Qh7BFKq2hWgm4yIV/av2iEoPlU6rce0Znx1J5vz
D8CuorZfFC8SNy5BdBY25zMeb3qEC9jbrylVl4xJbkAgR9KX36LmcP/w/kNrPmHr
Hr5ZDp09gvteGAbixCDIL7U6hn/ZajXnf9yHkBf9bI+/BrXhPMhVvb+lVRWNI6zc
scueLheUvVMdQcZ4c8V58kcP6NCZcnjONPRNAtT0K6luMDhqptar9DazwRmMeaq7
IJYyQ9GUfJsLrnFWRz0l8HuRSu4P3ZQx/Y2G2J0iZ4r0fjoXa4/Od2OfAvj4AS/W
cjTPlSYy/kcv4k9L9vwyHMACriYTrv85wI4GcrtE0Bsx58jlQlICXlnToyEtO+/2
/cCFP+ydRXpF1OMkn5rsy3AaEYB3xUT+nrpIIOdmF3wCH1xtQwzWb0OMrRf3TbrG
Kdu62oLzXly2Z9UHw8YKiHliyteB6yxrFe4n9mJ5kFoE5cMSTKPWJGXWDMLksd9A
JtVK8SY8s9/7GU44Js5yLuOKBIwdrT+vHPOTkGM0wA1AtifkRiDpGLHbvr0sKVGp
MhpbNXEuIWMZA4uiGF1TM5c6vIqVlcHhTQGuIa5Shk7tGMlhSDJPOUcKzpClo00v
rtaBCWua2FcY8lBaz4EgzKDQm6LnCfkakKtXpnXaIPZqFjAUodmL0k3hI1TlC4Vo
JCcD7MB0xAI5zvbnGfWg1A/oEJI3u4M2mbMdp0+FRdT34VCLdNfDJzeN3F5PqjKP
IAS6mdvw0tyP165lM/u1w03oFoM3pNjfJOUDfMEK2778aFcd87ZJHbEA3B1PYIIw
uZS5uOIL/6p6lLEytn/8uarTiMNhh9RwT2UZeFyIU0rli2G/7IxWILfvx+fYWkCT
vrqkf6wFtVXt6+es7jOzxfQcGXvtrVtml/r99aqyvZuSzhXa1v8vP+3vJUskBzD1
8YSvEOAEPFP8IF7IWMnoA7gZUiogrsawXVrAwzMcd+JTcjKRHWFXZg/WofIOwCOr
sx/7kTBDidGUkohdRUfkEQYXNgrQz7tTsB8+gE5lXpYYLX59W0ERSF6ryY+CWD0W
jZUJT3OFjZEJAZCz/PjGLZus6KRZB16eejWT1ezWGKu9vfkXZyEvI0LKHgl3pQ38
2hCvOT7P3iAJePLYP20UWRNFV+ec4hdGua2gJd8jYeUfTcQjpDgUvxyfz6E39Kkd
tK1W1BU/vvL1UGwjxi/hH3IM7wC7wtsnWgfVNVEBRuEEbiUMihCbUW1h0an0UpnY
dJ9jJmlGp0ldt2SMhtv213pQfwoDvwGk1TyzKPTZZjGRcG1IbfpmxkCacvRZo2X2
v6WpT8/zpXi0s52cE551Uh8uXhBdyEMs8aVeHs0gTPRIR/KTO9JGo0+eTGwQcyI/
xbAMPHlsm+1mC5I0mqKpvRa4oht6lnbon9C0XVyvWVLLUWgdA9uUuftHWidu6sl6
xKtM2ri5vcBXZC3yXqSd9+9MWk0r2VJdoE/8XLUeG1WigvySG5tyjOwN+OepLdBb
Oi0CMYNoWmQ/C90Zgh3Ng3tvdBsh/Sz++mCAPefDHnfWAa8iWJeVZ0o8wso7fwVP
8BXBrRsUADWeMmFgbENUb/ycB2Zpz7UH7T3CQ9tUv0jEjA+3p9/F1/ncJmP5eucj
TWfiUOCETgwmMEcEkXsIqq2cI/qJn05lM3KW0CSvS4NxovVwYCLjrdX6RXtTzu8H
pkGqxJ+Av/hPLtpFco5LN1p3D+BOP0JVXdpnHz9iUS8LRhMd3wA02ccPHIyeGcFK
Lkcuh2OvqqX5PG04dAUf++d9pVlT053sXnrEH2wWsYndJn21HY3kpdWHsk404QZV
oA0BPTtE91eJKgptPNoCnXObWGEWPE+ZSgjA1Z1S6BMB3Ia3ii2D0AtWl68IxH+H
qKUzhIpCezD0is8usSmXR5YwqnrT4+SFBqbsgjp9dWKNi6jFsfmNeDkGFyVuVVmX
SGyRYGzw2F8eBEfhoOiZhhSNT9b9+g2pmVA5KpPpK/XiwaMYLx1SPtfUhqFJEWVa
wTTWbPJ9KMwDJybriBbi1gqbjQxlOkoy0sP4DebXPW6dV7rb60x/cSYSD1wQvMCv
18da2skWod5GlK9W9AuXSpBhYmvLES3Ifmc8ivN0I5MZD4gfbW4f48/mLjishgNy
XcwD2suW+74N2daZNVpOiW0egygMavS+YV0lfCTRB5O8H9lzVGUVb6OXwThCHK6W
7uoIUxiY95jl1SbZi4QWITX661veuarHGTvxuJHwstMqYy591viaomqzXDD6alkj
U/i+Gzc+3JHg3DeozugkxvYtS/9glyr+RE4P8yBDDCZeKBOclvVpK9rf3D1943ti
GQqdaNMt6u3VfN++3lzyKuJcCIQ1nDo0a4iKm3rIAwq/5FIgvLfZy0aOevx3qerS
sBfLF1g9wgBOf+vtv400uewPNKYxXTcoJs4An+DaFF5tkQ2If9uWlMjiSIrVgyTM
FETKDcxSH69Vk8Qi3qdkWLpcEu6bMbPlpKfkbmDpoBgP8H5Lw0IJL96pBBl9OJ3k
6N8n0/5zUpwS8MYUjxa8d35rEefsmckKIqQiOk0YhA76h2WFfsGO9rgYCuHNUxaV
7qsy3XTUWG9rT6fol6LzOFnY3FsWrBX9l0fmnI4Bu9m7rmL/7O6DJjLDQ+xfd9ha
jWM5hwU9kvxbdLRpgRD24fT+mV94ieqOkRLQNMEkkPSXyabRkSXMr8rUJIZWytAU
uIJ6gSLKv0sFRPSAcjaFgTqg/Rp/lUdkLg5ikbaBR9IIrs8zufIRIi0P47ue1Sbd
Ka02q/C7frUZU0sUJz+jFdn7ZAdmCFrTBAwvOjnX3+Fdl2OE3eGEz7bPxygNdjjR
ANmIcnlmNmYKSvg9UVEvEMbSyLKXIfaXNvAVYTmPcFrLjbjBgb7xghW4Da0b/Hod
ZOmVI0C7c3qJ0ii9qXxIUjNJR2jD+4hEjFoPqOr3gsXoulYxnHbR+FGX8iLjEy6r
JewpVBjdR9gcIf6Th9LCgmGkEnuWQRKSuYdS/A8ykTHclHmXHjyySTqmcqx2u3SR
aLz72E/tGEzDnBKjbfqekyR3INoqlY4uoUHe8yfqwu21jtlz0/8ARAV0BH1g6EbI
6T4dc+ZByPW9fhWdtmlxXW4CtKnfDseZXUBcOhenmFSdOGL/pZ4TwMihJKU7oanN
0ibZb1f59WyNFAZCkLxXTch7c6RNQknmz0Dm+knibRun3Z0D8xBvl3OzoGNuXz7w
jVu5326KgBhEf2rg4j/9UnK3ZjU31JaDVZqdUeFnmiMI4Zy+CNuhyqE+ia8mXPj0
vxWZ9ojlPffkxmC2l5tIS6aDrY+PFTrzF9CBn3pVVi02IpKIvaF2Bdf5MRAJIu1+
iMGXUnUGTViWwnt2C3GIrN24GJpWwsVFG38JAjTjD5onWNpS0FudP1vRtACNfzas
w5/srNCfH5OoQTYlaXsuECljNKV6L+FuQ8spIeyzqVRZOnDuHRb7yKAAiOOEWaeQ
9XAn5scgg3D4BNZIbzutSbUYOpKB9pLybbUc4HHLRb6tLrwjw9DbEGbVNgP8MKaz
NBLwjyefDhxrh62oEexSwDNv/kHVHiSFniriS5+JncRtEBF00qR+9mOCb/6LcK0p
SfoI7DFsBW4TVpWIgWD5kONZALW4JYti0cRtViZZnLW2cvVOHMrEAHFynI7LT7bp
CMtdDt6lfSvxpuUXGLjo81hAcFdYGrdF/5n97EtW+0ebUsQixusI4sipjwJ3vTGj
ByCp2onSbiL+GjJEM61Zv8dU7SUhF9UXMkF+/BlF4gb2rHzXem1XPDjs8FQLp+6d
i7adJl6Dc1/K3mZUhHrI7tN5EMOzJvkP77Ie3KVYZR8NYbkp6r7Af6iVYsrZvNDJ
PwhdT+EXsAP59lzIf4P0SvVCingKos4oPhFnUUMRFuNmRd1CLuBR3rUCZBmOCft7
mjqEwFbQnXHxRMco7v7ZSdaNEwLNWJ0EFZdF+9b4Z7YwWq2CJ7vt7HCcA6WzciLh
n4oNWrHRPNtUa2S9QdGsuzsDVFrSfc+/ntqWQQXmsWpqAFL6AZVb0oV/teWwLVGm
4H5kqVzZajXKI5tHxXigJeie0InpR35+UJpGtGFoPFLdJrUoro5vgAIHPHCNethP
JEgdvNbOBW17ycfziAJZcz5RKDvunS2k33MhmuAf/Hcx+Rv4QE2aKsVbnK987V8t
BnIEuazeWf4aKrY9/z48mhDrTC23lStQId5HmnDFl51YNuh7/WfTTkTplcYCfojh
HmeSla5WEChuvJh+IxgwWYVy+GMx6H948NCTH5XDx/lz8ZK/EhK4fL7jseWw3Ahn
sCZqzo/t6e38NbwBvpsX8HzepBsaFIxGprzoRXbfDbnY7ZGDmW+Jfea5gtLJN9VG
RSTcBUp4JNcU4hvnWDMeqUsHsWwnNRn5G3S2czZS+2omaE/yqWFMTlubFfz1DQx2
c6o2bOAvauBA0fS5i+nmEdiJOBiYyCp2tayF7KIysS8WLMCCH6H9PNSC6bWNucTE
Dj0xkVe48FybTtEBUxSJoMLeK0evCWmVaf+r9hujzWIrXrb1E2mg7Yr0W6/Sh8zw
q2laCFpiZYJkN0+Gg+AvyINLqvRCAxN+IChd8eFfikb3QcVdO4JoenmZC3z/fTsP
REXGyPkcxnoBP9bM4pWaqeGnKihVCc31gsLwKeAvRcKbUTZhgsqvjXhuvMJth7p3
C4B4iBd/HkVsBVQgcwrmHZkBOip6spDbXXJXKchuPUfFrC/lElRcdyFaCSiRqDM3
YrlFt0eownrrdHZQq78LnNU/OLUmWPT+pjSQZddR8mlf8b6t/dmOO/4a6qDL0tbd
TwOuTRdZyJxR6hmqciFM3VIg7B3TthFxO/aNFLPdS6bs83AaIqPbQtnB+kj0ArV6
Te4Um/tpeUXiFYbO0w6zJASVYdbXk0HV1/O+Id+uGZcu8gBk00kRNWo1+HOhFDMq
v4UM10oEy8a8VA9caQv/IeSZfYWSvsapQXhL22OW/BV1neUx9biCK9XnUxObJowR
1WbD/DuYrYCtJV+ngzWyaCjXC/MAQW9AZ4vt3P0YIqEKdcqw6pshro5+LFj6mUCa
gQGhJNAnJH3Oium6aFYdNZdkdb5ZMpTPk+m84dTJtaJO3y+yuB/EMJRP9YxeqZZ8
y3ZlmUKiG8hjVa6wdq1TsQ2XdgKnpCS/graryKT859yPyW44rwoPj1qJB5ckt/Iv
qAPSGAQXLDZ4EgOiJPz0CPG1Ajo6kwhnYNilJbLlYoxje6yV2t9w/EBB5RJ5LwuG
87S6q1k2O1w6mFi6O6GyZkVCmiOITFL9XJZjUF98M1/VwwY8EjMLMoB8opVazpAQ
Z7neoH6SMGy50PI6CixhCeLUkf0DmgUp86ri7bWBOq9wwgoonts3LpPXZ+8QRihU
zBB0KU0HQkrpRiAKiOKwsWP3xZKMQxWuMmtFWs5AC6JoMk+Q1oYsXFeQXVSG9c1l
QNwMRT1DoGChkvrLSxojpWFk6LXjpd7XGmhxdQFwi0KuVBfC6vNQO5rhogHP7wvE
N/GvuViDmOJjCwjbsKhReLEl9BZNdhY7Np1YDX65w/0lbBnHSNc8CgFlsLyDgN44
g1zOkhtwQfhJ8M/6h54gIz9JpDoxiqMeQ6GfRiQ21penmHssix43v3aCgh/LvFb/
NwWe6Q3Rb+nySqziOkawUwLDcj10Kej/D56SE7C7w7ineTLmLmcClU1FW9zXb9WY
nT1BIvHS5mkKVq0sC10WaRaRMqoDoWdnt3/m90H4V/98h6bKyQBChuXASvA+m8IR
5oYiENB0dve0fGKvkAt7nTfV9Lkerj6mgAm/Km82h5Jij6W3hTndsf16MrY6DgM9
gesyXBnZ2x+C7cTBfM+isOaP9wTsI7VaKJeMcFea5f2e6XPGI0/KYzN6su+/kklK
dK9qrs+VaqaFIUUgpWoGVemR4/E2OyfjUTb09D4TfMzpkrzE7Iz3fusm4fVE/uFq
XSlO7blZHKBu4dKnuzVkWUBmqUzrb2NZZkh4fWR/T4NDxIEtu9MFgwBXVAJQPdjg
/DdQLiRQNy4Q6R1CkHj05ULuyQEb3cwiB4GVESWwrnSdXpf/IXFZemPHpvQQsji+
AIKsMFLpkHlgPYZ6rSQYTlRr0WiuLx8Y/jzf3ke2TqcSN9f+GOk7TV660WzlCDpr
YuEUlnyQo0ubHcMSBkJzd2rXWyK07qL05uweolMGl8XUPuwE79SoPWGjDWeMsfUY
mvMfeoM+/6j1If+Qvgk8DM/uCOTfGNwkplp85CQiohutVSPbtkzd2ln7BCmwugD6
i3xL4qVVCj+3AcQAA/tarOY3mi/9MHREfgBH4zFpx87PHCuNVfjqLy2guYBe09SF
kqLTBdS41H8BYEte4jyAUcf8fxa0tYaHAZ/1a2ViScQBzGkriyllaj0rku5uCXgm
JxnNoO8l7zDUj2Vd+s32AH9CzEVbyXXrDUbb5g8IaS1eFAwwrRJ3vwRzDUS+6Iah
pi646kss+jevCb4Uat9Hr8Go0WQ425TdsyKHoDOIa8g1zgKh7u8IKRG+zZjpwd6V
V+IuMilAG/lHsfOYeDweMGJDBFaxuqvtW5VH31Z7KPjRyYyQ65zBSMyJUQ2UYQER
e8hbZE5hg331Sm8Qzf2rNIjoXvl265YiuP170Dpa0DwQKuJxcaZ+UKzQBKVrnrMz
QPoKYPILcOlpWAALPJNQxw1yg+Ll5GymRLK2RbgkUiZQypwH81ceb6K5ol5EmSYx
f5BRaRLP5uOSdwqsbpn/ivbpoMy7ueerRG1x5rggHo8GW+boMmJHUAqui/dC5g8q
JBN9PMghfNrAXkOQMdBWg6Y/jDgm/vXjHGK4mUMwNivCc6D7I1NwBnwpTdou1UZp
VCPSsBLfOIyYPGsK5JejeE+2kmhwxSfsap0zSH1qV+/F7DB5cfh3s4zEYkqPhhXm
jd4dILACYpp5iO2A5FL8KKeiLTfqmhqmL7OPMRFav5bnfxA0j7zxbDvQw5V42mTx
xyjU6iqYGDl4B+8xIb4ovpsWeV/L7f5OrdyDfhXYc5K9MgIFj06f6tjtzxEMzmeT
WRtWHNsmhdLZiF+hKOM4aZxc24iaMAaUdjhKyU2gAtRFDqa0dsrFq31lswyP+UJR
t+aIAnQSZMRW8wk+TShwFN82U3qxBtUWKGmrHY8kWjG4u+DW00a5z/Z9roJlergH
7is1I0yxe29xBhRXqiMOFosJZCa2ns3pron4Jlbz9IrsgLRlRdeI47ZPj5x4u18g
PoW2eaVu1VlNVEyUZ1dACmADCU0pP11za0/Pk2O6Wtoan9z2LIHwkkSP1pSRxHNi
WQkomMvPRFYTuIWRtxmNQwpHIO45qwpLUmqh+HVS0HND4UU+XGAbVKzAa/CVjoch
qL6vKr8i14zE3uuE1XUTlE4rHs4aBTIZMFGTkA/78IJzcNmyDuydwTbo5ZkIGZgD
AycvnNHW5UnOHKI+gQCswxM5fnYLRi9ynG3RS7O69vYnKB9OCR+DWrsEzD/l4TqX
AeDA6rXsEi5Tml0SZkJ+8B5OSeZHMYZFl+G2OHi9MrBhS2MtEMVUFLfYFs584G7R
mdZlw59hyqK7sNSMBalOwOZK++FaAN8klJZCD2+2m3dYCvP2ZOOm7mVuma0dKDiO
Afkae/iJQP0PcQzOoAJJdaGekjn8Vp9qf1NP8H3v1M/fcH0ZVjLFtmKotjKw+pms
QjRBSXHKyIxatlIsDGRmOdNQACuAEk88IFxog1rVa8ueRnBKCrXxQIOvCnebaOEk
5vHwXf4HnrnqvbBlDymU4ErOSmrIf7Zk4eWO5H2xqIpfBBaaDbxI4kFWC8XPfjdR
K19XY3oJ0IJ6H5eg1Wf5D4kLyLOvvYSBaF9NtYudewcpY+7yUz/TEL5mlyZla5Hr
7DdiD3Q0Y4xpQBrUOfTxRFg4X2G3PmzfC0Ml40udtCaPzDW3OmsR6QvBfamhhvqD
lbpYjJHGRmwJMcJsIeVOiRxG0pruCO/NNHChUVLnOSpvhA3IXl+bZubfnsCkmc7F
IdDxp4sI6surC1N2v6Ar/HHKQaYRTJ1yRWLVaf9/oYo4uSD/CD15b+xrwVIva1t6
25hINVIyQLuIyHSc7MkoSobrdUsjvOfRdS1CtgVYkYeUetaFLJ9fYLvrtv30xUEE
IkAz8gs32+yTXVt+eyOCbkBsG4XM2HAsy5lCEWSXiG6L+dsDeRGR8QWw6C3/p3AE
YhN0QsbY6VJKmadoDLmasPcblTMxbu8MwBlc1Ps465XHzrqG2G1C/cK2YQuuHT27
72PDJH2VB3Kf0ccG2hA9JDEJpUHi8dlSe/G6+QbE03fURjaGVgx8gv2JNILlRr5l
C8/JSJbD962/1wkdddBYRbCuX+iS20nrKqHxIZOSd43tXK412jxylCemp62g8Q0D
JNitZh5TFKlzDqUcN7eutUYk3MNZNFff1y7Zyxx6CsPiy+G3scNQqPsvxYbcBMea
gmOjMrmpXc+mQAz6lHOyYnN3mTeMdtBhBN5quPtWM7i7caIpdasYv8BVB9Wn+0hl
qBMY+3VlR51VXdfxd8cDEVHsi3A4MfSjermrTu/f+ojkyRXxKH9p1GXN6TF55CgC
DcVvmWMb5/H9q7bHdVT1cpsmh6Jx3qV4/q2Sj/h9ylN0vJ3l3J7Eho7QDSj5JrG3
P9P396tn81UE07+QBNpmeyGL0ZMBqEUrEC9RmiOeBeogr4sjFlwGs1FupVvSVKj5
rF3LbdEkGlH+W6QPVlAROHA77YBTuiqqPmFwq83F7zXEWksTY3VVQhzBgA2pVxnF
HQZzzAdN+x6Mo18tbStzrh5gvVM2Sf3FuVNArLPAX7TvvGnd8cL1sU5PvD7vikJj
vZsL4Iyir9PfKY+llUhUPcyY2i8Fiykdf2N/AsWZ3g4A0UKXeIfapfAOj+ZSkWRS
Lps083Gk6n9i6CKWygzx579/yUB7/AszqoAz6jwZsU5u1yjmbTbAyEubmTLXybus
55UM4PnpxeHFFyYLkAYpTl4MO1x7GV44o8hWEFRdATH7PStOv5gKFvthBObUSeT4
OKYC0Gr9C5zwunwNeBLl7ENkfqnd8wI+X8nzsL1LYRJFPwoTUhBdIoTxodA0TfiT
KwKk7p/UkOEpoyjAUld/0GKVYXxgZVLGi7DAffloQcr62BuL+WQB9/RHtCEEoVP0
7z/IdPkrHOpW7o1QiMKBy+3CQODZ5oyKrIv33nDDMwIjQ2ujE1f1vehelIklYJ8V
GXkLKB+VFG1iZyfZU9hMt2KnIQzsQHfklcQ2mWPTyWhWR/frs9+w6WEETfbHG0fZ
J/bfUrYraAgSEc9VEWDwWgUhpWY42hVhMsnzLzQV7WjelME+NDWoEdQ4Oq2oSn1A
huAwuySVHBOPRPA8P9fsZ22u0ClZrQVU0Wjg9H0M6bxPyNrz4n9HEBCn631wM+uy
T7qhSF611GPdepMECXHJ61f8YN9Vh5Eet7GPHT9l3wOZO0mjUFNXg+siCkS14f+i
Wjldr5PhOzRoDaoOg8eTO7dxkzppSl3uo6woWzcN8i9Rt/ajEyUQOcvSpTFwyO9U
Xj2hqmLl6+PFA0o4snPaVqNNWZXHaNfik4ajcwO9JJ+8aE/GeZQm+yDQ3KSDB+sE
0X90FB9XLOWvjmhKMv/8+SxJUPzxa+UaaFFey37ouVeI6sr76+aHG7PgKMd5qMFs
WGWasUPk0Gw9veGO2I/JsTPALpBKTETcJZMquI1KvkXYQV/qn54x5P7gYt60T92k
6ADZJBvUNPgLMoHuTEbbgOylIVps4r0a9hZxL7EF6FjqbZA7Mix5D6LOJGnyf1T9
2m3t9eA59FdR0HZqH2phLHxihd2qMVUSVXaMC9BX6PsNtPgHWrtt3D72VafMeKaq
U3ajdaev5lPmIbxTd1QAZ9yTeXKH/NvnsVH517tu3CEB924lKUztuz74XWvsijIW
rl6EnF0wy2/AgSPLlrZjfukaIYWqdv4C8C4Kg0XrlDvxkMtZXDN+w+NgRAucrxDY
BI+FM8w7K7NXpLFG5FR9SHH7PKlEhm713cNdt2XsEPMU7XGZNoOKE10hUXIj1T8B
hoUIp07f6vsvt2u6xFiHnFaAizQwdriM/bQ/Wm9H5Vfrzg9S7DaeZwrsJ2MhZ10Y
fi8LQ/7EjgMeqNn/ncRdx2zAaBkdncJSigxo0oGdC1fqpv4evv+MbShd1Y756gCn
t5vB4duJE/r46sGV8fjyQfu1O65OOMpciQWuMc/B49jHbx3ZxtF3UEm4L9rpiTnp
ZAnvbPTn2B1u+lstkTsZxoH9JcBq743AbbnljFLgCSyg3VGWwrKl9cg2mu9OWgyh
UnjMHm9n3Z5zKWQyi/rKtFsRq5AfVuIn1FAqK3zF461zhGXMP2BmB4urmVh/maKh
3rNVVQWY8yz8NmugdVTwiGkTaw1J8b0D+ppU6/NNiupaEbiE7Pnce2PVQV3c0yqf
d2EuJYW98zC6C5O+gwo+j04FqaDZ7EpybQtyxtCNMvQpXXqiU9ok4Ks8Eg0o7a50
6JkvbLorQSPmygW9tLx1Zs/lAZd/reRlvv4BrdwZB/XP9LM4hHI8L7O23e8zVg7V
e4duqDdOAAylQbBjlmf3HnslEfL2heyg6g9/4XlQRVIn71DYAkFsBRLSBjSvsDk3
wqkPlIyPv64s35mJtk0dcHpg9SxHBJQUIL/LxI73sy9dPnMdjnuvUYbitSUrAYfn
omatHcl1Bew3U949QfrCUb/cBkT1q+be619AaGMsW4hf/8Y7D9RAtBycffFTFU8t
iNFRbyTrA7o7JA0+fuqFlwWiviGTMm63N6rlUHjwoeIFdjZ0GqxpBILEMfw1nor8
FyAqybszKoQ/q82PFDKmDPJ3pchL+VL05DPRKmpVROryP7CcFQfpbBLceMolR81S
VrCplzEBCM76gu9WOCDWUjo4j/Ru2CUHJZSHtJiq8qkgLCRsddfGYExlaYtNUiRY
Ylq589PS8lUIrbX4Qm/LkbAOR4ko2RFMvAFba6rBYngQPya8jQSS0q/un5TC6+SW
ViqUJwYpJSM6AXIPvXWSwQMfzYk3GmzLtcU/f17P+k5Aias5yx7EpFomTQZdezGD
szmw0hP4UbDEeJhUb5r/EY51LeY1l0TT+4d57Q0K34e5pSdilq6yGY28o7Nh5kpL
Qv9hfSgL0NuclcLC9q8g3PJsoHSGkF0LlA0z9FBVGp3UvayJQhrJy6+PMZ0xxmP7
PxBXp87I2oSYc05qc3Wbyn9RIz0S1LS2MiSgEXm4mlB/4Ji5IU7euREg14bUF+15
Uf7OFPxObfq7HWNWqQMvVrS9Gyjb3MgnGnUMdMcYqR9H4PkiIqMXvgFuQLe4AJT2
QuWQEB2t462diWpJpCil9ydY/cCTIYHxr05RpeVVXHo5/+DzC2p2gcJo/Z6KqzI1
Ll+6I5N2PSMRPJGWrbDM7IulGsy4JgiKUi6H8vVCqWliCkfpu8sp+m8xuTS2D4Xm
PViw4efXyRFVQ6lP/jAjuCL02bwzeRrh+EvgnnwFGXPMXCegeSV21FjpwDDL/F+9
F247AzdxkSwrOIYze3M3xBKdc3LiXBt9W3Ahw6KswcoCQjCsWREPnux/1lW2oobg
Cz8z/7AGgpd3B6hMRqcGIiYEEtgzbwzi73OG272dpK8l3GIH9BfoT/UtLHBcUyVD
yoXQMxKV+A6hED84QCQ3RZeV54LidiDC9+3l36HPbTksRJox5PH9BuLvv5O7C/gA
XtHphVbIH7O+DbIbicLdyQjH2IpYHekm0vdq58xQ3uIiR2tFMTfBhRVSPd3R6pst
eEU9JDoxrymv/mfGekF+buMRiaDqLFMIfWxu2ALtxgQYLujSzv8ZX93Btat4idG/
t/YXuq/kAI7aO86itb+681IwU2dmwKE36knarsQ8Ci2qeHyFBITYckd4hBaSzwQw
W7fcolUmcJO65szQwp3mmOqaWC4ReY0Bl7OLmjT7eNZr4erApC9XuhzlCGH3f4m6
y20fgGfSbaTVv7v1LV1KL9d/Ou9M47fr2wbGDgXBsT6SIpiD1U0RCgg1/xRMc+hZ
u5YmG63KvSePGE04kCx/h4TAAO+UvAtzzYXCyxM+SkHZE86vPopUbpHYH1qSYYkX
BH7zy2S7w9aIRB4BPjThJFY+k/pdoO4x29Rq/wigPtMHwfaEZHlzBd/m3odNnuAR
18j6UAppE20Z4k3zF1+4KUeYC9uyUA7Ni616i84M1LxfRIE18wsGW4y0mMUGTjEv
+TU9s1kR1PKJ0bSPPHOp5A1NfbTuWc+nblPBHXW4PqNKfhYaeecKCnaJrW1nJSlg
JMydni8puwmySJf9rEC89n4xJbEZ9zN7U+x0gIKfB49Yx38ZDy1yz4MFw1NJuGXj
ZXbg5vyAF19tzoMvFobr8fhGCjT2h9pmI30KnlHS1CUM1IdTK+UJUJyXJcexGX6i
aR6medFDWhE/r5+Mc6n5lVlxWfUD20hp4vnByygTX8dgeidUAR4Ff4gnjS35tPvp
99opaY7gxtyjEKEhuPsSQXwII6TD5HejFp76xpNIuZ2bxLixhnYrdpeEpeYLSXmf
eg5UONiAJcGq96N5iHO56FL8UL/KGNVNuMFOOtpTYp7XD2XK08IW+Iv65kkOJ+u4
wZtosRm8XeavPwGN890++qCT9sNtlSdx6NiaI6ihmKx9wqYDrWXhGme3y6TZ6ou9
Q5nzL2j1k09fnnVmkfZ+EtowbhthpdTI9p6uZtG1kjp+CXiVr+ehGN9gUJXgunsp
ySCmXQ2SvyNVctAJKw1JPT9xrhk4d2WryQ4YDfZETb5xer0LcmpFsugQPNjIkYIr
9/qBzQaMrsnwO5ifP1dvr64FxpfqXEwh4he1WZ8X9s56gKNcmeDOPZPHoPjpoHIC
YH5EXOJ8nxizQKToK0/yiNkl5ktw+w3j8JRCid4i6g86OlDvush+hlDwio3wR+JD
NFkFFmfS+BhmWwOLBM5JUgETcnUG7XWupHVMLww5nm7a7/o+9iTr6dkRRzXcy0BL
gUmig1dqBK6YZnegYV0k4cqG+Oq7n2wkRFhU7dSnENx/H+3fhBUf6AQQSy5wzjin
vP1UrOvms+hs4nZfF7MDQTBYmogD69j5xItnZS19hDijE7OlFbkGxY1OuSZA5kJZ
MnXmzcKFtJKwwozrSMQeOIxrIqqzYbMeECsOhpGwouVEwq4WAJ49A1g3OA8XQclA
mPX2H/VcMO8D6KpX3pI+ZJ9NZ6cH+i9i8TYDeSxSV++VpahfL7+Mtswzs/d931tI
gcsMWTkt+6SAsk2WL6hzJ+LdrTIlz7TsnVC6xhwvLARIuiXbRO/69hhLCgo9dfgD
pk28To39FtGijrI/S1ICYqoo680jR0clg3Hi9h6TKETntol+joc+QhvM65q97ADl
Hxvzq76KRuztaOrsNsvg3Q9TscbmByT/WMsrWQ+UxY8afkqNSDGw0K5jJKdBYDcV
kSt4LXGNKUWN8+yWTlFdYQU3tRuEYaR2k6L+PgtKMjsF9RYSYK3uMV2x4WoMtEk9
tPgABJV+wwh1wREVWf8MsW7VIVgzfyGYLOrjX/81k4hn6POt3OIgRnDk5w23gm7L
cQu74mACbPq0CcjHfcoSmQ00ukhE5tCA4MvUBiWIvtBt6s1ikPPe3sGHwkHXNp2q
MIRPpRmajstmTjDP8A5vigxDlQMR6dy/IyzdYZgJ2S6cVjGeR5kVCdI9QYvZUb14
OWG/nmm4bNpTx+52igAFElKjzl2lvIl08/a57nW1FZVoAL/hXvbH1ssa5NKZCMw2
q/PGMHe7LeR0AgwnGpnM0guoFYrbruj1sR19g2TyZghyrtfzszYl6Y3gw5kBPrIE
Ng6qESZQBzYqEtv/nB8LPMh86z7kUIB4oNsvlhz91B9ZrCvnzD5/BKSQgkH+FKNm
4cIiL4UKJDdxrNrb4cCRha5GgIHvQ2V/0Wbl9dR49Qrjc3EWwuHezqHyB9JHQAru
gu/Sef0ohN2j1YunWLm4UpZxgAUf7aCiP3vXkzBg9Ubep+8RGhjZuxjl8eCC7bLm
jEgIRNerd9ayV9S83zcySNGe43nMtZat7CagEgRXYTYnyNXgAj+gH3BaxFPtYQ1H
3lPEuECO2eWEe22fVmOhnWsK1fpcuFmk8WyR6ZbVKuhSakVvymeGIZBvZKPLSK8o
LKXOITZnIVFUUHeFOOG+ysJLfuaSZVjtyUFAE/YZoE9dKMfI69wE5V644kOZugeZ
acmzpaTjsSkmg47S8X906/yJ8Q0O38hqvAStvBRV53u3WnVJQvHhbBJdSWj7BYhj
q1rVmB4ifah+yfShFZ0suI3S4p1q8tdA2LWjlAZBDbgAQlER8P6u1hVAnIJ4o3fD
B/fuzYonOmXtWaKKuXHdvEcsA7GHY2oCogXPNzpoKiGN0sIFvHBrm8ojK1eNoYG1
N9SoHmiwgSD+BaZcqdUwThKHpccmI8/laxxO9ndj08Dd5j9inTy4gLRzIpKp+Vxh
bEMGvHAsxez5B/0saRF7dW02kG9vZ3LYk0psaHyfY6oO+EsX8muDtE7cCd4hVNJi
xoFGm5bWI89YMks3x8XLrZcLxSpZkVMhRc23d4Pa6f82dUqcQy9gdnXcMSpWKeDh
ZeU2jsmbha7JIDPCl0C7XYonVubsGlTIBi42zIoRJCYVFPQazfttrLbZ4siH67Hd
5lstl7Nc5ylVUAtTUxfoFUSg/elw2wuNNq+laGg2KM4fToKQ8zw3JUW0Z/RYkgTl
yqr5t63N+RpXqEWwc5Zi4B0C3rQIQUC8/v5WU+7GLpcSfQNUwgBq9XB3vYgjNajg
FyZPsWCD5tcjPI2IJ41n+IutAXRjl54qADH1WKb7kr9HO6nCrfKJZwddlhqINNqr
E/QVvCpSRGer5GBBZJhecu8kGqngPpwUpDJ5Dd25zMVzDPLmf+Glny0yxLICYDYG
r1IWOWo1T8UT3IZw97wKhi/Qo63HYEyE5ZMYNLZo8z1OVYCchIqR12MePUX40Fc7
AlCZ3aKhGDl+E2oWdsnK8AAud92BzhD4fD1As3dhWSnIYZykoUG92zHfHkrYn6Du
0y0tCYVzEw1EDVlmL0xJT23pwmoNdo08OFg8pavzRgdgba0GACZ35SrZF/QwGtTi
ODoH9JOclkyRyaxtbPDt2/v44ajtnjRrUEUqSrnPm/CLMTPlzzzECt9i9GuihKbh
BtdCNTWbOlp0IAqsRXoHL/FPF5sgzBV6LJKLc8m5D+bA509L2hjnXVPQStYb1BgW
svLOckpGseToelp1DZurVjf86Y5qf7J4NQC4ywTn/fX9UHGArwxZkkjNIhquczLh
/gabcx8hIYZiFQcBymqSGtjEFdeVo+aDL0n///U8A5SVLxLPKhu5XuQ59R5j04xL
CbAEtRj+aCzH89mIE1hbh0lMLGZbL6XKOfqUv/WBtwOk3yFmPXSSNksHHopaqonp
e6pNffq6oLqCIn16YDbLhCO0cKGJ0pzzkn5zITtARdSostvHYfO9qGKG2/W4Ekey
Meml4fOAT6HbpxbGaUCtrRTPat2gnIyVaOdi2WiaoHbudWN3E6Y/LbLI8sPsziz1
7zi6Lurk7KVHkgtOtIerupYtSybAq+l8I+ovnkHosaCVEHN/cURVSfyCKry80ZMe
3HgkmqdL9tVjSxFfx3Rk7LOh3gMYiA5KBW59Yo2LhXtg1bhQW63POAnlAA9J16QA
L3vm5o6+1d2f7Sm97N1YYv7wwRafdiba00m4MOBtL2LecE1viqC7tDdyp9eMa7Ho
vFqu78cSqd+T8FPfUhhnQ5UJ88Co37w78SGbLxP+l3Rc6hXGRlZ1R1fzTnzBBDaB
6CrDL3yyXoZ3S7FgU0CQWRf9JoltwWygB6zNh6n20zHFk+LjIgmAf2MTNdcY0lcd
9ZyFOcR9RtS8XptfkCKJQPrN0AMK/IfpBAuU/n4Zorv0DYk+80ua0nyX4HGZ9RSD
mUUcWIEOPXElvGGmMT9pLb65d2DITQnQ4rco3FIxB6P9OYUJ53VNm8FMLCct5N2r
8UxU3v7h1xldR1+nXDfqLnxovvh4djE6BvmBmKMxS/l1uNY3a/kmjX6SQsNo7qpw
cBwbKe9gT0hmVYQ5GlJL5ddnVnDTq/J1tk0yOAb22suwvfCQAvKJ3Yau16b4oTeX
Ic9JFpLbVT/7S+K0zXSOdcNX9T/dD52f/e2mF80Z0Qv4R/P11bDoZacNJjOoGTMU
t+Qx8UiunRzncZ/iUHUF92iA3aoj063i5j0WvSg54/7r6/lQxiGQTrdt6ptl6Yqb
wpI8/8aL1q5q3alsWIhraAHAu00kw2e1wHYMqUu11LmLcV/h21Cp8KLgH/VSvksx
KnCdFVj79CHGZNbd76brEZu20adEnqD3nY3yZRZFNHnEbq5hIyVfF+x7XFxAptHt
OBCdENxfJMHbfJBGBZ6US9SG+DuFaEf86BRn/6i6BX1g/xuCbb71nadajADSyvX6
HdaPEadc+5tKXaYK5JNu3QsqMRcmGQfTbHGi5MDZi0iX9ek8Ym6d5vNMyQjZQ/sm
EUYa32xwgjVGV0C+3b58bvJUN///umt6S6l0wazSt/2m+9f2z8i61n5VeNiLoTq+
5N+wL+Qkm0KgDrFFXwQrgBxX3/wTWZ4CePUmbyRDMT+qBCBC7UVpi29GAEuwgu5W
jISQLPGGoqFdj11mt+91dI8VIA0k8hE9fWbQt5sbHc22QB8z+XV7OjhRXHLhvFQg
Gw9/eEjNbDY855Nbp9BXyTNoNNcYLuhvQIgiG9Kj73ahJyTlqm+GmQrh5Hjct6TO
baDfQsv0Co0FPRTxglupyz1PERtomZgf0gB2JkA90mRtw1ZLsvKiBV4RAOE/KL+W
vAjn1k9xIsesBGbkrP2HhpZq1/gxGVz3W53Cy1u2EhGflhvTPhDEVMobjUrj6Gto
UUggyWgOgy6AgyJVE3Wi8fSHhXY8jkfiiQNdAuelR+YMVzdv8rGaOu0GzKdJ5+Sn
eEb9ljJZHnEm6/Xxlnyr366jxzr58BUwd6NBjrVpZReGuUstoDGIxh4bpo1hXnYu
XrhfVmZb8IoFfEancE+8Uuq39pCSWN0u1Sg5TT8fLLfXv9z6O1sasizcLTfRN+dH
JHSvG6oYdqgWPVL6SZyNryyyP74HHRYv1TGjpSVlmUb6GZCywBCHvv9PBpnrJ/Kl
mZxkEaoabkbgyTTl3+HYTRguTgZflaFbsqDD8yx38PEdH3M5mfe69v+yi99ZrFK/
CfSQQRJLsEj7qXYxtSF+f5XM5R4f5xhwcq286ZKwjYzB254zZd9sot0r3+llHZpH
NGIX9tuRMiteehz4VF6Ru4J2GShSMikUdvOztTiL5DYKLJiDZCEIIZi7v8BQI7He
S0f+HSLIAeMXFNW3Ie7IjRmvISPQ4mYd5E49q4gVBY5B0QhrUzcvcNN9S4aRxDsK
/BAVpWYt1aowAMXZ+gWTF0+u/GESAlW5p7DlL8lcxy/zfMtoPbqRKqGgPMCsuTdG
Ni2vx8/Rv/elJbStPYxS0M8k7O830OPsQoYu4h9PRmltViCOzEtZH4PD/2/ynymW
Or5gMg/7ye0fw91jJkpjTbYCtE9BXjuY34traknxLyy5QuNlocUuXJYOIM1cc/zr
sWIM+0VqYq7uhyFzkb/F7oYoRqZH/ee1R89K2aYobLkt3cHfS1cMViVKG49jUqVV
J1mhyzvcohVeWxAz8XuWOolGEy6JLfF17b0mx2eDAEB9+7ZoO/rcrkCNrhX5Xv6W
SyVNd+vQcLLFMoJMM8JwxS/U9j7a5u2FYYT8m3JiUwC4plZ4svkJODuuE4HY0zQ/
IGMjFI1/oNH/4UbMKxj2gxEeBro2WO8yJXBrRUaOgf+LE2r0Z/a4uqxLfsYE3y9k
yefhgBEMsmYsQG6KHuYnkSFM8yHrRdKbtH1WhYvm3ZqyLgLuDBuxNsp/5JJPUXjw
cIg2G+wjvN4preXzE+jLJI10wkNVFIsmwnEm8fTwbWBxSAmysSRG04UCyZPvFT3F
OBZFo2aA0vP2C1QxyIVGKiVu0jgLstx5ehpfcx5+sgTyd8RHhMBZWjoU6bk9f6uc
3hRfqwgKm2eXpe2MN2LMKwu7merk+bAFGis7pHWumz2kwuG47FKJMfqhGJ0AE7NY
UxW8qW6ugO/87Ze6RG4LPBrMncBsKhw0ZOx4aw3lTcfTcDWknfBz5dwFcFUTTsRx
fb3bmQfwlZNw0cbJ5fV63ynduo8G0TiEvb/ELHuyEW8xC0yw9o6hTMO8oTHaToen
dWGf3eZOqSdJfYzMhG4h7LR/qEI/Q5EA6Jszm7DkqlPEV/jwZsly4vRTk3HF+eW3
kEaZRSwH64r2P9wdV9Q3KOgkCLqPyEMzBAtQyKLrDDK5dc2czhF4UReyoG4xBrKB
SVx8Pfjm1zM07l2tHreC8JJJ8x/CD7rUAwR4pYluKUapZJz3LPDpXCxHxqffCqrC
y4I+8t2SftqvkOottGRK+ir+uY3Pzj1udpx5ARgj1zya5bXh0HoqdN/g5m7O9fop
u6bEDSMPU1YS+Lp+nXpOY/YJkOZ/seNJ/l8D+qfbOPDeFbbDoIzEB1ECuhtkOFrZ
Vbo7LzIDC67t7QqgSEiOO8lxJLF9oTbxa+e2Y1HGYMa0Zbj0em8IKG/LQLoIuNiw
REuobKlB4HZELY4iC2yJgZ08iw3Ta+GP5M35i8/Rag8nVWzWy953qHg+tmjGQ5Yi
9OeE71hTmPefqx0G4tsnqybPCqKjM4HGnC7jOH1fxXEzDW1KAZXPfaq/ZhAhxo+q
RTcomgfJ2nCXTFtSfAsxxYnepgNX70iWnkX4PjMC75fN6fO6MgVDlybLJ/5+keo0
DZ+6JeUFbq6RikbAZW6eCODB7KwsZzYjY/AnzJF4xDdUXMHgt+cnBzgD4m6zxFdy
s+x41R2QA1N17nBdkJcBA7xXytZxJmvX2Hpo0TBQk3yBvqmQnudSK+W33qby3B0t
viAJKzM4xhFclbvwJ7xMGgA4lEG0YBRfnCoEtncc2naSUHAY/cV+S6ajR3rWvXRO
1U/HbeRIAFz2itF4PKpD/sOvh2JRw+OoXjEF5esa2z5EBIhLgtl1oJ8n/duPVbmY
5R/HwlUWppPEY5z4u62FhB4QeAtNgA6nBl4hgZg5nvQhLFkYMfZqFqBbPVSjPRDv
MEr9Jgy3THl6g1ehbyuexW4kNujlcW+Zi/XkXf0sdD7qTj5jU2Wn4XLUMzArSqkU
N/eS+yGBSJD9PIbSmCb+TKe0edVo3NCrsd14VQP9dhzx6d3NB5sL2AAQQSCTdA6A
6tudHhriNgbLRdzlmWGYOdeprOn4yFZBxIc97gPKM4MXvBT2qZzJNkRwOTmDT7Mm
68phi5ci8znM98lbjA16LHhKHBbXIMb7H2XHehkqxAjW5So6vRHWSQzXOZyOlmAM
OWLqCOb/afYyyOkd1y+fdKmper9rBxZG3Y3bj5YY3mZ/SEBE4tBhFgwqrsxOikcT
FZMZ625VJCjq71AjNAzqwJiR7AIM51RkPUwzkQdG55ObRFLgrIgJt871dF3PF597
h7WAJml0oYciCcMSxS2rmZcHyBS7Eml1C8Wt5ZwiqTFZ8692fWjrkqm6YPXQv+Gq
ZnAeZUgwUkuVaMsl3cD+RL2dINdI/EUwPLWAl2FidxkKFXKI6W4YmE/7Fy+/V/4A
v0F3w9G8A9+udxHnFDpC7H+3B59Hu7U85nvSE/k1BuJ8vjiY8ik8YhG/pJ+o239g
OvRxw+2gW+/OzBbikyqOaICWYX780u0dIJ54lkcp9M+OgVxzemLq/j2NJu6zneAh
v2NzzbPrcosBVVBFFQk0CK2oVJehzo5fEY5z5A4bs2Mds7RKnfiEuatX44eVJsv4
5TdNHjLs8IJLWNwP2fGZ/Se1GCK5ynpP6qFlwgukZFlWWvUEhbq93aX6TVOFQZOn
/faTF/0EogYmOpzICU/krsgCU2EOXLx5xQzTkNkk1I3aZ9ZJDHmBi+D7oB2OlcB5
RNPevhTgKCHvSTHutEP6Y7Cn8kBGNzrPSKh6iSTFk+v3yl7G8/ct+n07NKEl7z6r
OSZ/erqZ7mt2dusMHHbsPltkZuy2mi1diHFjmNXytbpNzRXYhuJNYWOwdLb9NBgb
OJ7iV5RPvOduJm+1PLr2alJL2fN1un6aOqHaAowgHKCz6uNzFIyTMrCwCYqVEc92
uoKKo3oA7MWuN6gKPFrSfbbq4/z2YzLrurwlPx0/yMjzeHdCYFGbmKneMS14O1s6
LmWNYqHUml9N+TAyamuAWQYTd1qtecy47kakVv2m8MYpSTMFqeYNNcgRl3lV7c8b
IOSM7nrAPBlkmG7Jwi8CKtpHdfgKX/GPi1sNAlueRd8aMYERMVc0CjXdcHb3c+CJ
kE7/G5kxyoSN/eNSJzHkzHOYSajPCXMTz5I9WF4DkcVzs6qnmMpe6HP8GP6zpPR7
XlRvE+Jhx27VNlftLGXx0X4/yJPBPd0BiJn8fD9jSy0IJYBO3lf+xWNi1bFJXFu3
GB7qb3M6yqVmd6bACHA35+kZ0/RDr8K+hA5sJVaLvkGU6rHsncUgUqNj7prK8WyZ
3SNdoRnnkA48O6oWxR5fkRTCLUqFTgBoaIBowFXhUBco1Ydq9SENXtke1bmI0PAf
bmn4HR3rWABQs9LI7H5JEXC7sjMPlwBYN893BXL0VoOVBtfKI8XuTHCMI9B20uNj
/sezyLSE86O2W69dlxlcCZjuCvKBedSOvC5d/z7PuP/roVAFTR24IWF6FT/SP1n4
0F9IpdNPFmgXsUTcQMBYn6GAk7bPU3+5YroOGSdf8rgjlJNTyxNFOW9DKbqa4yLS
bgEq5SGm9LzeUvDh9k9myNugq6kO/VI45aq56q3JZ3NEGh1IQtSawLEbpURuNZl8
Ln5wa88Ld+igiIMRwBSRbvSNnDaXRgnRY8KnoadJzA6ad1ishMdiIpzYtWBt5dg3
V5q9BoTXV08GOXnhMjycVIetsRG481Qym95InJEcOCuMYhyOihNb3Y84HVEmHEjP
hIajEpLMh/qm+Nry3sbP231DCfHZ3LmZtZlDm5LGVQe3ZntjbaUzQ8me/prJ4bht
i+U061b7mcxHeN3AJJpM/pv/9UUSB8PkUkUR+09q0/bVSjvVrFWaBCpdNFGHZUIt
joIe4mBPxpVBOE9AJm2ISUdThVvwXJosUn2MQR36oQnE14DEwsbYX62xqRL2PwIB
cwTBEoi9siA5dZiLXvZXoWur2FP5gKTeERTbvNriUPpzkB8s1XvsFoqjmfn7+Uzi
5b/VK/CWzw9xevCk/C1YFr5AdjfSYnB75JQTJYcB2ii/EVs+vB/wI/TS58qZ3Nro
AcJd17U3jgjia9YIX63gQ220yaa5xz1187kO4uADeNez5YHG/DflpvscTn5UCzeP
CNJMmKZDo5VFVU6B89CtRkbBtrazDJLPjSr+sIUHlD+YK+6ZrH5cHDPduN/LouXT
Do7modTSiGXuIk1dLZ2JyPxnsI6/jXSd2EQAVOeng6t5kR88EWOKbOi4NcSgOfNm
vNvrFUcuPfotpSnDnfU/w5i+F2BPxJZme2WNRGkXJ9WU+at2xCmX2i97T++vMwNP
rwMTpbbXPXb7yMaoom1k3elMpdfhNPr7CXpSlNpCxXpCIUJ+pyNwL9dpJO2GEhQQ
PYQ6YzpkNIeBKgdxaIiFyYzdX40mghlEye+yv2HnNS+2tYRcl+8Am/hwsLK1mdZk
n/XlNnXYNJUY2eiEHlY7nEsrE+pmgyIWGenfXHFH+BUchY58lJBLwGSiQYepO9QZ
jdWbtUvkYd8+ZobYb7UP8E9Fy9lzDspMebqyOC6UL47UBPr0MbDob48xdFTi2sHT
IfAziP0n/P3iOfPlWRvaJem62L9ZVogFW1nNv8cUQ5h8bvb9VVGSRVQ22Ot/HY+F
Q6xKKYQQmx/5eJM9PRvN1tdKQPmUed92ipYmo49FcYsZXPIqQ+6KslFLlj465+4b
qE5rFR7WDRsGgm4+ltQ2+lgTJ4wYktVuenUAjFbEImHyv1z1WJkb8KnkSccXQ4sj
5tHFJA/MXURoaAjmf1tRQdcdeUGSYBk4xzwsLyrVsWGQwtHPFns1eUF8icpHvYH4
V04vlm5ElghzeYBZYAfRnQZYUoQquMIitl+aXP6wiDAz+ZO6l9VJq2kQ6Qbe/ekx
i6Mh/5MMYSErdYTyBeCXqoLhMSsTeGmlDkVqE0RdcU+UTN8O9p9g8ZmYro6QRbht
5dNHjyKsj2hUDPvZcT68e1K8gkhFvYAp59kPe4Y1tGNAXWO12pVvBW9ry2JZ/CCO
Zggzzkk7etTFvu+3kw3da1pzFwLJtEVmq5xAVBm54FLeLC4sBBD2oqn9XhQIKlgb
CPD8iog5IKecI8zC9qPFModvVo9dsl5yJC2Oas4yfriRIspPcURAhrL/rILajmYG
9OGHIzkAlehIs6dw2r/iCHl2WAz9Pli0CD63X1yt5BEayaliPuTc4+eleQcs1ryg
NksqsL7BtzyAlINXIoZSHIWkGWwKAsv+Lvb+jZSTcHlRMFbZMHsPYlpFp2cbej0g
rkZK94z9LoybqNMNMRYilM0Br/8ErpkO5bcniP45e2yb8VzVxtP2h15eCW/xpOAR
QG32tT64VaLr3fwaxp1/QcUNV+7ujhVd2wi9g3fmuHfPeH4B8HNVuWxxvzizuiQn
hPE42ZAc6xQom6PrIPsFaYU28dF/NhxNTgbURDU9voBP9tEOeEMMkbhixNZiIpQl
MRHyTzEdRxs24FupX0VoIAJDij1hbkowdvJjEN5GAsTWq+otsvg2pWPoIQJ8EpVw
vGrfq9T5iOc3ZETPUXOLHFJyFvYwwUI7Lrfu60h+j123t7H9INZYqFA129PGHteZ
xlB6R0UD2ciBM2eL3IDtWxO7sIhbgm2jGagt1BmiP1bpWNhcDFGt2AwGfAl8nGQn
mTCJ6A6VgVlgE9tXKCmqNoVJzU3k3qM3FtaDLn8UlylLX5mhrPZCk1uukIvXrBjB
sEguE3OgjL4ITGcqrd9vN5qO7+V/v0AGZplZ7BjOSZn+r1Mht3Fxq8Y19XOooU1t
BLY3bZBFDxuBNVf6up4hcWLc/tiL7AcTIlNCkA5HCHMLAZfoMPpgj3skIEoZRY7t
fagNUZ8ESW37vu9FjOS/manBcj95CiAkvpo5s+hS3zlqBy2dyyk6delR762exsVO
lggMoDkkUn5MbV9yJv54jI+gJj/1pp2neFcVmaiGmgxhhTdwhcTGRq2iWiL95FnH
43EkdVVUR2p0h4xRP0ealX/1RIhQA9/jDkQCxNL8n2vN1do4fDAK4UrVsQwJclpn
igFS3A2sv1k6DDf6MvJkxjjcrdStgjFmgrI5zVJHDCgeRnRkhQPMPeQVP1bOPU8V
dMMXAsu6ozsYReRQYSQzlbC88KaNb8aN5131BRaT381JQCEyi+5n1S4PitTRBziI
iXIEiJh55TjyhORkIJIv5PIy3ABS/1S29rU8P5k27zbznGab+ewNGR2akkPOZKdP
/MJsWIrKJQNIsYvA4lyzF24BfLh/A+VC1C6hZNiqfvmRoBQt8uG90uBH8d1VPBeh
mwmkfBGzSS7pnTD78vstjBJt6tR9tU/a5KPIgYbOOyJPCJQ1qd2yiGy+kQSXwuUC
3RC/Kz04FmyEmvOVvlbZCHgIvedzNRm+qvp17RJsEtbGuFa+S1+IQlsexgC8Ulym
XPredAoA+IKqoqtLqLVtjgukhrANZUbmRHfZTKglQ1AUHESPu5XwzxqrLHbTYYYf
J8iEJ1aO+uN+iCoZge7FQIpQ9YXeYeqKLVZZ96jdhSCYTvWlZ/9WexVrXTQiR+Zb
t/iYEYYEgGeRypBznGIfs5P4IoNdGy8d7RNrR63m3lSsk2ArTgkBUrw3yOThQspb
hDE6B8Xn6A8fLC178IALuPsSwzE/bRXYpTuoMawTaK9Xol57pSXbFRj4RhNhEWVU
zR0d4i6KJwCE6q3/6+XmyKLu2iU2ZIYRgnI0pEWElWXVORQG4aWmzz4ICDAX89Nz
YWnV/J1nfkvqnbV4csYbd6rbDauky4fBRvhvp3uxpYGiBSqK0TNIer+r3eMEC+Y2
dtL4HbIyrScpoJlA+OSq5PlvTmJNhG7AMLIZ7t+N84ILKe43YzgwuN9EsAfMkwta
Hfg2EkRC1KC3u8OtJZ4Bht2/v9YjMh1HR6p+0xE9vq6My73EkL6TSO932J94fwlu
KugV7awsOSGKW0HJb9P01qNfb8nogz7plV4aDNdL8oF1MErnhonMGVKUvdscjwti
KhPD5Er5/vhQcKAXJM0R9yijv74OP/TrsK6DX16vb5D1K9KZzDacEeTwSf8jctZt
nInIicbdPdXGOEer8533xZDnVwMwIb2+wb1Ray3RRfWEb2C+rNC1FocNraMUAG/S
7OT9KfO6pA+9nueYOaztzaZT0exWsE/mQLbvvsTpOFZBQvlEiOIkt0OzYaKz11pr
eRX9URIJjff1QyOaUiMGsPy7IhFurxbQWli2lla0AsVujPDOVx+v//bX3kcTzZwc
gghYxY6R2S+E65hAqA5KTVeHcVpJ3hc2bmBIS8bglAwPJOhFbMLkQQdu9CLq5dfL
Ed1xDxhobO7EtPIHhIKbFOZzKMCbOuz0QhrfA+MizWwFrexom/MRThN5xjcNJJSD
KLLTUbGZHrLG/4lhGfy9jziFUaaL7UaqKv8k2cpDim9b6yBHB64EYGAFJWisDWCn
pRkkPImrDMxRj1p/FM9jlZD3V8MTp3JTIxXRVs5BiFeFL76KSkKsscDMwxBHAA9p
XTL7fkwUc/bLXLPXrd+XK0Ym0YUsbtvu+52JHjGGToSilWz/YJP98NJMGLSjTCiq
WgAFYrWlR/tMyK9Ak1LyVcomtJz7iFOM1dVj06Ccqrflnm7ksIzytRCnqZi5aUC6
wG0tURR31IEf9KS5MKrgjMyfNVCnPdOnc4z4uhFnfcN5F+uQEK8Mq3kLD5CCV9xt
9Q11cjC4QSP6VYVgcpBU2axclpUoYE1AYeTcnFdqRclOQs0ao2Zv2Z+kBI38YszL
3MZbemZW8TRqHddngCFaIAA987mIzclI71PgSeV4duwkfdEuO/z5b/V5Z+PpGVz/
eME5Z0ilEnbZO5pVq5CFjlc1oC89TLOUBrR1qVu76hZVEJUtUr2wjqRU2y8SCk+O
YGLX/wuMMNGX9fTuB6eOb7JSOg7YhXUy83NXyN1Km/2ke4CU6lZIn2UJ7H3esByX
ym5WBxJcIG8g60GbHEHl8W+24eGalKZyISG3zz/otqk8kPMDw6RoQOEdszbAxGqs
0g84KKj/lwuL++B5Vdtub0GOYBjWfhj16qlu5nliExY3+WOJc/ua4y9QDRyiMv6v
K5lFCC50VFqtD7x0CU9WyBu+8z1erTDVhYPpAu+oFlrixV3V7wIVxYx+6bhT4V3M
tRJorLAJM1w5+C4Hh10hwrBVn9YFQvRp773PWh/JZq+Ukew3miqY8u9bdM47Ynm3
NNxiDzIXHVyrQpV4VqqHRMHWIqBEKZbPLQ8SMEBh/QUXltmTq8ONczBxdDFxCAqT
RR8is4tvImwj5zhIxpVcgUdih6m2qdZXL4GVoEsakvA4ElA2pdZJMShY7fVCtqPi
YSVjARq4zanzFOkZYWKGVizzOUDDkB+l18VO03ZuTsDBacxeoy+yN4rrzgTUrmbE
FIflFu1gteSbhnu8Zf9bYYPkKSEgVGSrFrCuIT3mItr1fRjFsMdMfcrUpPec123g
tWeG3lA2xY0NVa5Ytd8gNDVc3DojoJqy1eyvON0g/4HXXEJgc0PAs/yPqeDxc3zv
7HDi5ceay3ymQIcxGBhVyL09RGS1HZtqD/9CCPaU7gkreX4x9W9sfcMVE/B/nO4z
iFlsyOUNd6v+fPoNZB31KjduE37RRIblbQBKirONQL1fLkPP/gUM7jz8qPLxFCv/
UQxmSwYxgAbQ35Oy/YmJjbRp617Osfh4x6a6vEHvYWnDeQMJTLE7mRR9ENrddfef
ct2Pl7ym/tZBrDxm6pCjYhT7xH6BfWrTFkpmnPvr752eNIW6z7xyB4FVRShHjXCg
r0sehN4geXLXAAIHbbsLehLSdDd4W/oecmNGee6/JgppznoOC95AMJ0go6h1Vwxv
7+4JiZ2ICLNKyMZWiQ+bMxd0lC2OKWRbLDuiPOmqxpXnQY9TvzEfILEPVm4Or9GZ
NLlOHAv+4h+NkFlyV0RCN1QxZyX4AxlrkX244MUtdmEva1RFssjaGb57PaXBSbgW
ItN1XAznL3WJNLLNvEaEJ9QYAkSEJdRpvRXbaPQ9S4It3YLYC/5CkOf6J4P4aU2w
ila2fDujVCqmIv8eZODfibZM23HRuewdcn7AaOasP6Q4l9iqVYv0IMuvLrjZs0tY
oQhlHf6MOitRp5UwYxWzQnnDkpLad4p2aqte9KycpetlHnA7ioc5U5XczmRBEjPP
pBWUe6XM0uecV/ABSnMbjxxTaNfsmz81A0/8Vll7OOh8B2byX5pWA2CKgDHL1e+U
nl/YhVAyjLPoiDt/qeqPfKZ+VcMUuxBpRcal8Ca7+e5Ixhc4a3VSrVWvww67rHig
obl0F/pujMK72NWNJ+ugQG4E2RYpPEcqQSqXnj5RXZuBFYoWmx9mMTL4Lg0imILc
gYjgCxCF9Bda4y4vqrkIsDzu/YkGfTkPwL4HBAwy+NOuFYmd94TapXI6lM64EG5l
lvDZg/S/Fgv5LU4YjQcytQon58yPkTCzQTq81wX0aQ97kRyABIBfr9cN1eTs6QLe
V9g5Yp+5I5F0X2eRo8DMBz9qoj6BpwSJ5oU/N6twqTWDjldsH2/VaeyIhJ5LyhQR
M5MKD+Svfdz/qIroo3c5h5FiqEpD4TolFDhhdO1w5Ld70B1dNyb8sBz1TIc7CsBq
T0jogHqjhfg0HbkBgV+dxKRu3HUSqtKhQYq7VQMLFeyanuDEFZURWqs6dE53xblr
eFYtuOATBcxz/l2310ZxUULFwNhYXxLQPZGBATArgix+kwysdkueCxH/tf/ju4uE
F6LsjyxVIUVRMgMqyid96dB89ydSuYd+gbURv5SESLO5K5jnTDt/YJmSa5u+Zci4
t16j8Lu7dl19oo/bv8Bj2WgOX6g3PQ64ZDDI0bxBoQfE+9ul9sHoW1nEqeyGArOh
pdEsaCJV0web5NWZvp1DVLx/pTkxcWN7iJXP85VcDdArYIzConTMCYhS7Q24RL7n
2hSECuya/7vvVGTpymwvchnBpfqVB5Sll/QhOtEE1kNxUKpgeIGcO+sh1Pjr/RCG
/IUAYVwiE2EwE1GOWt/slNS3XOndVeOreKtlALuN94iR34LefdTHqhYYi3puOR7l
s6NBmM7XeweJ1EA7bCQr7UxmAJlHiwrRMwx1Z/AJOjBdzD1pq1zzuIZSEyla/iQY
fW7L5sLSFMAv+SA0KV0mHBnt6ZabsDFUnOtDrCSC6eE/zX8CTXo2LCoKWCYXa4+U
LZrJyBMjDXCbMRGBLDoHvFsNMrsUSnAHcFC6KfbS17FaNU0JdFmwp5NQhTKEPfeu
45KXTwurr0kWxtoLU32M1vBqTP5GqA+F4J/XB1uMpxyxTaKBuUM4Xavqv5DAtNdX
llcj+hiJRuKd0QgSwXImmfKh+05G2jGtkJFjo0KjntUwIPHTL9+8iKMhi1954/Bu
THomb0u5fVhQ5/NtIa5mCs2nDUGQoHeDnKfmwvYvJZIra36e66JPpA1EZMpB9OKh
993JNJ6RUkRD4ItblllHDzdfTceJn0P/YlpTR3JjZ6tGwC3v/SAjS96OE45RBzWI
Yl23A0+QD2w7CNwOougbk9hgGqleMfFDkYPqIId2uWbwXp7zFuk3G77D3ttJel8S
+kiY0lneIuUcMnG4UfqNOW9yVtOBPg7pxeqLLQGeeHE8xobkTo7CmII4vuIntySQ
sgt9O5bjk+aCMv3F4hEz6y2EoKO4lKBH/2YNtulpIzfpT8N3oAqGAj3kEbdvxU3k
52OXegBooU4ux4uwwvzX6VytzH+0BwqhPlbfkCXncsX5nehWekXY7W+/kNbcGtIK
qXbHAMGYOADv0FidPHZob7YL0JvGCNFqFwEtl4rX7boUdFG7ERC24XzS1m/r5rQe
BTYAeJyn2wiqKcE14KQp7S3vZcLgsuwI7Az1uS3b/ggfU6Zq3DRo17OexVZbB8Tu
6KpHx9LibZcHVMnxpki2ibrg6ci4d7GzG8CbX7Y+cz6KX8YKxlLm3zy8DMCWVuIr
51VLWifdsiry2fBd7557/NXk5B8Im5kDN5wHtbFAksKKXIE7aQkFMO+hfGpklPnZ
JBPGdix/spIv8r7lCk7cQTbj5byzPU/gYrUI4kKFip5BV6nOZS2/TpJ6t9Xz1hDS
iq4bHqZ5nzpHhuwtLH+RxhYKhXkIQg0CWf1GiFGT/LbtMc5GX/lHqlXu+Q9LUSb7
K/pnurZVFq+yXQHd2Sgv840ww37b/ilGkTTGRuREB7JTNyyvjPXvQzalnKquJzRN
ES8exb2J2nujmzvmGIYo10wmcNZQ+g7r/vZCV4xYnpgpu8wpnhslgOYIlP9WENma
EBwC9T8+VWSUnKKqjBaKrj00glwki4swvfwpzacw/FsZmBGLPv8eT6bfwayJ+qr9
z3gjOxaLZ7Ph0lLPD1bMxqBvUkhbkY9uHQaDShRFWwBMVhWJ7mSYS2rjRYA3iLwq
D+sH1XOmfhAXOwFpaj5IIeo80ySPdaLVT1RPx/5YTk+Gpui3Z0QVsLsSJCHVfjm0
OSbhL8RwcVIHfuZFfdnPF59X1mB7xun0QwIn9tQYJUax8JAb3S7bIJ2mCAuZQPSH
re1ecErdO1EJDD3T8Vhf2ykc3mUXz5S5o6Qi6UJUEDUFdHtnzjSrXClDWQv+fWAT
+OE7gTINiApuLf5IlyHAA/ht+u5zNerA55h36DSvsZRS5HCq88QCP/cdH5d0XM3f
Aif9b5VcUpIturFDdW1ft0l1nZUWCi8IAScg5cJ9GFf84cTunAKyCAz7oP4CL79X
jb59s7gnRKb2sXNFSuCKFeCQWqF8AEcfA8B95dDN7/ojZCzieP+iaIXluG00gT/m
d5q/kzD8fzQDOMqdRtejs6Q+wDdLmU/UJkkaNt2lNx6kZIDZqngHUiNE3nBgSSqk
4RosrEwTSObl4gOws81qUbYe2AWSUwUP6DUPJLEmyFWOV4or0wWItsNI1MEZ0BjZ
Jl0fuqxkZmcTYbTdsY5Lz6rfOIISeRInyiibqEN2rIh8hbDkVBzTGdxI69f7btjn
ULnlT4IEfV2HKx8qjvE2Vv65mBvqTjO6v2nE+yqYOwYwz77TUHioZECMykAe2Q7v
jMG5rBJ3Sc/yPL7x6tCbPPDSnuYr9TBJWNQkT2pJ+uI/GCX0y/FjDvrQUpWckgom
zy+vePv1Il8tZnTr/TjaFSqbuQ+P32Rmi0rPXOm9gkexnM9t9cOoVvGyFXgKVKiA
tfQg3pSIoangQ9rSLhzuK3UMeCj05bQS2oJrLiNCnKkPCIZ5i1HtMmz1vGG7Qy4i
kJ6wbVah4EVx84ia46gpKGFwc7shfqAAWhlOkRiSmdXeG966PcLsAORMLzCP++SQ
2NMSQERjKGeGj12gTllZ0okgUg+3IGmo6finVQLEwxik9UQwlD44Fej+ntlQoVPM
QSPx4ED4J24EAPFTXacEPj48FS8Z2q4vrhYeYJhtv+yhbwK/WSdQeD5MLDystWxs
N9i+5MRbkYYiWG2HIYS4N8BJBCDHRcOKs1V5bfk4EC94WEEozE4olw9iEDurP2w1
zwDjUtyJ6XgqCyFpHE/n8RuWYbqtMlnWa/tBmCfdNh1oycA4UAZpB82O923PDJhW
Ot+LnhGDTVZmNb31W3zVas7JG8cUqVPFNov33B0IuuSb+onkUWGR1t3o43HBZOs2
tw+lGzK7wfoOTM9lm+sRNhk4fVy3t4Gsck/cu8IUHcDbOKa347o5FQ9z6fLyDlsf
HeOjlGGwKCvb7jVdxiMN6g5cfH0mg8iMEBh21o9T9sLSl4RUKhqtpON3M4tcNvdz
pZwSv2Uxt8BfGkTYAtX1Fe7ZGdEJBuG+lvk297NpkCRYqTqQ59x2dp8LdaGOUBa5
GfSX7E3Z4cjvlKNhxcmtH2TopJmn+yDYBzzvkhe7j2tR5Y7/JqJtK7Th/SxmF7Ta
b7avnTLk+YpfLGSxVbr1LoKXOH+X/QM5btCSuzG3/4Jfbw0SDX2HZklVR73GAm9L
uuJ/IFdu+Pl2jvukvspNOHXuDnUnQTF98rUzS94MRrm1AGX8rheTl+0MQqQVPs7Z
LeBXUJdYDWVi/a5Dz7/ulz5QANjkTw30xWYZ7c5FzEhbrPrQl4thBB7r4yWxWg/r
BLlXfsYQAwbqukmmkR8XtYgSCDjs6eNKWf3nK/AjCkiEZX7o66uAENUdEdm65OJV
WYZx7ImPxmMUx+2ke+wv5dilFBuxTxRIdan6M7/zqlkqVz4xEKhrSdXb8Gt0K9t3
FwmNTm9XJy2ItWpJbHwXIX6xGILQEnC6E3cdQuv51hJ4kTK5tABtkD7nOhJZUhPc
LOVHBKVTCdl2CYpjOaOFJxi9QtmIQ4Svl1dJzW5u0/ZCZr9Yyb+QY72ienzfV7Gm
z6xJr7x+aeOPFQTgVTLUa9IIS+c5qbRQOyPik9fnXsBDr8KqPn4cNHVNsLBb9sax
3GfwHTEUFoV3z73Nk3qKdndX8VnQITawcnbagsIo1l9OdZ79nFM15j4IMNnVSm0q
lrLoGZQdaN6rNOm+mE5dxYp29dy9JzflhrfNVqivIa4IYn/s2ZgvqvNdpjXHCTNv
vt+jt+6Yp+j/nkA6LsW449lpYirZM3/NeAOeFIpWewwlzwEutXQOF563vvcQPdAw
IhFZvcC+QLIAsZU80BJgOuj5yI1hFhfzRKZIDTQKwuRRiEtXHMEoGSQ+MwcJ3YFn
/YOjQOv1PtXH8Q6/Hp060Jll+260/yL6Ro3NxueBVrdLBVtmxPAA7vKeKH7zIvsx
YwnzCEPsEHrCzI2rmPsQEXvW1PUh/ECtNeGbweOqj9cbDV+HtqYppUv6y3bLZmiA
0+c01x10DPUtViTwEz01jnmJKRG87N99GOcPgTpK/DyweEL/UJHa4EBkr5Lqwps0
3oAXNj0Zy5R2ogZFmW4fXf/IgaTv8AIvOo7HO6fqP96utAKs7Ff9g+/V6P5SuN48
+ZRZ8Ka8o5TRYh2evENVd4xzP3WlGWxsoXq9KygoxOwfbwFXzsr+pyTZJoDfQIWb
pnO5n0tljuZtsNuOEw+qIRUT2VZm8Q0taQbUHQKqEa66We5A8LnMLbc1SJIcFUTb
HdP605GuNMq4bVl2CM4Ks/aBrJ7lr6RDvUYYODYjEteB0h0pfK05RhRhmO5S1HmF
66uII8ETSlDCdUY0P/p8tCCBUbvdlmwgBIwd//RGbYVwVNJ3RO6V39jHwai449gC
sFyiO3zD/AuUoKjnbpKUp37vOqbF2n0kXqn+lMgCG3+sVJIyabOi7Ia3MxQi6Uq2
HA3RwBknfBB46XP8B+ULfazIfVekheFDb/48lFep+eT5WdnThv5kYGKpBbG0RzPI
m7a78DABSG4O3VRvvTJrgYJt5yP3EtQTbD8vUilfEkS7ghkgO3zFCh5iC/UjMpMN
qLamcudfeNT9WUBpNcBLLEsmA9jzNS6TpoOCnpd6bajkBAgx0b3Ro9a9CfBSfhFI
PpTFLPZYR7ikLgRv8JV1exxnZ0gSNfQWVQmp43NefFz/t0+6340MoC/VeAjhb3eC
+rploRbPDpLFuRGjK9P2lWb/i1DRGMW2sdtwmXsY0SwHSiv/0CR3ZjeqoQz6miTp
OeM7RkLCNyZTWADJTXbM9dCcAlHx94rfV2jx5BoqdEaQRh2alPZViIb+bljjZH3w
9HhFd7uMS2OOIswPMxmWNkedEJ2My20fjMZ3TSU9YBU1W8riEHsqFEMoldbktSAL
y/eCSFBDA1o5uJi2zNoKXzSrAUP3wu6183y6lWHr/fZSz7q+kknOk0loJxvwU2ZB
U1xDIQvpoP6okttrXOvpKHtR+xfyRQXPKMwd3TACOs14aU5DvQrjuGujyRMopIFn
1eDxUdPyHtGE2QlKEhjHLhfWnNQmDjBnH/rS+h8r//EKUlo4GfT4J9M3AJnS7WeR
xDm+8IVItw/nyExf3S1zs3gkCwjA6MkIKUEztjyVjhSr1e8QQkcOxqygcysDSMzg
z5HCJ1rI3zDCAksw8xYbnpNOzxGwDrC4NjQegutFRuDTVXXqhLfBh1bof7KpG62W
bJWqEuJ8wWmnFVntyswS67XpgcAWRF0NxrF0/wOg3aRqUAHRFEt1iSN9d3ilMQnD
XdzJ4ePuPMUIcB8xGIl5YiguMaAy03rgac7ew/MPDgP/kbXH5BYq9uwB+Q7dCz7p
JVG0k+x3ouP7zIX6ZWGei7aby5XsrphlmSGefNzLA4aAutf/ie+5OYlzXed8SR1s
KvbH+wNIIT6RjMRrIarZtIOSjp9I0EnuK8Lt2nYRm0cZ+/7OKcXMXD0p0hVBeWZR
0udJFXGrLPuZFTkxldwaazQnEXo242QL+Nj9pyKNIPaN+QuNqSnY2nURH5HD9Ijn
G17YDiwh+Nq0qZDee+X3zNB6jYFK58yoGWth5Ah1W/xiClxVPUj7SCDYbdbCvpMj
eftW/8GQUzvnQGSoTVrff24NJSHaxtINTc1q53g/RTd4dWxXbsqHV/ULZ1EIDuMJ
05sDfc/x2gb7xbvTdTezb5xVd57I1c/d1PTLd8wPa57Np/E6NJZMbkNtPLYKzUdb
y03MIEDv2oFgh23rb1xW/Ih7/zk3YgJ9CFpgCdYjiST8v8q78oBGjT4P50+7bxNY
LxVvW+sgyTqSdqG6smXU9MCYw1KHB5zL1atIPAJYvznrypOfLhko2PBk7HC5MAqE
v6Op5MZLX6iEe7SgBFMleky7F7HnbTu4sPcnrHFHYTq45/Akgo6djwCuKKQBHBJ/
7aN619vpR5lfvKJBLRTzOYGuf8wwqiH8Ka7eBl0b3UhvTEGZG8Cw10vmyZWOIYf8
4e6Hfo66QlgI0vqhDbrhDU0WKe6fNozdoThogTrabAgKsatBLTHUKkd7sEkIhOMT
ZBV055WdWcRpx66pjEox5yd+jm1WX/R3FQ2Y3XLNNqUFhhvPP1E+EIjt9jBqkeIt
pD6NfXl9e1wENT6i3mikOPTnzfqM2Sbed4I4a542snmZdO4aUBKMOexSwwlwgPz1
oHz7S+1gwOJB6RPwlinWWYhB3SIaUFblpt7t9nVzxPWb0ui7q1GpyHMvBbgCZrzw
7XghGM2xQ0O87IKrIcIDetb6qN6OjJsvKHZw+UdTjzwJmloTv8Uy1d2SeUFw1ZXk
wOuV879SdHj4Z/nNeD7RPSuWhSRGNm9EnGypp3SQ7YsgG6VODmIuQtoi/ap1GCH6
PG0uDh+yHU8guvvV7stzTXoni/TJshUarsxQC6S+8jqsaUHOTgsMxwY3PU+hrq4M
Iy4YaTehQ8VVGN88P8eMnfEO4+vOCuwzT4TLhrMBQk6ybtkoHypv2SJfQ8AQLZ19
CCvYEBxduDUnYMBrMEDkcDwHou9uUYmWlBE0fI4R7aZTRGr1nGUKIMlbAmbj2l10
VytkFYeJv+eOzFJnT20C0bZI1o9YVvLw98kiWhlfBHzAOwg0UAABUuWiO36qx+9H
vrWyTNAQ9UNt2H4whCxlfNrb+ZMoXRCtUSGwdvrLKFh4eJOtO6gC4jLDxUGNorwW
BS0H/IJ06YE1L8SoJHWdJMxxB+3CpPQ6heNOrhZBdl8UOM4lPuyXHRCT47bIVv/9
gDAErjWV1wuWefepMGjuRLmPHq1VNF0l710dihQHA9F2+fL2raDw/keY/sdZnXjQ
aw/SqWbMoVDXd4WHToqGxLOgVhXAC+2Hsw3wVlXGIIAnxNChoXX7VVcyrAh0oMXp
K5WIN8ee/Y+k7VWAn/feFjeaqRQyY1SV/E4yUTcN70xI553SNVfLycq8FVtIeO3g
t7ssT6JpIG4rGAUqmwsg5DGyATyItdCKSCs7/MhOsKby4eKmM/Y7407hA9C5UEE0
82XUyJ67Vvh2kE1KPY4Mhwab/TejaGj5lhkDCXeu0i5sMSRBXHD42SuXVOKQmscI
rNqJ/24Vjx5JnLjn8Ooxq7oGWJJm3bEcYZ1OMXwNHXKNUoQORQd6WWY1lOVic/FN
N5z469erOA1PVsbycKC3O0BuUyEyxClIlyziub3+6xuysW37gZk6Cx23LnT+tPEN
T3W+vOzCAYrc0luw7Hw8EED/LbS2aveiGnkAZgNouBDGXpg19n9/OGhj7kgWZ9xu
h6UzJGRzIcgBFzjDSi/gDUzvMFMtUSx7uoz/qTKTmlb5ujafeW54Z/NlFOB0s88y
y2GVnEXvRZHM+fhgb3+QdE53/Jn9sZe4eraj6RPzHSaldbcJSw2tDDv2ry1sCJmI
IVbqw8VgyQ5K31RJ5ir9ro0WOMFK34mS/4/NSGIp0+1XdFlCx7ZfJLc0u1F6AmlW
tnqaYq1G0qPwCcziYuY2TFmvkg9gE2GoqOqbEoJ7oo7hzajulrrVVAGDOanFvbwa
V/o5ASb7+pOJtwE3eFwPu+LCTnzToC97UQTBcBYyIm+w2/lHOMDWU2n8ZkoArqwh
7n0I2OsaJjDEJgQu5OAkMEqb9AESUpm4nIL6hptD6RHCXPwSVS7OvEcY/x8P43zo
475b0aR8o6DYPtVu/nT2xr1cJ0tJr+xvhgqorMiIE9bpX51xVAk2A7J52qPbXOFE
ZJRYH+6QcZjBeVfcUtBSoX2h3WnyxUcIfxpk/z37Ry45fbfMHsoJMt38NOFValy7
tmSWvzBvGfS62PPYkrSZG6nG7Y54LtWuFjo9ye8oAoANS5rs8JFYeBxZz7l4v3Xi
+5VeCUP9fXpEvSLKDuRcl9rdFHsp+4CmECD4tNNfMkVSG8gRB+BCbQCcjqL4PSIT
VWhsDdtC1yLGue1/ZqGz2bNx9yKTId3ge5yk8s3g3Tg7Xzmfmsu9k2e7/EvUKN0o
E6XKCvsv6txRKzmME+KfWEU738PQrS7+vyNTOPHzCKN25S1z3EfR3r0loYWEk6c7
nHdaYEYdsIOqeVflhdyQwn4ArhvBOm1GXzMfUHzASSLGSNNOMK0GsCm5t9FVfHp7
Zx8v1zHNHJfTf37OuMfsUpAkBmdCl4TH3h7td5TBfISgHF/yf4ytMQxtA7IdCZx9
a8dQnMd5e5QPmYxX+AstUve85YdJAMMW9YamN+h1p1r5JYIYiOXC24r5/QtyOA7x
CQUiC3ps+mRAkP9anaiiSYYgH3D097PDw1K+t6bb5PmblnB4bWG7/WWvdrkDYTPW
Vix2R5MJ1+zTsGnVMZB02hAd3zyGv0G7WMs7i4bVLkwaONMxBEzTYzAgPJ9sqH7d
9H6azWDglddy3+uo34T/I0usRia2JoeNlNp++Q5o4k6X9hmnlPKZyp39SpnPI5Qv
fWxgzjlLEfnM8dJsswSfYCyjuYR+xrF5yPWEMM+IQDBUYiaivOgigcoqIj6pgvsp
ZvrKjcR2IuiarBGA35LoLYkUSj9oeUrOjKl3xTCYMeeN1vgCgy4FUDCLmvmnJzOt
CV9al6qQ1zzyJGXHIk9HAoV1+3JhwGhocrfeMkkuiS1aq4NdET+2zyFpdvkCRxSd
xNjKi9u91PjvEfKvBajwl3V7su9NKa2nNWZjTBLnc4MX17cJP1HK+xsDFiQpFYJJ
LQcXAm6W27cDkpXJjE2WTFILdUxq8g8Zdl+23NwFD1njb3N4y1ZZ/22RQ4I8CP0v
CH1pYJQAUIiYR5swdr9XYXqVQwh4H3Jne1FAdeTNiaNw1AxHGcC84rxS9liAg3vT
3yWu7KVrknY0lCgu3nCvcQi3LnvNT+Xkzy+3ukulr8Rr81LKxmt7XNA46kjUrjc0
8PRiMcfjSVMVmRNxWy7RBLAOv9ZQhvgU6zSp/Rq1XVhNlP+DkY0n7suOSWXCNOHx
DUtoDpyQdmfrLmoDvQ52b7mFdKAhRhX+0ydp1BNGrtIRCivXmnxGgRIYMSSfAR6l
1bMYZ0r9lKU9AzG54QDgkhQRKKe+c8KJiXRuBSlx9fDZ63TH66wsCpgbO/igHbSc
d+eYa2Tn3U1guKKJeRWrOpOS/uqoezqj0J4R2DkmWADuDfBYxZPSW9aWWcp0R3xI
YVnY4R191mYW470a+9Tjc1deeItG+A/X+Tc+O5hfWKRT5TnMo4xHB6dDgxVJUNTs
EFi9e/Xnr4Zwp6b6/jyLvtk5e96MByv7XBgGTRSbA4/dDWsjmLvV70unYAIX1zAT
INQv12XloIZNLNjhX1W6R/J4cIyib8O8DiDYXcrvid9Yb7LtksVV9LGGIRLubQMk
NVUXFKtiBiyrdP9/lsg9x7i/qwYu86tn8daSrxL2/LthySp9Iv2UHglA1on1Nv/U
OwBeakborAYJMMbqOYIKsHpu/P+8uLR8zqoTOhfiqDvFI3mmmmrIE23JX0giWW/r
lV4Q0ZGdDNyrZTFW2rIJXrYKGkhsmixEXicSM/9VrwfjCfZZQKOg0v6OdlXi8pJ4
YDMZPoBRevDrsd9V0N/ri8niA1mr4KRhV6gcP0xNqBjRjzM6OvkYL5SC4LqF68P6
+svQGCJ6FGO0F3KgT0SbLX1gze2ihwUGixDPKkWO/XaYhB9ATbihuZWv9lXa2f6H
9MpS0N8miPh3F+xcnYCeKcaG+gpDRi9FR4MtbWPpLfpdt4aMRINdQEX1AM3vRCs2
nMShdQI+vtLRgbTE7vR1JzytuNPibjVZPb18nT8rG3Wiwxw9a09aM9SX3bBIcnLg
CAPvk0zCeAefcyvnJob+wywaxm0XP3Pe/49Tw15KUXRtD+cjzJ+gFd0MIdYE5GLG
Kc4nhtjGtNW9xwmq0SAEldZEPkB8MRM5GKLEGWFHMDHBscWFmz7eXMs3yhwgKntx
A159AKm4tULmXFNTXb4t2Kc35Q2107p0c6Sku9CVO20bbC8a3UAFsdZXMG1fnV6t
d2B1gpKsqVUsSNvDdwwmxr0yZgfNXRAWXEYtfCbxlFcRdHiX/1VfT0YDvDnmhuKw
zqxWxgfTkE4ph/mZ6Jg14yMiHt1fnG6V5cWsDu/zAYN1EFSYzh+70Y+cCgzyQlgO
yTAG0SnYgp9TIXodvT1l1UeO/DMxHmjW66u7x7baPgysLt+eHpPqQIbgDChmwao5
fmCxC+Y9xPNVirm3ge3xy4g4oymVlHnk77oHQfk1Xn3USM4hKmRf9a7rHmeFNd+m
3TO9rLVLbiKe2XXTdOglOhROJixZ/T5ILfb58iJcKeXek63V548ms9nhLSewQWYG
afg9t7qeLZGQQ02G6eANi3Uv7ZWrw3wbXmSTSj++uf9hR+MKhsTFCDJkh25o9skX
YKZBRS4+tkRMhI/YA9NXq2m3LKaG/br6qlABQhZilsZS8jZLYBEUhwoB0aCkyRbO
i+2G6L1cznzOEGKsQWoC+iroTFIgdYFDFdLsb4Qd8yExd5k5R5zhbrn9sLooI0PB
lGvPWlc803PPoNtdMZqH/65AEIPRJFy9elfEmFQmChN8fzp0UHViA7xYlumTYAx5
WGZ7G5+O3Xi/2ZGON8OV01FEz0WOCG8P5o9CSUW+kO0wDRJzmKw8bbr18X0Padi3
fhMdGoh3x9DWcaSS3Fneh/ByLpRZCNcQUwf4GoWqaHTFn1ZYUgIZtCOLECw5gfg7
oKUo7YJJAxHkQj/0LkMjl2RBupUOw2r0sajzSrQgrTwU0ygbQHU/NsfVIZQekbBj
SLcsiyK1KYoDLgCVq6f15lwF7kVMwnFhvLhp47jikOZcnQ1N5ckr8jHkmgWKCD7e
GP3inYzb/qbB3t1gNNrMxtRaRiqH53JlgubRCCk6hwbhOsayWygrEaMfT1X6KEwC
dI9ir+f6RbgwCATHJ0Kwm/Lpk0wCFkL9guTAZLw071WT15UzZI8zORxEdq2DyyDI
b6SvVf4bX8Q3VhrfgzoWS0h0HJsbKayWG64bQwlWC22ztD5p/t1jldYgU+TCBXih
GF7qQZzDPBiCLhJCAnxwDck/ksKKkUy+ZlT/dxPodGSsmB9Dfs44kTI7ooPRZxjR
hFCUqW9JukOCaBDzbwurXa7BMBwyrBPdXoSySAepqcWZZzbH5oO9bR449XaWnO8o
zXym23dn6ygYYeckfgVanXTaq3czs1wia2AKTkHpL/vCmkjyyqm3YFzVLq1vV0xm
fuEaTvvgNefYV0QppGmK4NDVAoxosBrEoBXhak6s3DLO3Gc2g+Espttmjy338JZq
SNWnuB3z41M9MqhD9at6kQhZzph2wNVMBVpN0NjS9RrApo72qdTiycXF7oC+tcPA
pzyes9EZsdPlMnquQwu05m3DHLh/liOR9z5x5v6M4SN1itGzd0mEhfw0syXdZz+0
j8CZKsgPd+CFjOv+n2g1yoFxEei96ir3KtkcgQaiVxC+zxoYVJBG2Qwto1jhbNgK
lgozvTRp9Fyq3OyoBLsL0nNdSFfjo15FzTXEf7bwJYLme028I5DCHbAHEpQZNhWX
0v4gluW6Orr2T74m6su9vX/YWpePodDEH9hiAgFWXXMQ1xIZNIqsIhkKlcZ2cTDo
Xy9L0f6FOEpjQ+tkyjnb48cVJ5x/FB7u1DkY4Skwazce7OgKvz0ORYUedvlp6FRw
gTc3DYuZrn0tAUGmBXtOEAd5hHOp7o4lyKdXUlnFXjBkz5STr8xBf+1/cCYR/sBV
Fq7qE7gKao4nfPszHVsJ/jKTQUji+HfLHwcnViiV9XTIWXUcPF74klyg98ERwTNU
kCfsOiAR6V9RRqP33Nqu/U5tO7PFaLZd1xp+MQsPZM2E+pd0ToIDs3OI4U68Q5t/
o16oyfpmO31gKTnux+xF6ocUxcOiPd5LJzom/ruEf8L0qb3tm5W1tYT/C8O5aLvb
RpPP9w3Z6W+K97KNWUi5jwM99ZkcXzqhIRPHvcuYShDerZTo9KsTXwT/JSyYCvz6
nJgRnnuMtega4ssmIJwPStLM09w10tCncAYQMBEk9rloOrtiht8kzu4h3wseGAFm
72zFRQfzY8BTJyWWFfe/WKU1kjqmODHe+hEQ2MGdV58PNFSdrmc5udHpFYjzBLU+
fzuXZUkl2TxwecCkoiGwXsE7JkoA5aWWpMUZ2kC4T4B4puX+vNYBdyWTWpf3Gxqe
pVEue2mn6tf9Wps+S8rgepddL61oeTbrqer8TH3XJypUJSHd6ek4L0bNpe5cs+RT
jw/A1ZnizLGSqRJzdNXJRYkMIOkxTEkNqwGa5v4aAzjnzfhg6G2DWCjftkU51NAW
zZO/D8mTWSmEjP9yGxfoYjHzuWR+x2LXoooNdyJo+Rg2As03I+rdELIscdMw8aYw
By1Ya0zZb3DBYIVt7i1mlT7GB1I8vtgRr4W55KvYZezSMdELTjtEVoMoxlDlnm4Y
twaUtxqUKwv/QrsudryG2Qjz7mBjrbSe/asMHfIDOyLLbgaWoMBd9u4xiUyULm2X
OB2CUvGCZwP+cX+BMaSQVb7m2UCASb1GrycDZme4J6dBQtngm6ItOPlzW+Y0qtkD
rdINXbquDrx/sLPmSz0SuuNNmHCUO5N678WQ6734JcSqHE7ddVD/cBHUkXiRtauj
s+eyoyswOPURCXD0acWb3S9ixr/15J4BvEezurX0+9D+11C/nkZuU65DHb182TCu
lauJ+L8Wz2IpkG/dQ/5VlU0KX4ylOsqnDW3oWgCSKq+q4see/6F5nIOFNejPQuTP
VA8zALkJbDSU19kJidOUhQDD85YV7+Wp+dX+choaC2BtHcYi5X9LQ7970lVtyiST
thTQCs9S6yx9FcvAceyhGHpra+E29MaMWQsE6zqYHPalU5UmMrmlMHMj9Ga+BtYX
kYl3wWdo25TSWgjjpmFT3B3/wmef1Xx5RsZBzIya424mW1qUxGRZA8TweybjHOwD
ycOCEJYmx4TyYuXpOXrhu0ZwDcv9XGjpCrij6EVOSYQDUfj7+786g7c5APd/td21
8+EBpipQyVXqnk9LILOX1De0Dc7Jml55yQ2o20z6pcXLaJOFmTzXG7wr1cYbwhtY
Qr3RYzVjYnZWh8RLZeHvRYEI4f1fk8nS66XjNqp8zLHIO5KSbNyvLBI+bqHkEf1h
xcZFvnALpvhygVkdmctj1FRPNhz+dbQc/YSUUCpxd1bibatakD0APHunCoMnk71s
yRy3jpDVJOoRBFbVz+wzW3N+UzhhA8tQP0hmkru5SgshLNDfTnA5rW8ZtaKKYGB2
O+RlHNvpA+xtwLmhznmClKWHYqSHosZDsjNXmcCW2FlaTL77qUFR3hrCok/6WkLj
+IU+xYpfeglBtLV3DKZGhXwOAM0hcMiSnXnH3W4HW/EIZ3LPzLHdmkePLbk1zolq
4E0ItEggIn8iNUPaQsRm9PWxl2Of1nlpfVoQ7m8i8OVLh/mpxMKGH6JfApidtV13
DHayDlKee6jsnghW6DJvLLq/v+XMzpocAPmCpIz72CXRwulgFEmTgzE+8Mfi+dgn
6UMNiOopXrAlUdvmx8sDL3z92RRvQ5IW4aMcrbQmERx1R9vAU3UQ9TzXDRXvF3Z1
Q2y4DbgT3SWrxnVY54teA1H93qy4clTWXQz7XR/R5c+/7truLDbgXHdH5f3GI5LN
ckpkVB4iiToabkvF8uKXVkpgDV7rk4/NNCVUEdAE/uppeA5uqV8mkAV6CHXkhBmW
sWNkAOUUIsRbcYuh4I9GVu6bOlFfsKlTPo2qSfzhaneEscYAxeoTJwjx7UM4AaWd
ftiUYn6t4+P9Ljzf2y48YMwdjJs+gCbnHlWRg5WZL/GSHY/BBhyHv/VtPH93fGUW
yngurlcJjrGH4zpRK8/RmborZn/bsWHEoqxRbLw7C4rO9VtTzxyZGwhQdX7NdVPR
Pn+ojPmwklGYaOPlCD4erFSI2apu8NDzPqOVrq9WKACFK5XxME51zeY/4lHydlnf
yVCnvnusm5xlNeIU2/xfcnSw0vrCdwFbH8Lvbei+Tfq89GWLud97XNclBHAfyfwc
1qCPVF9ZUDfncyAiNUWDlZ4BJ4Vo6pg2fw/IhAFJlkCf6wkMq6IsJnyKNhB0p2Cx
QsW7MnQf6g1osr61kbzvQuG9LQmK4EQS23Hh/vDxm1yG6AWxNO35UHBl5ppp1Fap
2l/nX1nFyfZa08hBBfAHB9yitTB8vg33I9LYQ2cnTDdjnY+kpw/iCBAAT17Ea8qT
sZlup3GCLP57fBpYS2dlxMRxgWVexlaYz8QC6eYQRS036Mx5Xsx68lVUR0vzV+pU
OFKvuRdjogkk3aFsNjCuz3H/p0P0ozPruPZoskEsDPdwl6hpeEZzRcrBuvPvyBKY
juK33Mjxi/agLUgw/20GMpmqLVJ6MAToYktUgiV7y5ugIV4P0faP3HHwIrNCu2mm
M5rOf9iyefq3tAQoCYTzntu0YR05opE0553q/KISDuo5ltk3gYssMujQ2ouy1SM9
4IuCDbHbWamKVqooYS9dTFxF71+PLL3ZN/MvoIlRkVXKk9m0OhxY4e6Z7Wc2yrkK
M9m7SIJfvl8MrcfgUDImYBt+VCBIkn/pmta0vbwtGDWTE/IwIx/pIL7XxywOkbSf
4u73Zp6sLU/e6qNaQQeBlBZVCFRbY7a+0K+PQCpZsf6zQk67hyyELVa58ukY+z66
eelS56DS5WN8pxT8SgV2P43HexeJExlFbY4TbegBc6FmYopThXLbHTs+oXvBHe7i
62TBBiC1da592oRTTH1hSDE/jEmXgDwldgDanMKSt4UO7WL/0pqTdPxYovFQgEeF
Sn3ieAGpVs1J20j8JqLk1iAy8eXgEApsVuPXrMEj5Bgm5nC3twUQOWyfSOCdCnJ7
+AKdfNDkoC9qoxFr5vjXwUTBMMXTJX7C8M4Mcg3S+mjWy77crKZoz/NBGWO23PtY
qnoE4/Q4N77ktsJ9JJrb6S3qx1Si8ISXCkhhqSY3dvM6vgKMRQjfk/TK5WS3goMA
4rxPd/ky5WG/Qlv+R12LbH10MuFcFkXt49EJuy+UlxO4GrGk+/GqojSM4GTq4r81
Zg/EREcvywgxeC9oH1KgPX/LXAbA/9xeOQ4GLshI2Ht2MVFCm3SrSk9X+SUszmbm
LbMKijEDoD/IO7gCAF/KzAxzeXikEXLdFTnVbw4IixWUYPed9yF0NkyV12W7ma1v
BVGZf3UCMlxIQEVKnNMX0rqdshUfsbRUpR23AY3VOy4AFPallviJO8qMt+78Y5I5
AUv+5wdoPzUZET+6xgFIX3sjOeWooYPTYBWTZmIeRZLdzyVrGrET6t3wm47BkwvY
0vlMFz/yRKWR6kl+gdKdWmW3tCYuMVYu63dPIPIb+xbZ6giHOo8HcQ9o+po2WtPY
/K72dxebwYaZFQKqYR8NpYQziArwn5Vhwf6JmkXNbHrECnPpTwWInucNe2ND0+HQ
gVNV7vh3kiYOLUbIX6pmBTS7KOrGRF5EqZyOVPKwq8bL3KW3CDcgt6XtlzCjTROC
lBvxrDh5cEgWIfrxwQK6YK0qdP8kSh/tCeLyd25hDGL2+DYTFfGufFOtvlBU0C/F
aKdUSXqJJqyXKSi8Ytt5AMkQYjTcnnSYOnCR7TEjOPaGUzGggyeIKug4y3vMMVV5
HljaDX6SQWbtAMlZiM0kdJ+uWsKEbCmnXrsquJ3srkLV5hk5t9e88be8k3Irjwwu
2tZokx4zAwaUdJcumZmJnFth/K+B+utEW6ubDd7ZIXii6Nh14u7mXEqiS/7HirpI
QDf1cGkh7y8jUOyGvJMQa5eQikWOtuzB9uecj68js6KC0PBydkehK9A/lwYNjaV0
dzl7CVXF77bD4ydkOK9fl5b78iWKpsdzsUsjceVzsymkpWIOnRKOe2X6wRraTcIE
ic/+ui0jXHopvbsN21BkbRZrTIgbUlY5wkwsGJnAP/14SWb+iB/cCAzeHS5fcoOq
0usswgqM0sTBq4rrWkwOYl/QkpHyrkuEHU4sK8UsPlmddSRWwDIgTj7SLv/0yh7I
mslicxxLEbh4APV4BnYGKDAwxqHbGkD+gAUJ8LZMK2Bk+Kh4omT5shvLeRWsahN+
USzR5e1OZQ2GCJPOAo8U+v5zs1hgo0wfL86VRp2xyLEz2cszSZxq+/MujYOi4EXg
Y2beF/3qN4n/wIoymp8K6r/AvOkYIlbv2bZYUWflKR/jlgqYWqa3TzWQ9ZtwaArf
nObH9TMBByUpBK8Xl3ac8R/gnIrs4C+hX0NyLGjIvFhSlgy+h4jXor3M0lv42riR
ymMlPJ826XfLPb5x01Mk2Dvc7GPa7sG1QdBJ2wjG5m5H8JetXoVheZuEcgfWZ5pT
BFfxSqoqoxijgDJ/EPwJ4rVVJJORFMeg9mkwcSCM395vQHFyqO6vPTrVxv/el+kU
oDrzoZxc+mw5ukkyfIoSZ217mIl2oTNSto6gaUeu9VLzgYVm9pNOduTRO8/qOES+
vVX8vTSj1Qc8opT01blBE3xWDNz7372igB1alQHi62iqgjPfb412bI7pD5W6aasm
F5q5i9iV1uBfSAkkB2mRAa6ufWGJ471ChUBmqh4Guzq6G1Vp/sj2N/gTXwpdi5Mh
3haBN1SwBA2qF1Yj0e7gI6NnImZsmm0pDfYlbQ3KzrMn1Dq/+lurPrzsymaGwdLh
PpCaTofpaALRjEK/Y+mxCiwO4ycS6EwywcHbc675DLW0u31+9zK9aubgUzjnIiwH
nsQ+y9dPcr5aQFv+BFZtwsSQc7qkD/782vtsfuMkob/9gokTjZY+ht59OywS8oOU
jmtzxf/6cuetczSi/PCXrMVyGYRjem2ZuWN5IzkvQW6EZlmX6CrvstJXcbaGyiVv
lXIYOs6xVItCuv4VZWcUfVjXr7UKQIhOP/tM87a9P5Rww6vAqKb374LGbtZJ1ftS
WEhy4qiS3/EhOsEgqeo9b7OQRZ9uOuVXprqssjn4YSxQbGuDPNT6DPPvmHGJdBb+
7wNmykovRnxn0n+oF247aIp3ywwtbbfr6sDsgGG4g6JcVMHLTqqPqfHnUwH44Fj1
WGtQON4kkjOdSbhePUp4MMvXOl3wzreKTuu6Khmc9HZ2Q10S/wSLutX2PrgPDITQ
oYxpSurlsKkKTZiz3P4/qAqCZ9JEBKRAqpD+9HRhx6O58KusQhb6LGjOnTsGXwp2
jwVdZhVroP/w5OyM/PPmrQCczA6DlOKeRxdRSrxwGrRStHv0vrRf0IPtluBIHsr6
0o3stReMEW+NxPYTg7jsXKxKfJoXc5Sj8SekKQKBjgaF5Zee0AqEfjOFGcy0wmYp
BJKjJy/QR/oE4/hu9tAhrI9/Q19oZMXEcSZnx+Ob3EHZpBW0VqjoA/IwEaRmOuc8
V05DgZy3BvQw+2fG+KIRiVjFgOdcE3gDbrzSymgDSykAwUQMF99UXBZgmBvmK202
urFFkFEZBIge/F/IEqEApDYlUuO33MPiidvzSuk7nA/WOtp1RkokNL7oe8CpEVPR
LnNHkgOB8HlODNA/vx2qDBltfLniVY2taUkawHHvJWKJ7l5ZluRRfzMhg3/ofHnZ
rKNTYSSbL2SEVNwqrMC/9UzV0kvth/hvORLVo5bSfZqQI8dJPMvK2QJrNAMfbwQb
lgBXyb5jZfhfqwkXrcAKgVMAm0MPG16K/kTj/nQUkV6qM99g0wGT5ZpvodODwcEj
NSE0A9ifYredRWdZ83gbMn0Y8G+xeYd+RHVwjG1So3Thwq1xIO7mPxhgEiIBsTn6
yYQVhDwD1k2kRmE44fbbgwoJ6LJ7aipxkiIAX3RnP0fbjLJVHjcnojERl3TKruTS
qH2kwvdaQD2qYmDy8Eds5KTcYnBYYl6dVVRSMcex0q9xQoOngwrY6Ry91qgVhFhi
2wcNsXeURy5hA2X8M0+QFyGv5lVljnd47X/tqTb/rlBWc1ErByB3J//13PB4VSiJ
pWHTQYERV3dCGAdfBq5y5NvQf1QbhvvTBApDl9zLJETIGdqz7L8jNhrYu2FinSfq
BWpOK8hC2E3nbHpPpWYUniLUYFIRgo96nVrupq8lxGXflhmyX7VYAQZILpNg0N/z
0b9Hs9abiwD6G9VFzJVVqWyR7gYoLqIHxf/EmEefxBsLEdy0+vlVj6banOEkQ6hL
RgeKwMwB37PTI0QT0RtnM/xV/iwb/LOBu5iKS4qvafTE6cdcq7/C/piiAXwlEUVl
1XI6ta/u6yLVOWvv2lxHyrlEdcz3mZAzyqsUq4Z7Pv60BywMiFFEcQRvhMH/fvdG
QcbhqvaWSTHJ3UI3qvz9rgf/WWeFB7m4iJ10thAhsZKnZGDr4+SBuJSp5zio8LAE
ZCSZE7AbY8n2a7ommFZuM0ROSM4L8tBhtpif5e0oAWfMC7f2ym7XSf/+Jfnl29i7
bgzZ9ONrJB166f9NMl55JOg5ipyy2sxLbPxO06laa6N3RI5N7FXJiSuW+jYmpn57
2R7Bj3I7IkErn2aaulaILvcdltRB5aqsw/tARQgzRI8PYD7Vn+8ctT3HVg+pPxep
sO7mRrmuJZgu8WFk8kscpMV9xvi0bFkEDGWBxLu5P1k/CmEXbkTHbHhHNXyYtfJ1
HgUEiLJGsZeYOSvNHft0xO4w0j3emao1pWeO28PWkyAitnQhz9p6Yu3MVqvG/Xz8
yrFT+x566Ywy0SwZvhoBaMdxV/dN74pndo/M4kXYB8vrYh09GitLDzftiQxi0jW/
S50ZZhhHeC0WKL94DaCqT0t3VSoyWhk1FrDF5Ni2ZpbDPmc/qaTPFXWp2nO05bAn
eou2ZEoBTNZH+R5xurQr1XW0JUs6aiRVpP0pHX0PoIUU7J5uhcpqjt6o3D7aZ3pK
7kgxvwnGmkrij6JiPkQ6EFfLS2hNHthJlhmwo6uVKlPrW2S1iE6vsKoqXc57C1WL
qn64kGkr8+H/yB3JeHR45vQJwgd99mWUqul/+kWImRivaIvJ1j1NBY2kCCiGlW3u
pDrAFAWOxwtP0/4F4nBWJKp4r9ekY5UCa9nNLulGrkz7eNnWu/gqamCvT+hQGVcp
09/gVZI5QzDEZebfx5BIUl5BnHUXyvF6vdiuBO3aEFp4+r4D9ZaQ7f57PvNMU4+h
N2dj+tWm+3xDKKm9As5W8QtxaEw6jq8TtRoPG+QYl2elEp9S6ymigFQ52/pSkjjS
sHkYzQ/ATzExpst8+olNDCtLKfIOTfOcciRQwUmSTS44uHxAL86S+RPVh44qUaeD
Vq6deZmRYWA3zjeNOBNKeoj8oEbhJx+7eC8IpNz+agc+Y7rKcTnA9JRFVy20qnT2
VTIUId/Ywisp6VNuiQFhtaKkalNG5EkOkHUJOxPH4RzfoZ960FocLQjUBuTn1lbY
ZowTHnaqbycVsDCkvC5R6NEFIrLIAZgKiAQQKH9qFHZZYctGeGfo5yN/mkBDOsmg
6tCJiomiEGl6guAJ6zZkFtOqV3CwwqvHoqjPf17TWtp5ZNIMviEMvyb2zs+XuFKS
ixxDHGtuSfdyzRO6WWfHK37IV0UP4ac4L/jpv+0QmlMMLl1VEtLCg86dJlG6HHu8
y92afnZ66D81VzXDlbQbz5/09RWuLnktR3rFviasUqADAj0x6b+lStNmGyoGQ/r1
SR9+1lOSEuOil2N9G7rAGUA8Bm6FlpX4dH4cfLOR832RlMMCzwrOrC2Ak5hhwxvp
/hQ80NxFp5aq1rWbcqXRqG5TuCmR08TjK1LMjKn1MI8lJpW1p32a6+Lkk2GcNKBj
3mpaAwGNQAxImrhbRHeU2uUvCQj/v0/lHHBoT/M9KHlx/7wqOBdmQ2k0wDwdi6YY
Ls7pvmLNKNDuGd2Vrdft9tPi8OVr3O1Gw4pQpHYeLEDY0LTTNMGOI0UwKOK9BoFW
UqTsVf/f5uX2Km0Si/CTSCJtsV/ijUtgYhBB/WN/vsdy2I9AE+b/uATAd1GIwCMj
nQQgV5RC/NuQ1GeBYG55ieF/GmzqY1tjR64T57bZAA6j0KnU3dvO5E9Uk3tc8kNm
GaI2KAUVkP/V+9Q/iLbVzC8M55ZAFLA92TFQ4qEthDACH0+0sV+ZAokOdsisyK2L
qBtMxtwkMBkjYzO612TNkxpIVdAC3DHpvOUta4m1pfjEJTQKj0PCZOTDkJhLxKLj
ksNuzg5YgzK9YcaDzEND4M9o4Srsf/z6tCICe0B38xujTLmXbxfOdzXTgS2Rjqyw
9dZd48fLSuta6ourlckBqcHm3DY85kQjrrbhe3qf/ofg7M430noEG3Bdd64bgCix
ABaguUx/on4EUFGc19UVQ/w9DhqnQOl2XEpqZgypBR2cGQtKZbmtWig4gMy3J7rl
TzswArTCfLvS2q85pZTKsI6MYv3HGf9lbKyqb77SZ0rL296Y0K2C/Dckls5MD8wO
X0j6rb5oFvp0bDAPdiHiJJ7l+gZ1+439YkmUdS0w4w7Uaiqrqx/gBZyn0e+Ad0cK
mvyvi6LHfTexTODWQ/wPbGA83ofq6B6WJfXj/UmnLh99V8N+y6drRop6VCf067bB
V6FdxfChVkBI3guocYAZcYJV5tlPqb7j/E3EW9kQqMYQt6u0bNRMnNW0zfS7dG/D
uzU7qEzTPP3UhFmMTYOk8/iyNCu7ulaWlfPe2RTTU3eU+9hwzjwA+Oot1Ki7BdOl
7amCTJhDje1RPO5CpVyVlF6qqWWhfcu+CieadWAoH8u5WQwfoZCzuoax4K0cNAcD
qUll298DPEs0T+GeuHgj6SvwIwC31RL/C7PWsMTix6KyIsMiaAuAkQfuZLqHr8H4
WSeYHpcg7RTWVGL90XFFp23vfXQdQ0KUaN5Xj07wFRANXvnX4HVe8YqXxQ5/XOu7
ijJkxq0IjQ3dCoWQ3QZZGtgMwdZI6ogvcMV02d0diTliSgkv9zIX8ZsiNUSDk/o0
R7Z10iydc16OdOj9E3KWPNXnmjzj3HkGz/2fzD1EMqYR0wK+CL09sMZBOP04tpeJ
f84m/BaHQqeuwUNFiVMBBKGSMX3yOcdSddaS0UlH7z+zY4Y9ODogJteRjc4H7dBW
MYaLxVQ3YfSFGikC0Ahcfa1TCg089hCN+e9R2L+S0OeRu/vMLvzypQoynFBRS3+d
DZBFCzCa5fJC7rvVOg2UULJbfiba09qaqZWeIzj4WXBP2GaHg6EWzxLJexwPEVBf
xY5xtSO88XGj4lxzsT2V9ePhOdUYJWoj1AELSkolmGDxLFF2u+Wcjn1l4/bH/NyA
e2ZGwAAFlKPoy14qmnJfQSeYf1jE4VLdEt8ZcLaUWhrTUJEADu0ELnhattyCp+4g
AyBPgwJreD43lttFfSISGcwfnwztA8JxUhdMx9sSVYiVhyEQVNGKRxN5mrxZUv7f
z4tgnVEFX1Vuekb5zkumFTEn0r5DQ5+Pl+ObhzNVQUcTZX3dX5QLkX4LUP86a/az
g2YM7IuwBrc+PZYXu8Ik8H2bQN4gcpGhZgm+xtLQUefSi1efiC9WGFFx/eholKT0
Tbk6RBWvLnRAR/noVTLq/XMkyM1zvbQKDjy/iAW/FjJNsFPHx3JpB8lqYJaf5BtK
Stzi0VXwkCt6WlNP6dIG/WJMgjtsG2fuqHvHXhYDsxSGnr3xA+IQopseclYnTdWb
EoP7fNJGxxv/B0vCRP4TcrZIRTSwkBQBDY2wDYXdxvtJ8m+gyDG20F0G5bG5oZYc
/kWCBqLw50DP//tyMKvFGikG7AdIH+6yjWdw/BdoxvjOuqO0db1PvJmrSaAFuMuP
fDwqK3qSM7LhBcNqyRrNss5OgUeDs92C3ZIqAewVPE33FJ9hkwo5TCmsLl/yohg4
BP56n7fhB9pon9ZNxJPkPaKJeBnyZgm6axtEidyZeCibValtYCvZKyZd159KPNVQ
gs2px0Q6WgWR3d+CBhNK7eZMsa87gnl7Gzi+ueIcPcDFWr20HKHjsKt8ujuVUb+J
lZRKmDKsC7+UnkS3qXB0Yejxje0aY6HL3X4oBIObgFHlfY+PzVklHIvxhSAXMIOi
PtaC5DWYu8jI71Z1GXJOxyOZyL0u4PgHg8lyljTvPyVMDxToFJ+bY5/0g0znXWHf
cXhpXZBxlKLblnhOVLvELzxKSDHURQq/XdhXznHvnRAenpqz6mpamujf93f9eT6B
7DMU9tZ9ABrSQBlyKTrsXklDiQd5s+sruoTZG3hJSr+uWz6w3x8scav9yeasIIYq
8GDMeL5FDaiuXZh1J3wDQPaV11KaXz9BpyLBhVUYf6tRPbxQa5v1qy/Y2UgzXXRU
bcy1hKNaWOJHNxQN9KVe9FXejT68LHGuy4wVtUJ8M1Wzs6N3UUCp+G1QXY07SbNy
/EHMR65YpuwQkO8aAF7NwjKryjJDND8ssJPnTMMkbeCgmfphvcjB5qgAITd3BGF0
iSFYEI8IZdr9H4kdD8wmsTgeF8/BUCsen/biQiqRIrgPWnXwrS96IlsZ7Nrj9sSh
7fB64M+wdgyAjjJqXU3Ahr8rTrbqXrQRzdB7XI+8B8y12PzvH+sN470ervuiwRxR
jwh4Am4buZ+XgT7L+QkgCSmSRaPSFT38OkOFWeeAE2VBPwfBMZK2x2BnFy2kVYbV
YYvcScaLLOXNEHGAw5qjaAeahM9aq8QgcH1E3Ci3WgaRTNOkNnIztrUEqQ5bq1pA
4oMsM63ZbSGvULOamK5a8EksFzDPolupOFOF9wilUPtWQ2ZjcQb/ZJE6Gl8USJj0
9rfPTDF41HJj3cshapYXty0E9Gv1s+Q5jjK2pUiSQv7KR/bi2Mlen3T4stPSTPLb
Q0lHFwl6ircqZz3RCQvuU1Ys0u+cEILudcyI8rwtRrgudGhtQElq3RLEaGSke0yk
J/Aok22hU384P9d2cSHXxOMBki9K4tHGF83gpK8hwwTsnLRL6Rb9jLvGXuO+VW5X
HN3YsAs+oZnZ4wxyqUSr+BFwGBLlcZCDQWiBvblDRKGLbCdsbyIDzmmQF0Qv5h5P
gJ1zKCGjz4ZSM/V5QBBgFb9OWFssTychH9yQg+VxqD8jZGWU8hdg0HJylRy/bJIf
GDuwaW6lq0MHjcP9bZZHuGzXp0QGfDMnWGXsWrSnuqkqsJsfXew6v0BSZRJD/LEz
VzMR+zcoMDmhc3Me+qaP4JH8nMk2t5b/upuzQQo5nV3I1NZ1I0gFmdefgFmzKi7j
JBAGclOoRYshJUjfHA3AXVegp+JgsEJucpI4+9zITSsggpbFA+QqUKVKIE5stOPm
oZeaQ5Vlr6FZXFBAkhDFiIbdodsOF7/1uzMqdEhc9eYqvlKrS+fxMp6GkQ9wPTen
UFF74Bz8/soE/jDSWIY5KS1PRQw1SwShmT/NX1SNcD6ShlE04csQcWhDR6bXuEi7
pPU7WpHRXRXpz8HBBaZ5sbia7Nc3gLTg0IYrZSe38oOvZX9YTYOYB1Q2HAUh/Wgf
x1kTlXdVhV56hmbTm8vWlCuZ/B6E8ljFGZUwdW/tiMvTJtp3QpMZCSTMVX5pI+be
tXVTepTk2+Ywtwop8sWqyHVxhiMg6a3fHoTS8VfkKCLfFBD/7rYycm6Ad+6XAoRf
en9YEGlmQh3NaaNnrhJJqH5dxGJGgubXcOVUK9+X5oHXaHja9DW912gegmRAEnbu
sDyiKYSoicN4A789XHLi5Ji3eRdJGRwTqFRWzOo/k47QnLc684NmO3g2+D+1NSiW
2xf+1EA5Cxdx5JtkFidX4I/zW8TlcljrIs+inmY4schUQ4tXQOR6pD2sNmfrKhgW
h5ha1/4rUAS7+ZqU/4OSgJJ4vxS7LNCtAUXHUe8suT3iVhcOHLtu/XBnMwUGiN92
9cJ55ZsAF/oOfGHL9IY9/eTrZDOdjkj2F9tfSydEBRSvvZWaStFcVnCHtLZG7Csr
AEubBooGorm2iw+wdVmKZP3Yb1biELmv9+NC2kB354fAacI9WrlhHldVndE112dp
FlyGmlus+bYDKnGC9i+65KTXD1Qdcl73yusrvJGOodur0HGGuM3wUkgW9Z7U1Kms
SpF2NxF91uIz/UaphIqJ/H03emKM28kfq0Iao6kvzYQXJS8pR5aTI0A86VIBErnC
FMHsedT7H+OrxRCLZZ/TgZsmnFGLYSH5Ge6emJsQDfchAhHMhYyw1JiizbK+Pmn2
9WSX1p+Yz/Jmy69OnDK8K4jtNVNADUtFJgb8JO10yG2WMnDvmH+vwLRqSvT5kj9Z
d7M8FgZ7cgempXrKwthgJa+rTr8vTq2AzAP7p7hJJHAESnrfLHAaQsJYLrN+JFAP
HlJf7kU7B83tGJnlx1agQW0j60MvtFOqQ43m/CxAU/H9LZ2waemGaNaFmyyMjahA
idOp3XcwIZpc4Yfm57DZVEBjgixDtWhkF9Xz+YwX2yV9vKntuMwjMc+/4SRCHzvC
g2A1SqgW9wLKHz2dvTKoxZ4avdsnx8O+BuZ8ZTIMy+IJ+WUdqOtOlolxYlLWcrc3
EDgJ++P7ku/8PJxxAo7XCm7V2KH3EAoG9Qv0UprsXkHTZ5wOkmK3kCHovXnK/rdk
hzwnhWE/YCwLDh3YawzLySV738DVAdLmhpxsyKawfe6q8lANaf9cPN80+i2X05MP
SH8N9iVeDXovlC8WDA3YkNyiLStrXt6CwMRpIjhcwBz0ls41haG99BVdMWGJXZag
c9JgNLoZbtkyzoV15q0C1Q54sf4RjdEmG20mWF5ZQFlcHLd1FSfkDZl1frEcRcvq
2RRCzYIwQhlyZr2CX+dhKw7T0B2L1Ngatrc4Tnzm8xU/0gNCWjdffE5/p448hGeX
8kcog4oJGZ9ZwqL1c5MxsaaW59MfCcMkrqd5ZJoH+PY4BDXWzhLRBNAssj9a2gEW
tNlvNHej3OVfRn46EenSlDI/billMyRBE1zRtMYvrOVfquMhLHAfMtz4uR72Coa2
e/ixQVFQVDJTHRiCww/1rcUTqOHE7+NduksIilL/5QuEt9qy0xgxIFIjtLCkUAKl
iKIUQnfVZh2Y4wdPUuAdKvrS21GqQ5Dxa9a3IR3xtPHxKdTcgQoLaCcbP1vZZM2Z
Y20EArK0OW8u4B+XAVPs7ud2iJGU7tf8bU6X0xYAynfbaU02Y/+Qu9Alp8aBpmUm
FwTubLEniVgeHOjBusbwWygRDvHsL0itt//o0oaj54D+TLTG15e2V54/VhXlsvB1
0kKY9krPbZP77zUEi8B3RH6FBNXPNmU4e0AQh+BplrvDwkUqVmQ8awMcZdk5Ai6V
z3czCIRt8bpJkzqPBCNe3Gkukrgs4o2HKHjD6EjfOxzZ9VkQc7G/ntY/ERdU/QqI
QMF6lVszS4kIzLu7mPYb8k2U5ye7b0F0qlqCY9Y47sQ3Y7jNRTEIse/yY4hPJLWA
HVOhdJTYLB9g4LwTu5vLmUMJhnigat0oUcjvV3hj1jGXwf6MM/hvy/x2omfrCmXW
mE8pYHdFGO/BZsKbbY/YDqUB0dKswGyIX2CVb+PYSd6c2WROaWP9h3mr9/jc/gKm
8SDIok/rPJ9uVQqi58tFLgb4Y0hpnZSXYeHTAsDskY0u2Dv49NtWRO7tg6CdnOTY
78UxlnRRx0oXXVqGMzeUxN+TK39QlMsqlPpvDRgMJFZtAxe5ppNEh8aMYOJGQlC0
s/u+bJvgRbRGAyIwt9SV+MKrkjlzksEw1h3GdKCvSWYjTlC1foWfdUF7xhdxZGsY
h7etoKGRZNWfteKQeHEWrvfGtdd68T7dMfzl0bFkN9QGGKcIqKxjqOcvTUamVQ4P
zr9z6BtS2pO/OVjjRgjYarDaC0F7ldpkgua/dg9D+sBtscRi4kZbhARBzFJvFdW0
kv05jBUDl2gJ5EDQHd8tdlJt1XBnL6LIweNdEBP6MngvoRzCxeb101FHAIej8o+F
yxljxmXPkgkRn64+cK2ySK/Dptzf6lma74FX5EjiSoEA6YtmcWMAhK080UmMJEY3
4hF+3wbQxLUEXkhDWboAiLUhpOz1RAOPIQqBdCbjTAqbtom5t8WAvJY0RUBu9jXO
vTnieSjVUV1UBN8V7W/Jq/ZaCCZJ7H6hkZ4DGGW5Tf3p6EiejmZgx7aabAj/Crq/
R4oN9oBT0jjj4vN+DyODLf6XBQvzBzYfwSN3drAE++cgEsAA7u/rsh5iDmv+jSNg
zyQrfb5lDTtfRZh2+oN0SqcZRTmGkVM6GUh7yB/haqMBDDRE9S3m+Gj9a0ut131v
DXzV+ZQfIHKJWI2++hlrMbton35NNeUIM1d2cxrQ5cA4o8EID8g1a5brcgBkXxxA
eVbRXUFRhb0r7SMT9IsfI8EOVvWJDG8IodRv552eoZi/UbUNlgIRuhDBbv54gRzp
1gbdLiSEhZ000F4k0FLvkItRPIQ26rQIN1rx1dX9MP13Q8xHNSjVsuADJIUKbmq1
ca02FrXaxQtY74MrxV9NrJk2E+xhU8QPmt00Hb4sBQgYj9Lz1DvveR8se04nNnqb
P2wxwJmdLI83idkrE0XPv9ZyisOzQ2ChNzz9qNewKoredo3V0/HRwBNvYobxxK26
2qrk7tMV7Bof4FWz2GuKMBCx86YPtlvnagHc+qWgknO4lm/8kcd9kw1qrTgUmL7c
aAiL4LjsrbzfBVXAz+a3m4o7dTwr3c19pp4jty5MGcI+oA83lFnGFDOGmb7DMAO/
GPL60tVZ5HEGWOQzn7jrN9DehO4alb04Y/uF6+pTVu3wwIn3WvWBkpleSmvibOjO
/fZT7tYio3PXhqBcf2tTFoML7LpIWszVTYDS2VD/Wz+TqV3kHuOtcQRTdjzsNm0e
IiASFZifN5gxvTa5umh5HMsbidE5pJRHrf/5EMlFH3rw0NuNJeNMt+k/JHV9AtAI
Qjp5/hsc4oTtea/oUA3rvKsAIqd0KxdnyWJBt5tDiw1f96+n3yOmQ8szi/exKEzE
eG9/qhWe1vG+lZUEHD0I7lVJ7OasW8Xps3nVY8AHvjf8489wEFN/6dYJdxPSIkmG
91q4yfbxYz4QnNYZiyVRXCPnP4Xkfa2V4vCReBIvgyWkpHCdgzKPwEMGby9uOo1E
5iE/HOiOWXmM4KQyrEzclweuV9k+X2Ahj5ZkSavgQzh3/KqlE/lLd71Kl1A5auBD
exOmmeYmTsZN1oKdDaNXM32NfwTQyjvx2o0pBc6aNRLrcFsofwfoMb29DcTApP9F
kFkSVFot6OpeSkqLTAhdw4W5Q7t9650SNrM+/a2irx0+vL5ns9fOeXdhs/JZ7dw4
rWRrowNNWlu3yIHTsX0ohWDm3SbdP5k6aV2txkZNPMbaV/+3poyjJDrfiKWojne5
2cxTdNLR27RqUtfz0T8sSwbOuMFN74M9ICEqu92nMFq2l0FCKnz2xUdheGz5QIki
dsAvDFq9hOsgTZuBap1dsJcOwqf7e9BdylDYf1LiuXbo0o7Caa9FblT4Vt8P9Xcm
sfDYYFr93Y4SXNIRAmLUovndI/rq2JAOoSdvzOs+QFakR+BPmjwWov12U79N5zll
h4wRki73JFX9kjPAUzoqMR/k2/92EibRYeC3zhK18LSseYuJ+Cplh89GHpLIYu2S
URcKvYPHezkYMqCv2xG4LOsPsEpRWvqZs9QBtr9E+LUaF0/CMF1IEVOus6TdPfzr
xX9tv435csHrun+pw/5ni7Dg11azxhGrWVzGn9UjyYLYJ30j+ES41pXM5PcGQWc5
mR4nwThdAryvRxyD/6iVc5lMebkjLazeefxdAbLHHD0kZgdFWN3eAhbmZizIl2w3
9tcwZGzjhEAWA0F45xKxyAMEchfSiuCD2d/A6M9x1/tkqZv+vxtfP9XsZH+bHp46
RItzJfN0SCiKKFFoiymBV46nYpXGC1nbc0jgYlS/Cy0XrW8MR0Ige5TgMrqrD83s
+oTOPCYCikxHk53hTRQpP9feKuf7tP+GZ2BEoiUofKQofNCF91BwyIdP7do2fFC9
+9U3Qr1Qu+ANFfYKkLbYZTz/GrjwEmeVPdGhgUUcn9DTtuQkvza4X6WBnrSOOecU
ynCUSFW4hyccKBCw6+NZIR7OK5Dxpmos60UJEVVeduoVfMQIHQJB5Vx+r64Cn3LL
N5CjVLj5mKV8XJU99wlYj56Qwv7g2wqTG7oO/ySV/SZm7JXIB24yi6LBvaCJSKiq
rrhPxQnTK1mXGAt90YJR4ZNB3pf3l/2LrhXxrj98S3nAz+bwboSZ1++mjIoOAF+m
9V8tIYnlcV+ywwTmLmq6lcnEbVtP05nRECMAgX/435g5Mg16+8SwlUjirHfYWJhW
R5PA4222SPLaelcLvGjEcEYUKcGfxBozSGgkTm0CA5vh6Oj0rea/uZcQdLavmcqR
lb0ve0EsKxhIhUXMnjTbWMNS/uUpKPzcEwyFiNTcuknmFHfNULXsGYlmpGThJJLe
uBQkNRY7HD+RrJSIbaclU61YA9DNWvkSEkpW8kbMOhbS3qJihJZL3Md1Y50bo9KV
iaZCfjZU8dpfdafzzV3gU0WcnxcbensV8d+EVNQ8l9DAeqAcfKxwVMvLRkk5k8EY
nDTKepFhrZ8u/nmKkVtMvppJ0BtaCb9KDvtdf4Ze0vOOZSO7vPo4S6RlZ602XBHs
KLjCeW1tvIAgCvORVayXffcaoxYzfz7UBGnysEbeyIKv0x9zjTYha5rGzQE19NBd
GO/+hUHQo0rVjVkS+Vg3h7cEk07GTb3rcGbCV57ZTmlou0GYh2srojz7YXX58uQN
UIFcyHCL2nIlfsVncnGHOHhq/xPRieGw14avOxZ3tiXsgtQ9ixv69uO/BHZ+k0JE
tFob9nplfLNEd1VgEQKfO1y/6mN4xxwkrtHkYvbg2L4YlwrPEnOFAuYVNudj2Ps+
dtkK/RHFp/XX0DpABLgCWMIBYAYVWeqBuy57iO1MW3+l+ng4zr2U8o/YiYbFOjNO
EtTNFS3vuBjurHoIDx0Jgm6ClCA+doM2WJu/Oc2LgE0U6UKuVi64NKUq0OJh7Wz8
kDV52E8MFx5qfvgyvhOu84c5zfsVco19ZMOTcWELqL573cWRYpO9lPiijyh+cSSd
usTtSiuoeQTSFZrdzVXWUeRLXNcZZb6LhUaKviGOvXXVE+9ViTEzyNjH9o7RwpNN
RMksimY4dTjRcwdBhjGfjFrWz90EtSEwS7i1ZJSl9EqFI3bd+MjY8qMrlQ8WVq8p
W1X8aOXiwmf4i+/HTgsasQ13WN8Csyfd3lzCbemmedW8VtcfBoIJLdJfN6xUDSiF
gNGOLsO65UmwCPQQr6Cuo+RSkphvmNJM4xr1NEmsHLMt5bzvjGot//LvLCoC5Uly
6/M6hJT05aNeLhmHFkBWulfzdQalda+xeuLmPOWMb3yNeRdUbp3G7ba95EQ26WbY
7N9taYaWeA3ZVSmZC9nUg8bFPPXvBsHYmlUZafUDWifl1BRmGN3iO/LmbFblR2Wg
9Lk3d/oUr1X4OusmnX0LcPNHztL985HDVWoSK401XI2lX+OCxnpvUo7Gou26PaYg
8C5VVJDlgAdumOBuOBj4v1VBZbWSUakJIkS5t3LwKpoOLk+dEwgkJGKwnb/ukA0V
ZdwHc3AxeF1Jk2da3kujTpCouX7+uJitiBq2xoEk/MqeTCeIzQdbFFGwQkpRAUGa
vEt7pbs65IdI+K4fyKbX7Bl4w+6Mv+Gnw5M5aq9dQAWzoVWlMwI7Swwdh14C9Ms7
A3fcIvRMWKKXX4j5tY8dACns7ueEW2CvmqKx/S56tWflcKmYQk75en8d5nUor/RT
75N9BAHvoyjw79bH9S6aURgDxgQbd0AiQVN6zkJWj1s/FOvCE9mD3qWxdCD7jb0Y
z4qPDttiSxOEeYUee5+Tml1pVNhjgcg0aRH7YKJjmLye2mrPpOqfqnhbtnMBnZRj
4Pwh3unAJcFQtcDvQ8BbiZ7pvw4juGik/gfNu9D393/exOPZug+vgw6xJIv5xep4
EIjDIAoiysGPoQiHuJEImYkNDhkXJVjnQ0M5y4Wsq+DMLEX61oSigGwqAvg9VyGb
Z0U9rTHpu+u3kqTiil3Hb1Zpgpi6PR9p6w/2uY3oaJE/n22m/+Bl90iMmZfK9S54
39pw6hyz5ZywrPtxXV8AXD1zz9wNUDTXA3KKg7XOjygEAEnOzoJf9hl8mtrP/XgU
gwCQPvhFDejQ0J5JOeipOzf+3sbKJLUUNgnjZ3HPOcygLsBIOXgKuXfLgwbTjZjY
i/qwBpGYzexInnIxI7LhbRgSSlLLqw1+nM20TZtJwlHbGE/Uc5WzPTSuxbzGlcVE
et6dOfr9akmxL5nK9NyZ2qmoRNcnTyq2xfe2ycbsn/wyvKgG33uOTCfq2o75ruWI
u7SXMaBmEoyzbDJ8aFeQv9nrE9LimPKt6d/4p/vT8JeEF8qyT3R9OkVPu8I5lkNj
LU4DUJWtrrmUEWr/KYe8QramZkpC/kmPL+48xZIewFzYTwM46VjzgH2gSlmFTmmG
cD8WlBO1MAwyRkTkmFKjcPGD/v8E1L0Ago8ZYjfDZrMXv5ipbDt/PgS5EeWqd6M9
SOgpe0sJwUVoWHxrRjL9kXdC/rGkMCDfU8Da5w4PqcomEStv7YaGbotN8UXxyd2L
wE5FEUbOrlu18T5SBLnOwFJEoP1YW9wXLco00U6+wXCFMHKkvyTUMsAmVRhxR5LC
cgBhQ9vLGoADjEQco7bpx4z3N7EaGvxM08AE7Oulx41ZesR7Zxz8WAbK3rEJP6iV
rafzi0J3PCn5LFYvH5JlDmHHcHECZJBmuwtQKAlsAtY6/Yk70t5AmK68dHB+bqv4
kZNMe3lejhf3TeJeX1EfUWO6Nn7koleMY8XhAaClVmZFUfHaLpP+187kVcCjlieD
xMEuCUtgZvR8fM6N3x77oX/urlqpd+AuKcFGZ8jvI99zx/LAwbl24xWXqdQ12dz8
uuoHrxp9yIQZbcQzXZcGCFDn0XFyr5W1bXPVkTG+s0TBHZYGMQOHmBEuF+yep+cW
BrVtJKU+8hltlOZvOfsOU55HJVtaSzOR3WwvLegkRk2r3S3rervlTkCPJnuRc8Y5
bcPo1K0hDk1B2YLM8jFQfT0pROJ4wxDus2TY23S65tTjH/hl29KdrUeeU/lNkw62
p/oqC/KeRyEDfwODp1IkIuqmRBvz9VTMUVo665AqXpNV1ii8OMbSGzwGmr5sFEWd
DA1ew6iO7WmRFootipTLcMtzroV3q7CRjBkWcIimHCEkm6IbBTgialLhbks2+Aw2
Z/eNm5NRsJNkBHsx7tk154gWt8b9yQXmFkZt+a04fwDWQXwRVekUd9ZNOihtENc0
I/WotYs3TmTTud0Umb9axGO0QDkIvTe9Xmr2Ck7SzZf86w6smFBycAfy2w51uqjK
ECt/JeQI7VVMhskI099AOa//ui7StceBCttV+6kPh4EELTbPbrHHrvNFcvwVwvIz
L4mJh9Ik/Ly6XWCUeAcMyoaxeuiUzMeFvL2Xx2r4q1QLh1jA7JjnEqp3iCcBBqFH
Sns6uCzpIZCj24AMkuv9nneBiIhvBoIE9Nwd057G+GMfqjRUciQK5qg+YweGWxA3
S4HyZmaQ53OSY4m9yyvR6p+08r02Yuj2yOJVzwnjLmjmIT3+hCZSW1MhXHFl1pIM
d0/tDgqfmk9xMZSElWnHoMvPyb/7mf/+Df5yaG9AC38tiLRdp23fnnn9ggrTArud
CiGFkIvz+l2fXs3dCNHDmAmoSe8Ipw4Hqn+VjWujEBQGOUQazFqrL1r7DvG4OztK
PrkPCpJB9lsXdAg7+ES3uH52uiGel8CqfZg1f6y+m+xIWZjDHB6XYmQscyuBhX9Y
/8FLWgb6py2stipZNsnNUiSAnMdnmbNPCdnEli0gVLPWUO/GsdCaXBh8EbMzVAvz
s/jOTfaf7se0CUiyo72ZZfKC8M/kogt46OXR9x9I9iBmerM59LzyHAMeGfYQtw4W
rE+51lKSD1/JXdeAO3liVwT7hFYg5W3PFqTSFZ5639n63ZkgiDp1Y/fn9phZNklz
vXLvuIY501tr/Q+urOZ91LASsdtKF5jHrICb60r8aDHJpgcFSMRf9tERpkXPQ0u1
13nS83MwAiKQLfP+Hqz2bsbq2/dzCEIoXLrke627NeKk+rACqXtlK9hnexp/EOYD
WyvCYRs6jo9GwpU+uRcWI/UtLMbBDzNZVo9vy3thAybgTXjwWB1NRrSh2TumkXo0
6FmrCr+UqjsE99PF6OiwvT4aeZ+h1jpTNSpg4Ki1Hu5cjCmNjdPHq3+fHRxRZdfW
7Pmf1FU4jUT7e83ob4dkQ7ck5hyW5f9w6P9GyQVfeMwrYvpQ5hTKxHfW63pAvvG8
bIiAcaIM67e3wLNJWxefnQ3XL+X3Utc0v1XzZNWTI2IIGJKKbPlzBp5zpbAoBiQB
HJ9j/wL7evhJkPuGsSa/xMKWR0ZCfHmx3C2ogbHNti2s/ph+BCOEg8IEqVg3ZQre
2WufeUa9TOFFH9xBu+rIUHPj27+/9B7mk+T6cbLVW2muOFuke1NxwHYZDSoME7Pv
Nm64UMaoaq2OtN+OkB2r8Rq2ANxAH5SUIDQtYXH35QrDWq8qtlgNucs2yWf4H3IU
8uXUpMLdGxKRugU9xFAHfyTsmscmMH+qBGoiNRDip77rXxuHxQ5U25Zb+7vq6rrj
/qYA+RvLk4M+QTkCUhvet1jCrbKosH/L8kQZUPgOXJQx1lroSigRbO2qsnsJqk6k
13qLzuww1lk47pGVRx6YNVPAtpo/0XBwv2rf3pLvwgQjBLmpgrWF8Aonrc8ekznY
MB/e4rpa+1f54hrWf5WWaTuhQvaOFo+Z60WoAtD2YAus2BEcp6Qj+g+k1F4belh4
7Y+WuliBshQ1gyNkGSGNss3D8k/GzjW7Do/9909J1v2z6XhRUcvnomG8iuhPR9Pd
p5KKa9lmOCG9S2RIlMsOX10dHLfRbW0aDT8q6o1z65E8n4EBoGFC6dVpugeKBpX1
jt6HYvE3BNh+hKt5+fYK1sf7A9B6IDDyKcTnkYHn1X9gCEQxoEKMEB8o9xjzZ0+c
iP6zMZQglQlzl6LoMv1mbJ30e4QSx4kCF45tnNAB4PePmlEkd03mxcNSyhoxEEu+
zpfvwf2U9d19svpEEfzFpiaRRl1pQe75oBMdm5gpd6e3ukrP9uP5WcWUy/Mkgdbk
704VUmkXnGwAzjUILwHG4amhTddTgQIXWRKoEdyhXkGFsgf23NzTYklO9NvAKEoZ
DYQ4C0zG0yJvB6Os8XYSBu/A9gQ9bfCkM6EaoPl8RGVKn1b537G6MmGbiuSVgMgV
40bx7l9GCZ0krWLLRmbpq1lRgojghUgoRdk2LuDisSStsX2dnYNMqgVSpch0FTOV
UXbn8Xh2gRZB3FBPJOWhhlBqofyprHLIjdFlEgV5SJOisvo0LwZ/vIkTdluBXpmW
QVRwqzQZ6ktzNrFOdUR2Y1Tp0hZ7PoWcJUY8tSbXv+F4rHsJ8H65TsqB0JSJeLW7
0hkJFxzZMZeNuZ702Mi3ilOMjLlLIHwJigZnMDqhV4Fz3DUSj8msCgjOys4hqZrP
b9FZxCm8G/bNm6LH5AEPpjm4+td12s/Npz7vqR3ZYOGhZ7EG7z4jw+78/IATna76
+aYeunUTkwY3nm/R2kg2jMhgzrfcQ4jZ1mcYeKXFMFJu4KRQ2+qgdn9BB0hQdzU6
6D/yZ8y0s9TrEo5X18103xklW/AlhPi5VwkNvtcctHXk0fLM/gKGiDsJKkAR5F+K
dyy/jT/wCAIHGNg6OhvfsDPuN0xi2CF3w7wevVVok9gspa71KMGSCJHmEFLzeEZ+
j8JXXGBbD5BClRwsz1tKaH8FkBygoDkz3fDuLA72CkvAtcXcjkbcj/1eY4/9LTMQ
LQV96cdBNMjzmaJXJ3Zts2Q+ixNUbKeqFSxVeHGWg0rG/urr2w8BuDWFyCpIhM5X
OMwC6EmRagMuFhEAUbrhRKv1ScXNYOm1XaWmHCuTaIxN1VgnoFN4uuUQ+o25OCDP
vcoDw9dCg4fGtxbXMRwwOe1/aRRRhdP4VU1F89UUowhcKXE0UpKIcEZ08lMH8xG6
qy3mlaBkHqgdsaK031YYbXeXQLgnalYgt6UfHc+q9CQ//yqdzg+X0YyTo/JlbEMA
B6G7fGrSf4sE/c0CaKWwkWeZYm5N0TGwPcqgD3tqSnrOr0eYiqB1O1EneypZImO/
4pjT5MrPLzSKxRn4Jqcxk75qFUZojP6sXRuiHA7EuabJRHFWqt4YNW5ZydEhW7wU
33Ge3VpVE3cGzgTKT9L9xyFK8zOAtw5xMKp5fEroqjmH1aAyu+j8CZJIQskktd8p
5T/2eNnVNP9smhHThAo8VU+g2qaszz+6guUXa1pfeUkVFc65ZNJLrfu1Q3eK9131
CD+rYuz5YOl7HqDo1oLCrRMJ6QxKKPYpBufMnMo35atAXI32cFCQ+aDY9AzlzmGs
qQybPD5Uu2sL5XomSebrZd+2L/8PXbVVtoYjSHy3tyAa2wUroNkZNRgQPr1R9H4f
QOU1q1wVmBvwYukEIfEAT14GXSvcMoWty0f0BfIKTMTqhM6F2fNrAPMtrkvH1539
m4gv5w+TiUD+JiJfXJwTYPVDrccaIe2PYLsKUsUTJc/NNPusO02JiaEQGwNBIU0F
ruNHZt520ZF3dq6egJfSyJx8Mxje5ZjeqiaPWOvG8g3nwnmFvGrsxHT7KlWd+rVR
siPHSzT4CHOEaQ/rCy7pUKG/qb6jMRVLwEAgJv9ktttt4pgYRPRAN60XfFCe6QPs
XsOGG/SSS/rS2mWTaWUucsvMzXKzyaxIy4vSe0H6q29p0YTb81m0LHMSYrA5v4WG
ToSfRmxDTjmdq+1SGT1dZykaXzBksxm8nfl9nsW7ekRGLSYrspCQ6nBT4is+r/uQ
MKylx8E77fJe3sAt7CQfey91em6jW4YiLeUhWdhQC1bSJofS9Hwm79HkyUaCofaG
x89UhefN+lbb7OzHQ4gvmSuyGiLJddyvarHfInXyiNdsItPjRcFVJE1ljbDQfbrW
K06uuHeHYOgeXszAhhiw3VgyAr2jx/d93ZrmBSe8zp1/mXd1eoplR9o4Sw6+szcZ
X5PY7geN8VmgzeGwASGYGmb2/qH9Ygkrx97Vy5e9MPlyI0cmNXzrCs5U0HGhXj0W
0UVuKp8WyIqNWZ6upmWgqM42dd1o9dCkGwpCnP+gH3ctstE+Qr6Q8ZRejR0sQL9Y
ArO8k93JMkGLsH1Rgoc6XMRrQ3EGFKyMF2dvKYr9MBvohb3d5SdFNJiwLyHSTaar
/bqPEzL4wcI+i5nZEtsDqB9szAyqgPdq5p6vRd7U6xJ5uqBmpVDzWWI778QaWiN9
UdB1KNyn6ciSuM2+KsahoYD2k1EoZnGN/z4YtIBKMG/1YQ97IuCTgF5P9Ixd3IFk
/ez8LrjN9c7VXs9Dd3D/ToTyhY0QNS3wOmSZ/pvPF3Vzl3dGD4JYm5/DlcWwWtXM
b3Aly9fu3jYVypBdmmrKxXyo0av8of3vSCdJpSL+XYuyrmG7Uke8uS+zQ6PfxcNk
OwQTA+flaGLgn+Y+ag53gTKyTDq2oiWQaOwWtgRgNhrxY0dcwBHec356+5TOxz/b
eoOhBd44nRexpjnNKF9s4KvhKzNSi51cZgkLo3mTV8rfs7UQPBeB7W1YfK3aOSPz
SAR9HEJc+XPhxcM1ZQBzlHOZ7At9RZaX2/K8SgvGkTfNLHy7C5/dAtPMCQNMWNzA
/fph0/X20eR0ENDPGn6HVVuDry1kTw+ktQ8Gzim7q59BNjIpDOkXDWGj/Jm6WTyp
vTlOotJEXHC9WaTHxJRVmAoPG4KLfSCnjmeN+C6NvfIzLfNcER8n11iF2P8/WbIz
bgCystY1YiNNMKI2ciVlo4fHn3twTyinqSV8T4R+KtEy1lgis8MrP/fkeB2mHt+s
jRKzrqshP3QMDsmvi8FbNs3ZXRJywTHqvva359dQANnqmBQqC15z7JhjO9Pp5b0V
/uz1wbOemthiWibF3kowDvDHY6ZScym+dfWcFLu6Ut9OtXt+sNM81A/UzfhTxI6I
jNLDvJ+Hh5yiVTN7EDEKulGQXlOjpImMoXHp5+TMTgWLb9Qip7yrxr0aWQB8lTjK
OWCGq12+yot1YurJWcd7a/IzVDkt5rqkrQSxiB3vTq6MyrtYCrUEEM3rNPVSEaDa
g2wpR0B0MhJnFhJ9Jccptiif/K22BDaY84WWIL44svUP91zri9kpoDVRgnbXZZnQ
IL0O70xpGTK7hm4/mgJ/lVwSw5uskl75MOm314sM3wxP4OHdColhTX30v3A/qVcn
iXMVmwAxdzmP/GNU+M7yh/vc1lwo1onauGPvRT13ZTHQ1+731zY6yY7ZbpT/JhTZ
Ox+L4U6SlZnJ27R7nf0DVYk9AvP/+q+upfxfUQAkHUb4X1CAEUYyogDF8xnBb8Hc
PK7jfM2rXwELPVVlIxixoofdm1nxFyP5ktc/Yc8yqDH/woE2LZT0xCDEGAhwWj4C
MHr0Id4o/+dSOj2DcTZ5t7K4tsvNa6nqD3HlZWMiONBdinDKNFiNJRsSQgSJz4hw
dxei3jLRbGaJc8mWLYQZs42SWh8VohAGBc5ks1TSFvQwMFXq58e9sQQJ2+RUTqjB
EUW7dYwn4trdrHwRQzAuGPH0vrJ/vgkIMrDYi3TYcSNIFNgsbc8pV8yjRlqwJnOS
0TOksPxjigh0wc1b4MXOINgojJyB+r1bEmFoGifClz47xuBv+vFLtn3tR4gTLxpi
EH+IOFKDOxEPz+cl1JAB/4i1wH0lDexjbDcJfzEp/hO++dBTk/jWe5Lwr9KOUo4i
3tZ8OScdCRmS625Wz5kfyGisWyNEDMX6qBrlqim0zOyCJiZa/cCPripPTn039yzf
PGqJsgrh+eMohD1tdIq6O5J8haUUODxXWNi+jJv38E9SA8iQitz3etE2RLdQcD2E
3jTXTH34YODkUGG+mdKiedt36qH3oxKu2rdFAOfE0im3PfzKVCw+LwnQ4yeQI2lP
432BwfIUGvfU/xg1+J+HJuA05wu+rr7jYvZIQJTqSXt0z9LQDe/SRzL/MRu/ST/O
8Kgc0CuXoaY2/LS6SoB2ejLY9kOpwqg6Ds0/v5EoskHkcna3vJTtOxglrJX5h0kg
/trBgGn83S/ipDyvjgDcx06WmBEzUKXmW1O7puOQj038oeYzaHK1Yvc9MoJ5shLe
VY/BEHhYOmkmp1QZ+CZBhvyGl1ZRVCZY5nCBMfELAnmZ39Ert0JhkpupismBaLg5
jqAun0R5FOhE4uu/cFtQ4nq5vuiHoZ9IIcri3NliAdPbS/ygdAi0lwpRfDCQ1d8J
6lvH5qR+FZG2atfvXVKM7Eoyx36gOG+KU/boL2X9r8NL3kbTuFDXkmsByM51xZMU
mCJU/5FWxVLuWg34tspBjA5Y71GP56+bqBSC+wKmmqC4WxG+OPC4Rlxq9a2nc3mj
9ljlho28ZqqULnUgJFt1lVE2rpsqOuKUIm06LnnMJ+zhjXmotFql7Cx1WTyQna/p
onRi/NG2eA75uiSBNLDou7K1N4lROyDZGKmQ9sIX7X91KXHURB0wD/CZIyU3Pver
wbF1k1lAiAvVZPzNlQdit26w25m7p7ohLraKhZcQhFaKYKAHNl9XTcJWL2dqxWg1
cymn5wm5yU88GD/bsVYRS7mjs+TsNB028Jgj5V7vaE71E/4kDmFLJZQMLURigbkh
cX2T5FosFDmKdFtnHSvs+Iw/JonOv5kbJjwhd5mZeGgCkjsQ++h32qlNpao7Rcpo
igbiy0HNOSP8W9gGZcrAsQ3B17KK4rYSQ3pZCcoSH1FKqKaZ7dd/sMEwkjIG7Asv
u7yJGcdufO+5vmQAU4HaL2gGmFKNMlMZBSUdZ7Cmw/xDRAN/wBEZIojxJzPvk/9N
KLyLJ/ri1mJgfwtjaAugPlQMlNlpemZ0+/93eCWrYr8E+61LElwFVN6sXTxlJ5ld
Amozm0x7M5AHUGs0aQ8SspnQZhIl03x5cMXubNZAaPnvVwqKU/F9yRPprHfKgYph
lGU5hbMeoZhDkDv+/BPtWpQI53ycxK912KRZ8jPLnYRyN4ip+T1SePjAIsDInTBJ
9Q55ehFgOG4wL8nyxr+RgqHfzBXRofGbXukckq4iVw6ocmBIS7tvAv1nIm/8dND0
COB08gLfAZrNum55D4uo2VX5KkYWhO8rQLZzXPCx8nYXvClQd0hU834Gw5lS8rMI
pNtOoWighPYh7TozFgS8ZLmB4Dpe9frQ0XUUJFaqnmKTnNAtQligc8kepG0g5wz8
5ZPqDWKsNl++mO7gwI4o+0JNzLgQlSHM0YGGKUBBhlhuZK12ROk+SYp9yOLw/8KQ
WOOgdKPu+q/EcYWbsh+SFDtZsTSsY4ELWDTc1R1rpa5GL56ltH2BP7EF/+TxexoJ
R99Eq7zSJ+saTpiEbvGmUZM8FVlG3JW/Gs/dsRItOic1+cWPCeCeGXijTlGKldU4
a2/TPASq3rKas+bwY1XpCIwBMojvj8VUNvPYDmx+5fMFEwbiUHtg9mRY8/8+qutl
B1TXRrH6lwwYg5jRI1OAkKggrEPW0/daGF3ubWWR/2DIr8JHnD39mwCzNDpDCGa0
JrL6l5HXfYi6u8YCE740oE2W9AU8FGx1hcDDuPEFQSuZdzj5nuw01E9Rwu2Q2Eqx
XHpC7DHr4Y3K+APU237YxN8/Xan1Y6gqhsyPEgtbzbhtKUtsycHkSA4Cinqz+qar
rLDH7IlcLhejAvtdNJKgL4Z/3zK9n/DswqRsOkCvi2WXzANCNUix3WpYGsXeZuQz
E0nSqYck1J+FCcjVJ8OQtJJxxGGup0Q8dy55kArAWrP9rnTNNAMr1jaDeEsSaR88
Yx15SIIu1PQpMgfGc296VCsUGyy9hnY8CB7RUY/BEQFrPBYv6Xcx3TnJy+SrIy+x
9K4AIWguiluWd1SKhhGEA214oVBXuwQzoZn1NQk9/HqdRBqR5bVjpdJi7ScQts8p
veia3kbndMUWibeD0NFAWkuO9RABdV4cbMmAsnj1sDGUQUbxibTwJck7QF10ayn9
Gk2WdHS88QesxlYu+45eEJGr36gg6AI+VCFCh7GkIxtaryPtFhUdJoxw4IK/lGRG
7tEbTvj6b8xk81BiJ7Ej1XAxbMwU5VGIPxpbBfuw8faJdmgORMNeP3k1XnnVRLl0
ioWBKWx0UZgf6PPUmRfXCYBTK0eA80R8EXc5+APWWYzI9hsjwL7oI2B2ug6YGzTZ
LC9kIGsrFzs1f9QAlc0ednngUyi9Z/iHVgwHTlnhvoaRnV2+9s/ulkihl6Ant0k3
CaHZ0kiygHiIhsCK5i4cEN4Npaz1QWNrfNUKwJawJ9H5cScNqRjEi1cp8NsZfIjo
KeI5dlqzgqkOHVequ7i237UM5VlIGcKmzbMiWfwgdVdnV/2jI8gkc6/FC8HvJbWO
crP3Bkk+jqze9YA/yKb9xEoCLgrZ3u98ggP0vVhm4ujm5iR675ephrWF/X/pw67B
MVEDcfD7A/gUqUqxR+KVN+TRe1g/v8ZYsm0UxYaq39FYmGzwshgj4thBLOivgDWN
RgiRbyiCEalL7cnMZmv2q5XiaYMOxm5veXQR0cqW9nnaeHISb14Ud3wwIsuQ4syd
APYrhPnq+SuWZWsGm6Xy961Omhn62SEYFkStayxNWkAa+gIN+PCoZau/dOAV9peT
aPqej19f9hdDsLuQXJsx60+mQqPsnPSgabrJ/HPgeqGbfrVo/szkktxGAS5sMPem
63NGbbl5q3zWnpUd1plYRdB9GkCrhm6SRJg/XbJo7c5/1aB4tMuI59fxJI7VNFTt
D2cthkCHVqB1Xjq8hwg7MQ7XyYHstVUWLkg1fHWAH5UJyPMkF7sJZ6JWeHOuf7zz
sC3Ny1OjLrTuhHj52otqVkJ2SZ74s5e6AjOqbFoyLJmD3AE+rIo3ZbCb+YJdPR8+
GHkJCAc9WFM+GfTmt754vNg3Ha7h790wcPTc4lyWSYIhDlDvsTQNemBqnZO6w0e5
FnHrw53sSTZBaHmfJzCwUJ/rJNgupgCiubNEmNcRi5Fq+NaQLohfWfxgDRBSwmHI
L1f2hDysHN0jEV8RZCOjgpUSFku1l26Dtc57u7tVF4GMxtvTxJC/y46Oivp6sLx8
UG1r4zACcXnv32gywFtiWvun0TPrTEkZlvcjELWzIQ3fKYhA5iGtzWXcEaxUdYLl
GyOJQCbsg5EoVwhlAxLz3LrsSmiZdOXtPk5GP+w8hD7NxeXGs8y21nrt2y2skvVQ
GiGfxu0NkynnrUoxG2ReG0mkZ7shtwNTbiEil+8WLr2CypBsKwyLGoivGHb9mHga
SOtpgDjUffZKPMIwK91uUQQ1rtSdXTV0hZfv+xtvOS0m8SBvyq4Z48FHwONd7K1X
IEfgM3Rk8I6KTmG2WpRKy3nBpx6y1bT4Ic5UV11+8q/J2yJm4UPbaugFXRs/1DwO
89x1NBtGLppaFiya6oOXpwjlRtuel/VXv9j6YhXVT+4YMV+AJ50GRqhkaHsyBZ1p
PZB72LL8TmsyZGUugOlv4VcPkq5R9eA5t+UE/sN/wSzBrXcap64TunbU/ZtOsPL1
ORxZmnpPZ2kqsGvC6EQJfFXEDyNR1R03VfnNZ/JmccV/81CZU50UQyaOlFmlVsd+
Buee3m8CrbVTjY6GwhB9SSiuXRlvEofPZAOhpZFV6qHgdzX5HvPHtkUouMPD/UqW
f1yi09sbc9tCg31g9LD86uNOhmyV4wyy1BlxBDIKLSoI6Jz4TSAtfaStzd5vDQ/s
3pGAZzlTDks2TsTJH1LTKYzbyItyjaL+8daUlmeh3nI9KUvP1fhv5mf7gkyVQ2RP
97M1hZrXr5FJqUKmfQXepOm+mezQupD9bfwOlUIlVMTS0maVMrqsh0lIONBpVvRe
g4ySC+r1rVk+5G/CMOEdyi7Uhc4s9rLhAHT3Hi3h0lGrGd3nBbp9WFSD3+Elre2F
aFPvz07P1qbANA4hl/jcqL6akYfjAx9VOy4eVKK6BZ1WPOM/RGR1ElW/nrO5YXH2
2Zm3/hXYHeZMCBhTqrLCfHDtnZSA2T4q6TAqB1uo4LJSGCpGjtk14U24nIx4xGxc
+bDnTIn2SPOiNL/5Fao8vZuJrr31dyEGOikw3Nf6hnjClvD5xv/+1hfET4+o8wU1
RNLvpZLemayRC0AhfNM3HmSncHCB6shE1BoDZkeo4EYsofw8uM5NmDfliqM4U8tD
PWiOhR7bXW9oL4eZnf0e8cITCDFcCH832y+eveja1KHctv6ai5cdbQDcAKSfQk/h
c1g0p9WDe1hIIn7/XDbOmVCsuiBcMlHUgUU6q5Ivb9QgDx4Tk2Wci4w66eZqRAwz
3xMldMyPT2olEQ7p64NOioKrpgtK1SZwU84dW7kt/2qWmbrxcIJrvYbPsKAFZdGl
nWEWMRGcRYfNozlnzAL5UgVURStM7cSLXh2yfv3P4vvJB4banAJvfFwzpSrrmioV
9WOYIcCB0Xle2Z8kPNTy6ezwYZ6ykUjxFj8/fouOu8pjROBxSVzhP5jHgMjHXomc
ZUbZyiWPM+Cr/vZdRMlpUe0XcHv+4lrSkkXGLrN/GevS0wKrk/fWbdInoAAYjtvz
x/fDfvIwwLS7nswYVQpqe2lqNj9QUPCMIckR+i9T6DjInsLgpca+FBLFeqtftHYO
q4geVRAES6oRfoOBMbNpC9t/+l4jNtlxJDGGZN7xQJ74ILGMe4q19U5R+diUs05W
HySzEXFXdP9wV28aK3SUZMtWqOM4Bp4gtBizd2aoK017JxVvw1pOpvUUC8QUSy5R
jGI8yyaKBkPmhh5lnqcVlHo0LfLFcTJIznjFe8C4fnCz9YPxWGhTb95JHHNFQ1Fx
cBpqE7nXCUTvNBSWl/edl4cI4oFfKB+NRIW4fTw2HJ1aZdZwNIa2jjp993g2t9oG
ndFLPenrPHPDwHSRFmTp4P+4Cqms2WuWjrjwSdxtltncSy79kMverBJLR427T+Bv
o6fm9NpQ5q2fZJPuCNTT1g9ylpNR5Y+65SD98tPrXPT9d68sjT79eUh+bzCHVLd4
8cRHpwCwzoUYUuS6opD6M4tpPNVHhkLG6k9hpRRZDgT46sShTtwvgxMuqPFCma4I
UgjSqS+S1hMTgTGfZMPW/8axPZxuolblWStXBQAiUMXWYeLGm9HIDDaHtu3geeMX
MExuYPSXgUHl+XClqxTDc8qUGNVsC2z6pb2OVtPyVX/qEZch++6B8N5Ik2JNCV0z
lhuZm650Tu5LTEs1L+BVtpEg/pavcCEW4TP0KzL7P7f/d7c7LJgcrlyqM+Q2vkw6
QirJx8VajQzrYcLSBUaiUhaka5UXlYel1ctSOeOdknrMw78Qi2+cqjP0uouSPkp+
P6N1mcRVHMFJRCbwRz03ZlOdgBgzO9Sh3sLdmRgNXXSzsLzgbVwjM5DgzhR4eUwX
Wnn1w8IKtFtXUfB/sZN9zK+OPGtqN7zvcWTTRu3hSwspYX30aamWCUOuBfZPT0y2
maQyWpVT9F/x6Y2hUXyvH9MvGXevqFF0rM8aa+fruhtHcySwoGlvgX10wb0wdHLh
F2mqTqwqBt5foL8JXWJl4arzJP5Xxoecgy2AmRB9PBbpUgFJ/97+WS5uP9JtW8lC
RDzpV6gWLYn3QMo9x6W5TCY5oeKvcM6NNko8XzHQy+ROGgnttrgm41BodYl2/Ysf
CHlnDqwFIO2bHWLA9qO/XDxDzYnb6CQhYCqeGiUMuqQCti8vtLExzWCN4KZG5ZoE
6VISpPD2GxP1qGtRVajDplRW8sv+7CvHOWnYnXMesnkkwJNMRtZouwuSoJuhZ3os
IrE9k0TJHKW0kvtID7ztsyUv4FWv8/9UV3aT0T7AWHmvZpfANxXLf0TjY8FOiMaG
LL17j6OJ/kQU86PHISwQWZHsKkKZFozqHCdHJwpRpIFIxEDH/1KMbQnyBI/jL1rD
Mb1XH3c+hQeUGX1I4Oyk5Niv/EOXmzlH67kcBDu496c2y9kwooP8pPVU+C1WtVG8
qcf9r1IyvnAf42MDpqPBLmx3jhrPx9VJOiAXE4SuuW49untYZR3LACV5QJ4RFvSG
HvDOmnvbsoFgcdAkw8jRGKPdhvPzteZy3RQBngKDkGEWcBmqCDFOjLdmWhLUJCfh
nNtg8rXUcbh1JewKLhriRo4aERZZgyzis/6dPP4o6BxFrfQrmEwRCe8fznjatejd
x5WauHhHGXwamiGv3XZ7V5MVo+fTZ/XoTVzItDsvmb272Gxeulk1IIXbkmSC0K5Z
KD979+iJfZfyyzZ+5dWlyM5+4IEbgzAmGR9ut9dE65wpPaUSXoYO+PJdqCjtcMBw
NXN7W6GtW94ZVBdAdYvxakkkNKgMUZq5UuehtZ0jIG+bvFBBcRGVwCs1uYlzzknv
PDm+YZXXWzDZHyQM8zlxC6pdKwLQ5IuH4jpYk+gsGmnMNTs/UaKBQlWjGBu8cDul
Mtq+YH4tbHeF8GqbLS2Kt2Au6ua77e12NI+y1TLgANOdJF/h4Ike3U0RIzjhuw0D
SWSalhBADcHJymdat3/8YgFTiwD1nmFdqOYatSa+sx1SbZTnlKS0IEE53j8q+Ar1
dy9DFRdfGPgJURePGLFlfsz12tqyXjbQJgihR1IN+a1Rh83wUA0M1GVzl7cgeoQo
4LnhYJ+S1+C+L0MEtSTIewsrtfLwfYbDLI17k/S76BfWP/4rp7a1pwY5cIa+4CIw
0SDtVb7ZKGrqm8+kd6L0ZLkE/qLbolVbpFv+Tid893D+/nCfEwkL0T/VKHs7KWgr
EHxxvQIj/pDAkegQhd+k7dk8oujpX8yD0ESn2h4G59PYG3dAzbHwN1jcaGECm1wF
VSPtcTnF8NR7BX0gvcxCatvcUjCjn0uopDrrtMLrwt1XLH3LRwWxC79bmurCR/sB
frR9iwU2CCZrcSla8zbxfzxP6QXia9uzar9wT9v2yZAC4+V9FUc3q2dYo9z2ueJg
4SfR4dRiCNrBCV9Nan5tSeesIrE2FJLXmQPu+dkPjfUxMY9Idaf2KiHZmsr4SpVV
qEOLspItYGdicB7Vo5ifFM1oFresJ46eyP32ZJV5+IESptjhI93WHAx4BlXHLewH
Q5heJdErVhQevP2ilMbcHQvu2ipnc/A4Iy0lEfoiifLmDC77g4d0iRF5cyHVbCM5
O5oxTf5M9iDHE6leByDLuhQabuDuTVrF89xwA+vOT8H0/LxAp69FAiJRY9iYgBf1
wUg3ZoQiNpAJ30LF4eHFlNUfXv+dLpcr5LA2UCK0UP/FfAbQr3klhcSQGOh7iSDq
EPBe9LOCiYBTZeVXcuSIhcmjo2cUBMYU6DfsfEaL3yjqRX5nXTWbjVF00q/s2Htv
W5V6686ZzWuH1Jgtq+sJ0+hmFIOUPosDpsEK9MscWjFLHVELjNjJ8NGdcaeskzPO
epiwBF+y8I8igFY54+lMLR+pcg1wUsst7onV5EAUEFGe4VqJJanuiiEhPqSj6zvk
Bj6wKloNkzQjyQ9Jk+uBfqZ2TynP9UJlZW8pQJiPoztBh7zm8scMm1C9Brn1c1hB
Nc7SNE0h4Fx9fV440r2d6WmbHNSVhoandtyuTr3tZwIA2+ASFVBAubnDrPVwmRTa
sWYwIbA/xqtQ74CdIzfRjxzm6zFOcmBpf/oXbUZrHo2wW84xhy8OMnChb8D8BufV
zEI860HML7L51pLOsdNEZZ4bba9VpYKCKrR49xxDi4Oqevh5BKQ3ygxE2AhSEfSc
J0JUMVVS+3C30bwQPnmT59Sfq5vB1eb7qXb1pNFJW/jseh4SHhgjdwsOBBVY3BwC
G2jFKUfA2o/J2HALW83C+ooGSL7LmxVedW7NQUDEZVGB2ogP2NE1BWfogQF275LV
N4jlzp5iT5UsOT98RjNIGGZnNoKxSwyFu70nMSXdoan/Oxg4gFHlFxKzm30alB3w
jkR+DJ96a/iu2er2t1JKg8AReKVl8G/x4VLKEsMxnZLJckE7vQd05aT0kmTNTsuj
Caj66Tad1jzigS9KRY4U9hnJ1Legyd1+TYMmqcgD8xUXBztcRE2vs0pwyoJpqAC/
c1Qk26+2o3Dpu5IB2Z2ggtyz1ma4WEbOTUQelJkan1FOMUxAnvx6vnx04anbPV3T
pX+3l2yVXa9nRUCPS1UeZDtT9MzUTh+BsUQxRQRJ9igCHZ6nb2jr0mZCwvJ0QfBx
Wg/s9EHSmpsMXu2O2dlyidVBZep88PZME/k8jJVoTiKq3/5Es0rymeabJ+cKLhh8
+H4aca3CzYl77nOSzuMp4tMT23ZmtBeh7rs2yZsbQGS8t75MWrrLbiwmSkc8iFX4
Ms9gKyaYXN9ZfjFTtWEABep4fDLmconNJgbV3Gbq+Ut2P2an/mld+2CWohCrU3SZ
is8b8fF+XQtgSlzPFyYPvhgMQ/XaCzSMNshtlAigwGN2tQN5Hcpjtz3M9Nrnfe25
wOrqCFm1AL49CVLTErS2JcnyF8EgHWP6OPR5nYjV4JqyYx74VP2R2RbBZygxhrUA
1uYJ9GFLIvBcqbJYVhqYGZfBdG3YlzralEfSCDrOxndB8ALehXQ0/Cgkn8sEi0l8
KZHxrAq0rpFMNCUlGZRZqzVppM4l8o08qL3zJ7hqWkIRNAf8KJy1omAIQkQ/WPdY
qW9IVWltfGiDYK50ApjcpMtzE0b9GZX/ShM1dfrFMSHfmv5iPt0YKcLgP2OiKBYV
6szWa6ry9FLqh35oa5gMzOLGlaPW1hnz0sPGY3rO3olWJsyzhcVAWVzWylIT3Wx2
f2Ug2upsmpT1je2w/vkz7jmsx6l3fhcvCgn6wPjKdq5qm9dJBN4IKFgaduif3Qs+
qJaK+fMVbH6FvY4dXVagGLm1uBw8VhEfqVYMbkYyTZ/trvBsW0FAQjx7gDeKV9nT
MMuGEotMG36A61hVrHjs5vD7V7GUlayn25eqxV8VlQc1J+7TKB7kZ0C4iBsUhl6u
R6rWzRVPc5oBQ+o/gAtE/syAakYvPy+GmcPsMk8TDoHqESue5dCucJEAH+v+R9wz
nSU0Sv6RwXAPMO+3+MbbGEXfNEimCnONu72c5qvd6jR7V/mQj+uHeFidbtwPGXJn
+0cCPb5HBvtCI6vbNNHBDQrpvoFiA0uJpezTLZS9cz/dd/UM5QX0DvmQFeFrKnEy
fO0qN/su3bSuORCBmHvHULhdoqNloNjlh1st4q/womsI5bzayQJJmjUa0P9KNvAp
+abeUTvBZWj+JvZnaY34BFhNMsrN1KW32pCFScSftFuAnIv6tht82x8olfqVKPNy
AfaDT2GAN1eYfBCb9KfBgD0bsxKRm3ZpDnIJocEDQ1iXGm0GHFgNiWRqECvgUtM1
rYENxkOaQfn9mZBopRo3AZ3NHTabZJOclFC90jp9lp2Mi/p3Uy05NVtmBDE+t+Yh
zCIffc2q7gU+G985rpXO7XjgyK++UEKn5ePuqY0kQkOXHCSbp/nfzn+RlRIqcIOu
mibnWUBPeAF/j/AEqbmC0GtwwJGKeIDQTUrjiDZXWwx1pWO5PSgrANZW1NOh+4eB
tqgMctWVivV+S0UCWWncVeVDXokeODbcQlmMj4354pymViZh9vRO8a/jF/hXwYSw
hWDtBHHeHlj+NYkbpU6UY8RvCASuGMLeuJ6fTGv/sPQ6HSiH2myt6ZxyLSFgxdgz
48TeAVTcAvs3dJILoirL6hZcC/ruIRvGfyuDnHtaJ/h1u5AUXL6NrnNHkNdhu9yD
cF5by2tapSro1C1uKqmIy/UC0eunH0msp5daG0GoUBlCdIcILZCy9DDqRlGsK+no
4sh6AHl85a2WFukCbANgY0eSBK/7UH0YwrDHrCwAHibtYGC42o9rQc1SaAGrHXw4
zq6JrvbKwu0ouuaCkCFrpOOM+U9ppeR+d13nBTk4Q8wdVMStYQ/+X8kYEP5MsvYo
w8QYcRH0X7Qp16033lpOc8F0XOWrUqjw+xlNOYVEyrYurORrEB0YI5wSdbTue7BL
kWDfq01f43XJigf9RHdAvnmdjX3pSzcvDcckHGo+LGWX43zRr0qFfFhcHSVkmcTm
X9IuF/ahjyUJk8B1zfdpfRwb/KA3aodowPD4ht8QfGYnN3y4SsQUBJtFJhBCnOZ7
nX1TMiFWQ7tEJgS+HPx0qDfeQcWjFeA9rKfSvOcyAR9SaxOOT7/5OBOyGWNV33GS
JrZhswYpT250wfhSoa5Xi1K0hrpcKQfO1NZNu2J/rhR3pixRl46lQxX7vivczgkN
aDoEbxvgEFVE0xZLCiUzrzK3T2wWLwi1b9845NNRD8nhEXnQlaVMjN7xv+poRzPO
lKyAFdMnpMgh5BBoBzgyW4E9m4utB/u4tl30qdIQ6iIyQoqh9yMTUNJjAD2H3wyl
JIC3qlg9y+mKWYRWjQxQCdXrOkRTRVkR4XLKNzXWDvlUiRrUd8cs5iYwxbV8CPja
l5CPnfAwQ41xGdEv4bfM5GFu9lJBpo1NWE217UQ9HQS7m3yRgkD9hYYiG/O7e6Tk
42QY9IleeDKICYdS0nAnfh8ofrYS37DEt+dHdEEZTUtU87ackFMaOlMnRzdb6pOP
urfu+ZP65HvkuIDSVN1AzojI5LCIqdBdYHCQGRETGtFQKB2EogKEkvdI9vHRkIAb
NZwbGZEoNIuown/KfAfAch2ZRTQE+2XE29D4xvxsItX5S9eZcEIX8iJyTCXk8G7j
f1rWZhdiv8I0d2XECo53JNhKaXn1OvCtXIjjiwh6oQAdHboM4c7s0cJJng5+0YNu
2S5VNwzk9uDpL9yRFF56Y23LHncL0UI2d5P6xB3v42SaV0x2spOjaI8rpRr3Og1l
zf3vB0BrBkFRVXATY3scG51xX+A8ALiTOcDNrwwu7+o4vZLcmAw6j+jsJk870nDP
/U3ijB6HjVJ6ul8gMiuGnXuGV7yrjzc8R0Zq+6uZU683iZt9QL224b7PurvLthZb
pK1inBTNIiaLd+pX95Oz1p9m3AkTrZYE0aw7Zx1Az6kgmXM+mXnvq8E7QjHbqIqf
uaZuHcNgL/C/Aw39f74TqVpFFonq8PZKFaKna9m/XNHIUHSpxIfmHbR1MgfDM9wH
4U1v+YXVek/rJwdxXiBbedkPEkQGRgR1h1O4CzLb5yfnedf6CM5X4lXI9b5GR2aT
lxJ3b1KjkxTCWvlS8hYbPEk0sF52kthdJW4e0ljlHCPC9lHPtoRMQm0zS7f+xU9s
gGc5hNouVFMCpaELdRbmf1J+5hWkg+nAsRVBj8GmJw+BkbwdvArgY83JmFjQUH+v
CDbtu3hf/VSzrb1WP6hyK8gvw9V1c5KouMq/rrTS6fHEx8l0mBVx7wX2LUqEvgXG
4ZujqmvwBEQBbPX6ce6p4trhjN+YVb8HKc6jIn2XFjxLQ6JPZV9g13jYZNVpZce1
IN5LrmJ0a6eVWH8Z1dRhk0l7MLVbX0lqXmu6CPYqOh1kk40mCyRkITbBhAWnbqjK
0ZmC9QW1543zxhQDZN9yafAmRCyesMUgXrUQwE/xOS0QJMuP0OONN6HVw7cg6AwI
agYj/rSx90DeVazZPj4AILdjwz8RL/omTduso9u9BUS5VHKs+63g5z1TZZYF1tGf
3VYHxvtDNZUDCqpJkW//eJhHNvNOnqQYulddXZRSs3VpNg5yEjvHdh7zBAtngYB8
CmMIIuk9ixH5TEIXOHRcnCP74kxtyAnuUWH/7GiyvlOaLOviaNV2L678rfGiuZ3A
23kQaIQ1HU6Imia8vBfmxefBdN1ICMsDuuTRbhGiIK0y4pAJIxy4m1vMPB7LVsLL
8GqUEeESpcHb9TMwY4cDv8at1+viOdz1SXFUMu/qjMWeua7nXm2eTqAzjiOxhQyK
ozNSh/sCMlZK6S5TM23qktSInbJLyG4gq56ifHx8IxBWQ9HuxQzlrsOE/+qUjsC8
oFjxNZ2FcPP4TjmrEaxg7PHWPTjwJYwOgfEC+A88dNFWOkXCqXsTi96t+9uI83By
K4jo2JR1PtJYhy+s/sKMeI2zC5c9W4mDLIPTe6Wy2MB4CGwvNJmag+UbKA6W7a5Y
jOECXmqUThBd/2kdchf+i51whGpuoKkym0pjXA1Accvep89YtXZRhjcWk0oh5/hx
H2FA2b+Pv4DpOqB4x7jW2vdwZ9Wu01qhSWSjB0QHWYVR2pvP3KMLyI3kbGB0cbK9
AiQtjGJta6n3mKmn9TiJgwPNCXRMJP5iFeFGthG/97gGmpLDRpSIXowAoBT7igGG
2ghzm/f8sA0kue1UAu7D3Lwwxjk8DEnNeWqzlZhtRfw2uu6KgJ+g1AT8ROIRP41r
RXj4Al3emQcL5nhrqrGT/RAd6I4GqQTEA0xkyjHOTCtGtvfVbT+i1dRM2oKsnhDl
Di7XZdUFIEBnHSQyAebTVERr74kdL0777fet1QnuBIev/lzrFPcMHCAtY2GbYVDC
quY1z5iCNpCujwL/BLr0+Igf/JBLEDlUenaD/G2DeMtFt5ujBcYZ4aTQTBftpeBK
6sn9Pc7+pGfrPtMp5rEByidzqEjGT1ADwql4Z6lCKM7vSWItz1synpI7jGD2Tf4j
IBqd1uf6kh0hb7yGv1v4bLDcIv57yxJNioqG1+D9QmZ7tBFfQX6tF7KAY1iQI/xO
0tqXRU1jUmf8ehQ+Dhz1Ot3HH/6kAYDgPObatqixHV3iqLANnPHuEMdBEQj09zf5
RS6oliYUSi06cLpQ6dyqqovEYcZkSf2Luc+5nrVcvM8r6ip2IzEgximlICqSh7vz
/tiVGB78vqBy2F7NkCFAm/hrfn9SweitP3j1DeovOYMnHhVukCP8AovnVkffk5M4
6QkiJDVvG1P9+9FcigCVpnfhuA1giUmMpO3GjT07mzmpFpJSZw406RzySl7rDbwJ
bbXVLXgKnrkhwwwW6a+TFgo3Kc1mDt3HY9p2dWWfcKEuvlU/5MgCtQtwHrahw8jI
K6VyzHVQNenhtsSHWggResHuMhPo5S0z3haEXR2TiB6WhYc5k7ltT/UHc40rtLuv
xfs+gU4vz1bvA3ENm5wq82V/h61EkaChJa3PB4PAauO2RPFU3ErJpncbOyZSS/F9
ztvPAlxw64rnjbL6CSzMVOzXgjfMrFTapCtyubcTNtXr40SaJ4Qar2bzNmhjl01z
4GCZIjQkuzDUXyoTHocr4H6rAprG6VQJt6m9D+kz5Uxyqn9bvDsv1TcBkumz2Op+
dPP88n9rKuY79fHSzd1xwFrKD3QvxkDXA9b3AHIlcTzNMlQKFUY9zSNVx+65J4eV
xIyBGatFCPVjDpqtQHI4DQf5nOAzY9jyoMag4eboU6aWKtVdz1BkCNhLUdKMCa91
cDYylK4QE46uhuNXP11Xh2TIcmL4bxy0jkmHQoiMtpoZIgWHEHaxSTs45SwroAMw
6GBAowIBpDy2da67oN+QanwjLTAZPF2Obs7R/kAc2WhDGLdz9frjNLOKTKIsgOr/
ctfbCmOzyA8tzlxBOPBZTA6W2bYMQInFSioANot6gryGYqhwhyhDqAaSaIqBXt7y
3L4LWA+z5AJKijeeSJDhuippDa3XzoJ25PsikAEnOAtKkRQl71mPIPoCjXiBefnj
vvm6XhXEoq49qtb9zoYVgROVweMyOeZTGY42y4Fk6JCcDDVMril8vfBXVAa6KcpE
NYqtQiLQy6jzGNUHL8Ws4XHu9HabQXvXKJS67Km7jRwliNMdpnoIEnuqDzokk55U
dY9bNCipCFfu9Sug7AQqCCeVzYHATwgdYaqSO9pZeCmjlQa5P5PNe0IewQr6ql67
Kl0fys3FRZd92yvarIr8/WSEbGoDjwFKO9/y4fFDsT7hQHWttp+TZlFwrG2HOxs9
zzcxvG4xQ2Qzrapmmmi3heP+piHJScwrbax0Fac0f2cTDY272bKdm+Yp7H+zFD86
5VdKXm8V0FuYKJJqG0amJkaivoIDaF2eQPrggmeK2Yayls9j2HfUydLBcgWTTD9Q
gjsOcXg17NJotj6lhGz8rER4EFiyNJ+PiRgW55MKlyDZh/nHC0cH160n0xLvEvY/
0RFLKSJiaT5HittLLlSVwnGW16k+GLogkrMAnTkStww9hLdlBEyhNy3A8KuPqXrh
7RoiehTC0G1zNc6svMvBv/gvw/QL+9J+lRiGKEvMH568IA1ievWf5m/Cv3i5wvtJ
mAkd142efzFrUr2LWxBb7Dc6MB0sB8j6xjEu94aB+T4W4Pb/SVofRQ5fQoQ5ulia
lk6wN1EODokGie87wO5lQ+q8E8iEExlTj3S9ZiDcC263NldgXOWaTvEqDAP9R2sf
aYzBxQga+R8XHjfYlRt0iaUZ6VEmI5KjrRx9ITDhF//tb9gjF6wc4sie/xrUvBJl
1CDl+A9PtH8+1JjfRwayjOFsfQdQMJe6tfj0AomoZBVD/9rkHLYuc4Gfdc3pCqS+
Gr1vMsr7bTagZTnHuobRfhbGobJkyiUVBnw6Oo9e+y3Ih/kRWbvVRAT6bn6TramP
uXoYidMhGoa/k9e/sbFHyfSSsw/d2lz4NRUNiERRZz87Y8wc4qa9Vd2SUMWoxHYN
8rczJRf0Xrzq58lulMANTGn/i54hp/ryF0eIVJeN7TlEeEuzQHk90Oj5/bAs+yrS
2Mqf+L88OipCRd6/rGY6rIE7K8OFJsYi+folZVRF8IYl4tgfuVEUq09Cub8qTTQx
t5ILkI/KFvQy/RXOZo7OxNgCDuEA7LQ/9Q9Mz5tuFxZGvqma5t7cdX2zx3aOwv+i
OC8jKa0d8X0dTW0pP9zG/MoZqs/tgakfLRQ27EJo1pQbTtOoKlg47La+qGwr4p11
Rv3N7rYCkpkMf+l7sO9FI7MQB7WnQqNh5ihk91UGuF5d171WkBThR07F/R+X6hMf
dDerEwX/ClDMs/SnmwhSHU452RhIMYvEN6SW2Qh6Fo/ze0bRK9cOGCMkcj8W/j5D
vw2H78/WAaeCoYQpxA6meUlwJO1fQf/XFu/0ga6Lycnbs+J4jmmYPDspl236Ub+P
vWhKO53WNqgyWlSN9TAgT4mKosQ/TlOVGftfTGL7gwq7gPpEAlXhZgCcdXG6AznG
2lypljgUlgv6vQPm4/c4bJ26W2mQSMIg0UGVx1NzjJNbl6xvGB4D0o7b46Do4SWr
ZUYKIFsXE/T5SQWkKseAVBYliJ/CD8HyQbtdjeZ8ey0ykBvzR3XwC6JIWfGBCrKy
aYik2x25G18nEM4EJh2QReJ1GEx5rTqBr9Bv2gBndmpJdtUbPsyOeElNJcnYZbnt
BssNaWWeJ7/LqYoH+aefki3RKNYn++b3C5ZMmNfZBdA0w4i0WXF5Qi1jGA5bMF5M
efOu0ccD1J0m12Lyb/UTmCN8zRLQHa4guEC1xIfX8QEWMCMGJwqnn42C/kIWH5ZJ
l/UCSOcTHW02MeKAAi/zdwQhS3uRrEc+TssCwYsKqN6ML6n7mqRhZUnwCUl++CMm
v7ygct0ciA1y+RCVoCjTJ0iPYbRSYe3ddvPwfZo55CqJw6RRwEcUShE2B3KFFANL
Eu/Do91FjpNbJzpzXONtX0WI2vz1tyPromO9YPgENG1LuJwUeH1ccYVISc17YKfj
4RoMnWvlvSnLETo95vqcDpGSBAiCBrb9qBnjHdH+NQMr28gCUhPuHo9I1q8u58xG
Es5iEgVSxm2n0s9i2AeMy6Hs55MGlm0xLgvcULUIwT6L/0N+Kh9nr1jJNo9PwjAn
bDb9XXxmFiNsdtv1XM1tUfStnlajI/ETjVLHLS5FPh2oEgdfiP1BhDyMr9FeSxq/
w+JMiXPj5se33k1Fq1okFRKw9lKjTR7uDvVfhisa+vedOwhZwR9XjJyGxzsxRyEY
lsa41lcGgZ5R5YInE7uJU/NrGy94/LhcvDIFyJJ6YP7k99oieXeHXQMQoU9FZUdU
iU8ts3w78qWKqGaey88sq0KyYl7ATQ3ylwq2MZIeUv241eih9HyYQhIlvaZdJogE
Kz223S+0EVXqyvXNNeQTyPwpXMaETZvRhHhIisQIYgHcECWqj0Fpm7mxjlg+ze8T
3Xq20IcNNIxW8voqrdpqnRGSyaPhqrjTvPwMtzSZ+Bi0qY9T/qpLAaoOzF5Kz9Xr
vGv998zHfMwri0cL6kfIRb+KwwGMpXWosmv3S8eSOFPS2jp9qJAt3uVmOEbGD8UB
DbbFJ17gwWVYzRQ3W1R4vXcK4Y9u+R0324FkIEY9yNrHmkq0IsfIMV9R5J56c6pH
ERKo+VZNtvIQzphbatKOQk+twMSK/NrydsGYP2Rlqy13V/6A5S1FUgtGfoc8gDOq
B0izT6kYB9S45NeAhbDPk5n/QnbaEj+lZ+/bNocG2BIXxdKE/pl+12YSXhoyxUkS
RVY4wRirL0P6IUXI7A9/hCEW4MHIvz0inXd14VDniQ6ly5/VI1T4D8hwjAjfBstT
dnsPyIZbKqSlLD62mId6Vt6/AcqYyJJXmW/pZJO6UuK8o9VU0bd0fGFE20Rqp1ON
v65tBOpsfEopLyqkqS5rzaQwCId4YMpA5H2Rsl2hiR3tEYdw77c3F2r5GHb8e4BP
9Par4ZgkiR1g7bnsxikkEw2IAVSou21hJ/dJ5khG/YFatJEL8idY6R6gGUBAeY9I
5Be+8aLkUd6CMqijaFdpgNb4CO5FPx0YilwzSyjRiTkHKJ6XpyMp5a04XPi2QSZU
eVT5ArlS3GMZMxxtWgyCA+qo+25fdEXA7qvym9qDjQBF4+McIdHDCuqM0Ki6cWmT
clv00p8V6GfHZB0sgME7aEyw+JoEjL5Xjg4/tFAzkQRY+BECWtIZ+AEkKhsfwMIw
rcq3d3UhctULw4qRXc/MEgxv8FAVixJ3U3OZckbspuTm0XcVbL0cA4sXq4ZhxTry
A904V5W5Oq32A219YpTqiHYolNLMSRsrMJ9dn2bz1ZhUFGVDoyeVv0ndRaVYQvUj
4vlkj2wD2naSLJ3pWISOhSj4zQ1Urmi1vQ1lWrbdUzVR9IvHE52pVVoIXpaYwP1N
K3Z/OoWjPreBY5yPj+7+g4ZqAbHiXhPM4Znw4W0DVN0Hgct873eqQGdO5GB0mSSU
xZj4cZDjvm2wYTnacyKOKPAMQ7nMoRbDBKCOH3I7CvVZwY1CxkcuSjNT8G34LMDy
F0SZP465eGDs6N733yPen9JX8xAaR6BiMz0vKwEQE8A0BmOw23w7gcF669oDV5Bu
WDUFucYwGLQJWLnG3VhWMKB9VGzuVy15UucctbiT93jwPdDizulcgpTHzyu+GCVk
u5dDJGQXme4RDitRkfxzSmyfL8JQhgcEsfSrOTt249eW1guE7NcvS7SOlKzq0IR4
2RUmciSM3I1RpEtpV3fHOqWkTSWyDi8VLTWZXo6K3bunPKTrzoXILwIV/eA1+0rT
lal0RU/2V8J2oCTBfGTGJ8y+GHzcou6WgzqLm9eJHSfjAII2FOOdkLO431amXPm9
/Z/tlDZsfxCiw0sm7VEVk7r28cY+nMHyOnifSHwNJMLJimTQ+J+jdpr/ZPoOfB7V
DE4RSo5qldpkfbcSX+wNZiv1twFhv7A8ctBpcCiJRFTDnkZn5pd0TKLcKehdDBX6
vxVWrVv92Yb2HNa7Jrn0iMFRgCKMFFsXGRPuYPZrO3fSWvo0tirraZQ4E71a9pBd
LJCUHpiKvP3JIfmK6yE5redxmHgQr/843peZ8mwwPiYxb7jdwQNwKUHwYVnGCoCR
qyYUuamfGl1B9y3Htp8sEgJ8uuzpOIb65QqRQW1V9DwTiT9Mh1S+pape4JluaepM
khDSmzUlqBRE8DN6fbjZW+cYyaMpHLDgRVIvjmaoaPuVJJA2AnikhWxeh5rFnsz1
SStgruJiWDzVm4sHhh2FedKDePJjIPvVqBwyqJQLoQh4qWVplArMnK5JJenXRkYf
61VcXrjLGkkHmoZrzVKmzdDohThpQVTmgLEsJsd3hzV7Bs9yh/ZrJdXT5np3LWmX
pPLyixX0gNcuJLPMFovptbhmbThSsGnUAQHVPclHBtGMTmgV5hMyTUi6weigV95d
Yl6vVrEKc8v/LxCayrPmuwv6ZBby9REyv8pdUgvMHOcpnpEOKkUgqoU5U2fh0AqE
Mmfoj/espjRbfmeFGv/ElclCfAAwF6SD8MF6iAJr4fmWMmFFb5GvTYQ6freGXAwZ
iX68zYL66TKzxYUir+HNoRJkFyP5KzOHlu+fPxs0jvqNoBLRrhxtIdiy1tKHS2Uu
UfSK/D2CwRroAGWwLOlTYDw4oBXFOMxAScNKzjfNmyFZc2e1F28dfBWdaxWWyBzP
DEs4lIc1mc42Iie9ErQpHTYstOkzez7o61IA1nVWhNjFf2Q4DbTsZQqZb6RX5Mt7
Xzpr/e3FopgOFnBDx90I/y+O9RJik8UGSqoxW8ug4/w1YdE7PZazOnT3HslTpqzD
10VxBP1pB/8tw03VS8iMWKigoZEobWEg/iPVrBOaXEk7B7eTMOKi9V6uEcvRdGPn
uFkddW7hw3fTXSwBbNC3JSnZiFxSRlKjzwggI49dA+yinB2fE+EWd3qw/F4tizl2
nzKcGRh9sOjzMFKCZa+mMV3BfMC6o2nqlkK7jlzKC3XXY+JmM22wSVblUd0vPDMp
JlvVjNmurFEJCAB/EK/CojxPadcNvmoBzszzrzflYCtz4AKiazR/diWdGppl14ou
h5TQxVDfj0Ztk8jiaeMFj+/2+gt5edmXEBXmLJx53sayTfuvR+fbUzypMSPxeY9o
NEO2Q6EMJfRhZiAsPxBWsguC0wbWz4CVQL2hhtUWfrRsc6M3shrYk0eF9PtKIyHm
JmOcov4t4po3/k6+uoYIYSDLpV2g54iS9Whu3SC5VtaaaBNMb0yDGO9SXIkWYxHd
PFa7TgjS77whi1975GwcEptDA/Tj6AJaAzy7hax8gj22nSHG9fKveNwXljrgYITG
00OmeFW5rkb9HaWp8nTOXvfMklBtcUZkLmVTb66T8B19ppzNYUx0nwGU2N+7JGin
uahw1QO5F+boVbWVMV7DalRtpaK6HslDrf41WZF37ahLHQe+d2/Ub0f1iGl3ngZr
La8lXsICeyXDPudGyH/XpFUvyN6aI/xN1/5TxMJbqv7CZv9EHIgxXqLTOT1o7+KW
d/nPLxrLXofOfMKye7Q4rY0sHbGXMPK1lRc/80On6PeBP3/PmSD/CJCvieqftv6S
XBJrEkCoRT6h0rxh1YMH5Klr6aOkU65TNxOWiMYwiEqScCRYjyizWYQDnhK5iDbf
+aEJKlAq5ZUr9KhLgrBObI8IgJwX2PRA0i7mukE+bzVql8AP9iXGQleTfIAb0vX1
o5mzxHCkFNe+a8ResXew/fU9Zt8giYzHUhbuBlDbodt+fGs1603BSDfUrELXPkT6
0FG4P9yNOXY91jf5sKT2zWo6TggF5iUhKtz11pJaZpfYxcsNtBScl3P9FItyFh7k
u4zjD4kFaV5DWVuPEaOEMMIqzJ/SdUfRtpMV1fBfg7uyAwV3RdRKNb+TfrjiwJX7
FtVtJu+pB3EXNdSgxVLBMvdIcXAf1/qu62AHvGBbnf3pD0RRyve7FF1CyWmuxF3f
rSWr+G2Ido0y/2pZlL0KjikMGmWmaLMKd448hsYh8C4DZGnXk2lyYTaOsY0qQDw6
kR1zIDGiZ9qaIFFB9vaL2mZ35JSvyJCb4fiDO4ytQIl2L9I+4GJ8Wij1JmeL6qCm
77GvV095JG6eX+yzTBkbOClGQQqWOQx6Jy48Bpt7KiMoy8YDSKLwLygrNMA/Ar52
LcjPHavjsFG/abjvd+hiejgR3PM6OMP2wXnc1pavRVksSwwz2GbwdBvqspfqd8nJ
5Q/7o8Mc28NoPT1fvEFZwNTdvUf9Od3fGy29mp0WPtPGB5z4Aq7gq8iSdZyhyhzh
nP74+ZLsoEgzHxprHkYeO18ezeykQc1WH7XyJrADV/fLweN166P32r8ZBEy/YQ0P
bL1Br4XL4onIb8M54PHCc7EshsYOJs3HO1EqRg92tuP2nj1HrBZTdT2MtFdZoyMP
NakkTLc/E0mXIx/uCVtU63bb5foS58Y4dlMJZFEM/POj1u2wQ4wvXldtlbRPwWmx
bo1q/i9Q041Ju7cFbpDc82DK15OsSxgLLD7t7q5HhPOYU5kCgjrJdB3eRPhYye7b
+Y7mw1KvRe7OjHINjokl6ySk3z/1etXOIeALYt67Q4fl61O1IPmRc6aCLzZ4pEoo
T0URVCtv+oVLZbbjFgglHvY7whlPC8NeSVGQJrq4G+P0EGrJpJmmXtZqWisXDMde
yqHxE7Wj61E3dtXc8px2yDdAcH1tpF0uz2w9OBo8Xyrd6GkAouLsSvsYxuJjQ9/u
X1PRWHT9VhMEXk58K9SVHtiGP6JDahOOK2plk66c59tWh18RSfqvn+1vL0DZWxvz
9Sm0IFUipVwctJBHKfYEVE9a1B6kLasoesDPltXgthazgp6cOHEZ5bla1gMZg4oY
ICpExjGCSoPHktSlVLXECTJU6tFlLfQYXVwjeO1FQ3mK883DaTLXGvHo4C+B3VbX
duhK8zglReV57gEusRhEGfKiK5Nc7ikJzUKz+ke1c7l4q22vfbgSZVDlAUeRfHHz
mRsUKK+uwWw3J4m8+CBT0LMgA3x/P5CDmrygh5qnjkEv9igEuv+LtzCg+U+6blyu
7qpIajUwN9GkiFM4ju5kI78CO7X9RLQ1OpJmCIa9Jl77cgkBSbs6fMTUKaQRyBHc
J8ERlW/6tN9tyzXQwzTKSfeaMc1j4PQ+5yjTBRMJL/Y6ENQ5CmzJg1CJjnjU3jYi
6zasnLZpa1SNGs0RENfQM4DNB8yf5BCIhkKzOksWXD9RrK4mhrbFECjkHrgyAdRf
9mKXAXGXNtkCHYtsUWZ4uNAmGO+Jg61jF8Hi9mj/prfbCt8tQFQCzsqmbj1ZUeff
WzQfXacbr5mOeA1uPynn5tVkfWBU76HqLN9HT0F3e/s+cAl34g2DKjsGK3AugF4K
8ZTxt3R0MmP7ddrLG47nvvWZpt2wAMgzOmYn7QCRZIbjiHGUoQDMEkSOrYhKuDOt
F92/hOJ2YCUs7Z7imBZ31oczmWoS1yfKcb1DGKMoOPcCCyBUCDE3m1DeoaQ7oD5A
XUacEoGHtv8TTAtd0iNnaQNHgRn5UnX/KB33hG0sxHA=
`pragma protect end_protected
