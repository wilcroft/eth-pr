// eth4to1.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module eth4to1 (
		input  wire        clk_clk,                     //             clk.clk
		output wire        clk_312_out_clk_clk,         // clk_312_out_clk.clk
		output wire [63:0] eth_outstream_data,          //   eth_outstream.data
		input  wire        eth_outstream_ready,         //                .ready
		output wire        eth_outstream_valid,         //                .valid
		output wire        eth_outstream_endofpacket,   //                .endofpacket
		output wire        eth_outstream_startofpacket, //                .startofpacket
		output wire [5:0]  eth_outstream_channel,       //                .channel
		input  wire [7:0]  eth_tagstream_data,          //   eth_tagstream.data
		output wire        eth_tagstream_ready,         //                .ready
		input  wire        eth_tagstream_valid,         //                .valid
		input  wire        reset_reset_n,               //           reset.reset_n
		input  wire [71:0] xgmii_rx_data_0_data,        // xgmii_rx_data_0.data
		input  wire [71:0] xgmii_rx_data_1_data,        // xgmii_rx_data_1.data
		input  wire [71:0] xgmii_rx_data_2_data,        // xgmii_rx_data_2.data
		input  wire [71:0] xgmii_rx_data_3_data,        // xgmii_rx_data_3.data
		output wire [71:0] xgmii_tx_data_0_data,        // xgmii_tx_data_0.data
		output wire [71:0] xgmii_tx_data_1_data,        // xgmii_tx_data_1.data
		output wire [71:0] xgmii_tx_data_2_data,        // xgmii_tx_data_2.data
		output wire [71:0] xgmii_tx_data_3_data         // xgmii_tx_data_3.data
	);

	wire         demultiplexer_0_out0_valid;                // demultiplexer_0:out0_valid -> mac_0:tx_st_fifo_in_valid
	wire  [63:0] demultiplexer_0_out0_data;                 // demultiplexer_0:out0_data -> mac_0:tx_st_fifo_in_data
	wire         demultiplexer_0_out0_ready;                // mac_0:tx_st_fifo_in_ready -> demultiplexer_0:out0_ready
	wire         demultiplexer_0_out0_startofpacket;        // demultiplexer_0:out0_startofpacket -> mac_0:tx_st_fifo_in_startofpacket
	wire         demultiplexer_0_out0_endofpacket;          // demultiplexer_0:out0_endofpacket -> mac_0:tx_st_fifo_in_endofpacket
	wire         demultiplexer_0_out0_error;                // demultiplexer_0:out0_error -> mac_0:tx_st_fifo_in_error
	wire   [2:0] demultiplexer_0_out0_empty;                // demultiplexer_0:out0_empty -> mac_0:tx_st_fifo_in_empty
	wire         demultiplexer_0_out1_valid;                // demultiplexer_0:out1_valid -> mac_1:tx_st_fifo_in_valid
	wire  [63:0] demultiplexer_0_out1_data;                 // demultiplexer_0:out1_data -> mac_1:tx_st_fifo_in_data
	wire         demultiplexer_0_out1_ready;                // mac_1:tx_st_fifo_in_ready -> demultiplexer_0:out1_ready
	wire         demultiplexer_0_out1_startofpacket;        // demultiplexer_0:out1_startofpacket -> mac_1:tx_st_fifo_in_startofpacket
	wire         demultiplexer_0_out1_endofpacket;          // demultiplexer_0:out1_endofpacket -> mac_1:tx_st_fifo_in_endofpacket
	wire         demultiplexer_0_out1_error;                // demultiplexer_0:out1_error -> mac_1:tx_st_fifo_in_error
	wire   [2:0] demultiplexer_0_out1_empty;                // demultiplexer_0:out1_empty -> mac_1:tx_st_fifo_in_empty
	wire         demultiplexer_0_out2_valid;                // demultiplexer_0:out2_valid -> mac_2:tx_st_fifo_in_valid
	wire  [63:0] demultiplexer_0_out2_data;                 // demultiplexer_0:out2_data -> mac_2:tx_st_fifo_in_data
	wire         demultiplexer_0_out2_ready;                // mac_2:tx_st_fifo_in_ready -> demultiplexer_0:out2_ready
	wire         demultiplexer_0_out2_startofpacket;        // demultiplexer_0:out2_startofpacket -> mac_2:tx_st_fifo_in_startofpacket
	wire         demultiplexer_0_out2_endofpacket;          // demultiplexer_0:out2_endofpacket -> mac_2:tx_st_fifo_in_endofpacket
	wire         demultiplexer_0_out2_error;                // demultiplexer_0:out2_error -> mac_2:tx_st_fifo_in_error
	wire   [2:0] demultiplexer_0_out2_empty;                // demultiplexer_0:out2_empty -> mac_2:tx_st_fifo_in_empty
	wire         demultiplexer_0_out3_valid;                // demultiplexer_0:out3_valid -> mac_3:tx_st_fifo_in_valid
	wire  [63:0] demultiplexer_0_out3_data;                 // demultiplexer_0:out3_data -> mac_3:tx_st_fifo_in_data
	wire         demultiplexer_0_out3_ready;                // mac_3:tx_st_fifo_in_ready -> demultiplexer_0:out3_ready
	wire         demultiplexer_0_out3_startofpacket;        // demultiplexer_0:out3_startofpacket -> mac_3:tx_st_fifo_in_startofpacket
	wire         demultiplexer_0_out3_endofpacket;          // demultiplexer_0:out3_endofpacket -> mac_3:tx_st_fifo_in_endofpacket
	wire         demultiplexer_0_out3_error;                // demultiplexer_0:out3_error -> mac_3:tx_st_fifo_in_error
	wire   [2:0] demultiplexer_0_out3_empty;                // demultiplexer_0:out3_empty -> mac_3:tx_st_fifo_in_empty
	wire         mac_0_rx_st_fifo_out_valid;                // mac_0:rx_st_fifo_out_valid -> multiplexer_0:in0_valid
	wire  [63:0] mac_0_rx_st_fifo_out_data;                 // mac_0:rx_st_fifo_out_data -> multiplexer_0:in0_data
	wire         mac_0_rx_st_fifo_out_ready;                // multiplexer_0:in0_ready -> mac_0:rx_st_fifo_out_ready
	wire         mac_0_rx_st_fifo_out_startofpacket;        // mac_0:rx_st_fifo_out_startofpacket -> multiplexer_0:in0_startofpacket
	wire         mac_0_rx_st_fifo_out_endofpacket;          // mac_0:rx_st_fifo_out_endofpacket -> multiplexer_0:in0_endofpacket
	wire   [5:0] mac_0_rx_st_fifo_out_error;                // mac_0:rx_st_fifo_out_error -> multiplexer_0:in0_error
	wire   [2:0] mac_0_rx_st_fifo_out_empty;                // mac_0:rx_st_fifo_out_empty -> multiplexer_0:in0_empty
	wire         mac_1_rx_st_fifo_out_valid;                // mac_1:rx_st_fifo_out_valid -> multiplexer_0:in1_valid
	wire  [63:0] mac_1_rx_st_fifo_out_data;                 // mac_1:rx_st_fifo_out_data -> multiplexer_0:in1_data
	wire         mac_1_rx_st_fifo_out_ready;                // multiplexer_0:in1_ready -> mac_1:rx_st_fifo_out_ready
	wire         mac_1_rx_st_fifo_out_startofpacket;        // mac_1:rx_st_fifo_out_startofpacket -> multiplexer_0:in1_startofpacket
	wire         mac_1_rx_st_fifo_out_endofpacket;          // mac_1:rx_st_fifo_out_endofpacket -> multiplexer_0:in1_endofpacket
	wire   [5:0] mac_1_rx_st_fifo_out_error;                // mac_1:rx_st_fifo_out_error -> multiplexer_0:in1_error
	wire   [2:0] mac_1_rx_st_fifo_out_empty;                // mac_1:rx_st_fifo_out_empty -> multiplexer_0:in1_empty
	wire         mac_2_rx_st_fifo_out_valid;                // mac_2:rx_st_fifo_out_valid -> multiplexer_0:in2_valid
	wire  [63:0] mac_2_rx_st_fifo_out_data;                 // mac_2:rx_st_fifo_out_data -> multiplexer_0:in2_data
	wire         mac_2_rx_st_fifo_out_ready;                // multiplexer_0:in2_ready -> mac_2:rx_st_fifo_out_ready
	wire         mac_2_rx_st_fifo_out_startofpacket;        // mac_2:rx_st_fifo_out_startofpacket -> multiplexer_0:in2_startofpacket
	wire         mac_2_rx_st_fifo_out_endofpacket;          // mac_2:rx_st_fifo_out_endofpacket -> multiplexer_0:in2_endofpacket
	wire   [5:0] mac_2_rx_st_fifo_out_error;                // mac_2:rx_st_fifo_out_error -> multiplexer_0:in2_error
	wire   [2:0] mac_2_rx_st_fifo_out_empty;                // mac_2:rx_st_fifo_out_empty -> multiplexer_0:in2_empty
	wire         mac_3_rx_st_fifo_out_valid;                // mac_3:rx_st_fifo_out_valid -> multiplexer_0:in3_valid
	wire  [63:0] mac_3_rx_st_fifo_out_data;                 // mac_3:rx_st_fifo_out_data -> multiplexer_0:in3_data
	wire         mac_3_rx_st_fifo_out_ready;                // multiplexer_0:in3_ready -> mac_3:rx_st_fifo_out_ready
	wire         mac_3_rx_st_fifo_out_startofpacket;        // mac_3:rx_st_fifo_out_startofpacket -> multiplexer_0:in3_startofpacket
	wire         mac_3_rx_st_fifo_out_endofpacket;          // mac_3:rx_st_fifo_out_endofpacket -> multiplexer_0:in3_endofpacket
	wire   [5:0] mac_3_rx_st_fifo_out_error;                // mac_3:rx_st_fifo_out_error -> multiplexer_0:in3_error
	wire   [2:0] mac_3_rx_st_fifo_out_empty;                // mac_3:rx_st_fifo_out_empty -> multiplexer_0:in3_empty
	wire         multiplexer_0_out_valid;                   // multiplexer_0:out_valid -> avalon_st_adapter:in_0_valid
	wire  [63:0] multiplexer_0_out_data;                    // multiplexer_0:out_data -> avalon_st_adapter:in_0_data
	wire         multiplexer_0_out_ready;                   // avalon_st_adapter:in_0_ready -> multiplexer_0:out_ready
	wire   [1:0] multiplexer_0_out_channel;                 // multiplexer_0:out_channel -> avalon_st_adapter:in_0_channel
	wire         multiplexer_0_out_startofpacket;           // multiplexer_0:out_startofpacket -> avalon_st_adapter:in_0_startofpacket
	wire         multiplexer_0_out_endofpacket;             // multiplexer_0:out_endofpacket -> avalon_st_adapter:in_0_endofpacket
	wire   [5:0] multiplexer_0_out_error;                   // multiplexer_0:out_error -> avalon_st_adapter:in_0_error
	wire   [2:0] multiplexer_0_out_empty;                   // multiplexer_0:out_empty -> avalon_st_adapter:in_0_empty
	wire         avalon_st_adapter_out_0_valid;             // avalon_st_adapter:out_0_valid -> eth:instream_valid
	wire  [63:0] avalon_st_adapter_out_0_data;              // avalon_st_adapter:out_0_data -> eth:instream_data
	wire         avalon_st_adapter_out_0_ready;             // eth:instream_ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;     // avalon_st_adapter:out_0_startofpacket -> eth:instream_sop
	wire         avalon_st_adapter_out_0_endofpacket;       // avalon_st_adapter:out_0_endofpacket -> eth:instream_eop
	wire         eth_sendstream_valid;                      // eth:sendstream_valid -> avalon_st_adapter_001:in_0_valid
	wire  [63:0] eth_sendstream_data;                       // eth:sendstream_data -> avalon_st_adapter_001:in_0_data
	wire         eth_sendstream_ready;                      // avalon_st_adapter_001:in_0_ready -> eth:sendstream_ready
	wire   [1:0] eth_sendstream_channel;                    // eth:sendstream_channel -> avalon_st_adapter_001:in_0_channel
	wire         eth_sendstream_startofpacket;              // eth:sendstream_sop -> avalon_st_adapter_001:in_0_startofpacket
	wire         eth_sendstream_endofpacket;                // eth:sendstream_eop -> avalon_st_adapter_001:in_0_endofpacket
	wire         avalon_st_adapter_001_out_0_valid;         // avalon_st_adapter_001:out_0_valid -> demultiplexer_0:in_valid
	wire  [63:0] avalon_st_adapter_001_out_0_data;          // avalon_st_adapter_001:out_0_data -> demultiplexer_0:in_data
	wire         avalon_st_adapter_001_out_0_ready;         // demultiplexer_0:in_ready -> avalon_st_adapter_001:out_0_ready
	wire   [1:0] avalon_st_adapter_001_out_0_channel;       // avalon_st_adapter_001:out_0_channel -> demultiplexer_0:in_channel
	wire         avalon_st_adapter_001_out_0_startofpacket; // avalon_st_adapter_001:out_0_startofpacket -> demultiplexer_0:in_startofpacket
	wire         avalon_st_adapter_001_out_0_endofpacket;   // avalon_st_adapter_001:out_0_endofpacket -> demultiplexer_0:in_endofpacket
	wire   [0:0] avalon_st_adapter_001_out_0_error;         // avalon_st_adapter_001:out_0_error -> demultiplexer_0:in_error
	wire   [2:0] avalon_st_adapter_001_out_0_empty;         // avalon_st_adapter_001:out_0_empty -> demultiplexer_0:in_empty
	wire         rst_controller_reset_out_reset;            // rst_controller:reset_out -> [avalon_st_adapter:in_rst_0_reset, avalon_st_adapter_001:in_rst_0_reset, demultiplexer_0:reset_n, eth:reset, multiplexer_0:reset_n]
	wire         rst_controller_001_reset_out_reset;        // rst_controller_001:reset_out -> [mac_0:rst_in_reset_reset, mac_1:rst_in_reset_reset, mac_2:rst_in_reset_reset, mac_3:rst_in_reset_reset]

	eth4to1_demultiplexer_0 demultiplexer_0 (
		.clk                (clk_312_out_clk_clk),                       //   clk.clk
		.reset_n            (~rst_controller_reset_out_reset),           // reset.reset_n
		.in_data            (avalon_st_adapter_001_out_0_data),          //    in.data
		.in_valid           (avalon_st_adapter_001_out_0_valid),         //      .valid
		.in_ready           (avalon_st_adapter_001_out_0_ready),         //      .ready
		.in_startofpacket   (avalon_st_adapter_001_out_0_startofpacket), //      .startofpacket
		.in_endofpacket     (avalon_st_adapter_001_out_0_endofpacket),   //      .endofpacket
		.in_empty           (avalon_st_adapter_001_out_0_empty),         //      .empty
		.in_error           (avalon_st_adapter_001_out_0_error),         //      .error
		.in_channel         (avalon_st_adapter_001_out_0_channel),       //      .channel
		.out0_data          (demultiplexer_0_out0_data),                 //  out0.data
		.out0_valid         (demultiplexer_0_out0_valid),                //      .valid
		.out0_ready         (demultiplexer_0_out0_ready),                //      .ready
		.out0_startofpacket (demultiplexer_0_out0_startofpacket),        //      .startofpacket
		.out0_endofpacket   (demultiplexer_0_out0_endofpacket),          //      .endofpacket
		.out0_empty         (demultiplexer_0_out0_empty),                //      .empty
		.out0_error         (demultiplexer_0_out0_error),                //      .error
		.out1_data          (demultiplexer_0_out1_data),                 //  out1.data
		.out1_valid         (demultiplexer_0_out1_valid),                //      .valid
		.out1_ready         (demultiplexer_0_out1_ready),                //      .ready
		.out1_startofpacket (demultiplexer_0_out1_startofpacket),        //      .startofpacket
		.out1_endofpacket   (demultiplexer_0_out1_endofpacket),          //      .endofpacket
		.out1_empty         (demultiplexer_0_out1_empty),                //      .empty
		.out1_error         (demultiplexer_0_out1_error),                //      .error
		.out2_data          (demultiplexer_0_out2_data),                 //  out2.data
		.out2_valid         (demultiplexer_0_out2_valid),                //      .valid
		.out2_ready         (demultiplexer_0_out2_ready),                //      .ready
		.out2_startofpacket (demultiplexer_0_out2_startofpacket),        //      .startofpacket
		.out2_endofpacket   (demultiplexer_0_out2_endofpacket),          //      .endofpacket
		.out2_empty         (demultiplexer_0_out2_empty),                //      .empty
		.out2_error         (demultiplexer_0_out2_error),                //      .error
		.out3_data          (demultiplexer_0_out3_data),                 //  out3.data
		.out3_valid         (demultiplexer_0_out3_valid),                //      .valid
		.out3_ready         (demultiplexer_0_out3_ready),                //      .ready
		.out3_startofpacket (demultiplexer_0_out3_startofpacket),        //      .startofpacket
		.out3_endofpacket   (demultiplexer_0_out3_endofpacket),          //      .endofpacket
		.out3_empty         (demultiplexer_0_out3_empty),                //      .empty
		.out3_error         (demultiplexer_0_out3_error)                 //      .error
	);

	eth4to1_eth eth (
		.reset              (rst_controller_reset_out_reset),        //      reset.reset
		.clock              (clk_312_out_clk_clk),                   //      clock.clk
		.outstream_data     (eth_outstream_data),                    //  outstream.data
		.outstream_ready    (eth_outstream_ready),                   //           .ready
		.outstream_valid    (eth_outstream_valid),                   //           .valid
		.outstream_eop      (eth_outstream_endofpacket),             //           .endofpacket
		.outstream_sop      (eth_outstream_startofpacket),           //           .startofpacket
		.outstream_channel  (eth_outstream_channel),                 //           .channel
		.sendstream_data    (eth_sendstream_data),                   // sendstream.data
		.sendstream_valid   (eth_sendstream_valid),                  //           .valid
		.sendstream_ready   (eth_sendstream_ready),                  //           .ready
		.sendstream_eop     (eth_sendstream_endofpacket),            //           .endofpacket
		.sendstream_sop     (eth_sendstream_startofpacket),          //           .startofpacket
		.sendstream_channel (eth_sendstream_channel),                //           .channel
		.tagstream_data     (eth_tagstream_data),                    //  tagstream.data
		.tagstream_ready    (eth_tagstream_ready),                   //           .ready
		.tagstream_valid    (eth_tagstream_valid),                   //           .valid
		.instream_data      (avalon_st_adapter_out_0_data),          //   instream.data
		.instream_eop       (avalon_st_adapter_out_0_endofpacket),   //           .endofpacket
		.instream_sop       (avalon_st_adapter_out_0_startofpacket), //           .startofpacket
		.instream_ready     (avalon_st_adapter_out_0_ready),         //           .ready
		.instream_valid     (avalon_st_adapter_out_0_valid)          //           .valid
	);

	eth4to1_mac_0 mac_0 (
		.clk_156_in_clk_clk                     (clk_clk),                            //                    clk_156_in_clk.clk
		.clk_312_in_clk_clk                     (clk_312_out_clk_clk),                //                    clk_312_in_clk.clk
		.mac10g_avalon_st_pause_data            (),                                   //            mac10g_avalon_st_pause.data
		.mac10g_avalon_st_rxstatus_valid        (),                                   //         mac10g_avalon_st_rxstatus.valid
		.mac10g_avalon_st_rxstatus_data         (),                                   //                                  .data
		.mac10g_avalon_st_rxstatus_error        (),                                   //                                  .error
		.mac10g_avalon_st_txstatus_data         (),                                   //         mac10g_avalon_st_txstatus.data
		.mac10g_avalon_st_txstatus_valid        (),                                   //                                  .valid
		.mac10g_avalon_st_txstatus_error        (),                                   //                                  .error
		.mac10g_csr_address                     (),                                   //                        mac10g_csr.address
		.mac10g_csr_waitrequest                 (),                                   //                                  .waitrequest
		.mac10g_csr_read                        (),                                   //                                  .read
		.mac10g_csr_readdata                    (),                                   //                                  .readdata
		.mac10g_csr_write                       (),                                   //                                  .write
		.mac10g_csr_writedata                   (),                                   //                                  .writedata
		.mac10g_link_fault_status_xgmii_rx_data (),                                   // mac10g_link_fault_status_xgmii_rx.data
		.mac10g_xgmii_rx_data                   (xgmii_rx_data_0_data),               //                   mac10g_xgmii_rx.data
		.mac10g_xgmii_tx_data                   (xgmii_tx_data_0_data),               //                   mac10g_xgmii_tx.data
		.rst_in_reset_reset                     (rst_controller_001_reset_out_reset), //                      rst_in_reset.reset
		.rx_st_fifo_out_data                    (mac_0_rx_st_fifo_out_data),          //                    rx_st_fifo_out.data
		.rx_st_fifo_out_valid                   (mac_0_rx_st_fifo_out_valid),         //                                  .valid
		.rx_st_fifo_out_ready                   (mac_0_rx_st_fifo_out_ready),         //                                  .ready
		.rx_st_fifo_out_startofpacket           (mac_0_rx_st_fifo_out_startofpacket), //                                  .startofpacket
		.rx_st_fifo_out_endofpacket             (mac_0_rx_st_fifo_out_endofpacket),   //                                  .endofpacket
		.rx_st_fifo_out_empty                   (mac_0_rx_st_fifo_out_empty),         //                                  .empty
		.rx_st_fifo_out_error                   (mac_0_rx_st_fifo_out_error),         //                                  .error
		.tx_st_fifo_in_data                     (demultiplexer_0_out0_data),          //                     tx_st_fifo_in.data
		.tx_st_fifo_in_valid                    (demultiplexer_0_out0_valid),         //                                  .valid
		.tx_st_fifo_in_ready                    (demultiplexer_0_out0_ready),         //                                  .ready
		.tx_st_fifo_in_startofpacket            (demultiplexer_0_out0_startofpacket), //                                  .startofpacket
		.tx_st_fifo_in_endofpacket              (demultiplexer_0_out0_endofpacket),   //                                  .endofpacket
		.tx_st_fifo_in_empty                    (demultiplexer_0_out0_empty),         //                                  .empty
		.tx_st_fifo_in_error                    (demultiplexer_0_out0_error)          //                                  .error
	);

	eth4to1_mac_1 mac_1 (
		.clk_156_in_clk_clk                     (clk_clk),                            //                    clk_156_in_clk.clk
		.clk_312_in_clk_clk                     (clk_312_out_clk_clk),                //                    clk_312_in_clk.clk
		.mac10g_avalon_st_pause_data            (),                                   //            mac10g_avalon_st_pause.data
		.mac10g_avalon_st_rxstatus_valid        (),                                   //         mac10g_avalon_st_rxstatus.valid
		.mac10g_avalon_st_rxstatus_data         (),                                   //                                  .data
		.mac10g_avalon_st_rxstatus_error        (),                                   //                                  .error
		.mac10g_avalon_st_txstatus_data         (),                                   //         mac10g_avalon_st_txstatus.data
		.mac10g_avalon_st_txstatus_valid        (),                                   //                                  .valid
		.mac10g_avalon_st_txstatus_error        (),                                   //                                  .error
		.mac10g_csr_address                     (),                                   //                        mac10g_csr.address
		.mac10g_csr_waitrequest                 (),                                   //                                  .waitrequest
		.mac10g_csr_read                        (),                                   //                                  .read
		.mac10g_csr_readdata                    (),                                   //                                  .readdata
		.mac10g_csr_write                       (),                                   //                                  .write
		.mac10g_csr_writedata                   (),                                   //                                  .writedata
		.mac10g_link_fault_status_xgmii_rx_data (),                                   // mac10g_link_fault_status_xgmii_rx.data
		.mac10g_xgmii_rx_data                   (xgmii_rx_data_1_data),               //                   mac10g_xgmii_rx.data
		.mac10g_xgmii_tx_data                   (xgmii_tx_data_1_data),               //                   mac10g_xgmii_tx.data
		.rst_in_reset_reset                     (rst_controller_001_reset_out_reset), //                      rst_in_reset.reset
		.rx_st_fifo_out_data                    (mac_1_rx_st_fifo_out_data),          //                    rx_st_fifo_out.data
		.rx_st_fifo_out_valid                   (mac_1_rx_st_fifo_out_valid),         //                                  .valid
		.rx_st_fifo_out_ready                   (mac_1_rx_st_fifo_out_ready),         //                                  .ready
		.rx_st_fifo_out_startofpacket           (mac_1_rx_st_fifo_out_startofpacket), //                                  .startofpacket
		.rx_st_fifo_out_endofpacket             (mac_1_rx_st_fifo_out_endofpacket),   //                                  .endofpacket
		.rx_st_fifo_out_empty                   (mac_1_rx_st_fifo_out_empty),         //                                  .empty
		.rx_st_fifo_out_error                   (mac_1_rx_st_fifo_out_error),         //                                  .error
		.tx_st_fifo_in_data                     (demultiplexer_0_out1_data),          //                     tx_st_fifo_in.data
		.tx_st_fifo_in_valid                    (demultiplexer_0_out1_valid),         //                                  .valid
		.tx_st_fifo_in_ready                    (demultiplexer_0_out1_ready),         //                                  .ready
		.tx_st_fifo_in_startofpacket            (demultiplexer_0_out1_startofpacket), //                                  .startofpacket
		.tx_st_fifo_in_endofpacket              (demultiplexer_0_out1_endofpacket),   //                                  .endofpacket
		.tx_st_fifo_in_empty                    (demultiplexer_0_out1_empty),         //                                  .empty
		.tx_st_fifo_in_error                    (demultiplexer_0_out1_error)          //                                  .error
	);

	eth4to1_mac_2 mac_2 (
		.clk_156_in_clk_clk                     (clk_clk),                            //                    clk_156_in_clk.clk
		.clk_312_in_clk_clk                     (clk_312_out_clk_clk),                //                    clk_312_in_clk.clk
		.mac10g_avalon_st_pause_data            (),                                   //            mac10g_avalon_st_pause.data
		.mac10g_avalon_st_rxstatus_valid        (),                                   //         mac10g_avalon_st_rxstatus.valid
		.mac10g_avalon_st_rxstatus_data         (),                                   //                                  .data
		.mac10g_avalon_st_rxstatus_error        (),                                   //                                  .error
		.mac10g_avalon_st_txstatus_data         (),                                   //         mac10g_avalon_st_txstatus.data
		.mac10g_avalon_st_txstatus_valid        (),                                   //                                  .valid
		.mac10g_avalon_st_txstatus_error        (),                                   //                                  .error
		.mac10g_csr_address                     (),                                   //                        mac10g_csr.address
		.mac10g_csr_waitrequest                 (),                                   //                                  .waitrequest
		.mac10g_csr_read                        (),                                   //                                  .read
		.mac10g_csr_readdata                    (),                                   //                                  .readdata
		.mac10g_csr_write                       (),                                   //                                  .write
		.mac10g_csr_writedata                   (),                                   //                                  .writedata
		.mac10g_link_fault_status_xgmii_rx_data (),                                   // mac10g_link_fault_status_xgmii_rx.data
		.mac10g_xgmii_rx_data                   (xgmii_rx_data_2_data),               //                   mac10g_xgmii_rx.data
		.mac10g_xgmii_tx_data                   (xgmii_tx_data_2_data),               //                   mac10g_xgmii_tx.data
		.rst_in_reset_reset                     (rst_controller_001_reset_out_reset), //                      rst_in_reset.reset
		.rx_st_fifo_out_data                    (mac_2_rx_st_fifo_out_data),          //                    rx_st_fifo_out.data
		.rx_st_fifo_out_valid                   (mac_2_rx_st_fifo_out_valid),         //                                  .valid
		.rx_st_fifo_out_ready                   (mac_2_rx_st_fifo_out_ready),         //                                  .ready
		.rx_st_fifo_out_startofpacket           (mac_2_rx_st_fifo_out_startofpacket), //                                  .startofpacket
		.rx_st_fifo_out_endofpacket             (mac_2_rx_st_fifo_out_endofpacket),   //                                  .endofpacket
		.rx_st_fifo_out_empty                   (mac_2_rx_st_fifo_out_empty),         //                                  .empty
		.rx_st_fifo_out_error                   (mac_2_rx_st_fifo_out_error),         //                                  .error
		.tx_st_fifo_in_data                     (demultiplexer_0_out2_data),          //                     tx_st_fifo_in.data
		.tx_st_fifo_in_valid                    (demultiplexer_0_out2_valid),         //                                  .valid
		.tx_st_fifo_in_ready                    (demultiplexer_0_out2_ready),         //                                  .ready
		.tx_st_fifo_in_startofpacket            (demultiplexer_0_out2_startofpacket), //                                  .startofpacket
		.tx_st_fifo_in_endofpacket              (demultiplexer_0_out2_endofpacket),   //                                  .endofpacket
		.tx_st_fifo_in_empty                    (demultiplexer_0_out2_empty),         //                                  .empty
		.tx_st_fifo_in_error                    (demultiplexer_0_out2_error)          //                                  .error
	);

	eth4to1_mac_3 mac_3 (
		.clk_156_in_clk_clk                     (clk_clk),                            //                    clk_156_in_clk.clk
		.clk_312_in_clk_clk                     (clk_312_out_clk_clk),                //                    clk_312_in_clk.clk
		.mac10g_avalon_st_pause_data            (),                                   //            mac10g_avalon_st_pause.data
		.mac10g_avalon_st_rxstatus_valid        (),                                   //         mac10g_avalon_st_rxstatus.valid
		.mac10g_avalon_st_rxstatus_data         (),                                   //                                  .data
		.mac10g_avalon_st_rxstatus_error        (),                                   //                                  .error
		.mac10g_avalon_st_txstatus_data         (),                                   //         mac10g_avalon_st_txstatus.data
		.mac10g_avalon_st_txstatus_valid        (),                                   //                                  .valid
		.mac10g_avalon_st_txstatus_error        (),                                   //                                  .error
		.mac10g_csr_address                     (),                                   //                        mac10g_csr.address
		.mac10g_csr_waitrequest                 (),                                   //                                  .waitrequest
		.mac10g_csr_read                        (),                                   //                                  .read
		.mac10g_csr_readdata                    (),                                   //                                  .readdata
		.mac10g_csr_write                       (),                                   //                                  .write
		.mac10g_csr_writedata                   (),                                   //                                  .writedata
		.mac10g_link_fault_status_xgmii_rx_data (),                                   // mac10g_link_fault_status_xgmii_rx.data
		.mac10g_xgmii_rx_data                   (xgmii_rx_data_3_data),               //                   mac10g_xgmii_rx.data
		.mac10g_xgmii_tx_data                   (xgmii_tx_data_3_data),               //                   mac10g_xgmii_tx.data
		.rst_in_reset_reset                     (rst_controller_001_reset_out_reset), //                      rst_in_reset.reset
		.rx_st_fifo_out_data                    (mac_3_rx_st_fifo_out_data),          //                    rx_st_fifo_out.data
		.rx_st_fifo_out_valid                   (mac_3_rx_st_fifo_out_valid),         //                                  .valid
		.rx_st_fifo_out_ready                   (mac_3_rx_st_fifo_out_ready),         //                                  .ready
		.rx_st_fifo_out_startofpacket           (mac_3_rx_st_fifo_out_startofpacket), //                                  .startofpacket
		.rx_st_fifo_out_endofpacket             (mac_3_rx_st_fifo_out_endofpacket),   //                                  .endofpacket
		.rx_st_fifo_out_empty                   (mac_3_rx_st_fifo_out_empty),         //                                  .empty
		.rx_st_fifo_out_error                   (mac_3_rx_st_fifo_out_error),         //                                  .error
		.tx_st_fifo_in_data                     (demultiplexer_0_out3_data),          //                     tx_st_fifo_in.data
		.tx_st_fifo_in_valid                    (demultiplexer_0_out3_valid),         //                                  .valid
		.tx_st_fifo_in_ready                    (demultiplexer_0_out3_ready),         //                                  .ready
		.tx_st_fifo_in_startofpacket            (demultiplexer_0_out3_startofpacket), //                                  .startofpacket
		.tx_st_fifo_in_endofpacket              (demultiplexer_0_out3_endofpacket),   //                                  .endofpacket
		.tx_st_fifo_in_empty                    (demultiplexer_0_out3_empty),         //                                  .empty
		.tx_st_fifo_in_error                    (demultiplexer_0_out3_error)          //                                  .error
	);

	eth4to1_multiplexer_0 multiplexer_0 (
		.clk               (clk_312_out_clk_clk),                //   clk.clk
		.reset_n           (~rst_controller_reset_out_reset),    // reset.reset_n
		.out_data          (multiplexer_0_out_data),             //   out.data
		.out_valid         (multiplexer_0_out_valid),            //      .valid
		.out_ready         (multiplexer_0_out_ready),            //      .ready
		.out_startofpacket (multiplexer_0_out_startofpacket),    //      .startofpacket
		.out_endofpacket   (multiplexer_0_out_endofpacket),      //      .endofpacket
		.out_empty         (multiplexer_0_out_empty),            //      .empty
		.out_error         (multiplexer_0_out_error),            //      .error
		.out_channel       (multiplexer_0_out_channel),          //      .channel
		.in0_data          (mac_0_rx_st_fifo_out_data),          //   in0.data
		.in0_valid         (mac_0_rx_st_fifo_out_valid),         //      .valid
		.in0_ready         (mac_0_rx_st_fifo_out_ready),         //      .ready
		.in0_startofpacket (mac_0_rx_st_fifo_out_startofpacket), //      .startofpacket
		.in0_endofpacket   (mac_0_rx_st_fifo_out_endofpacket),   //      .endofpacket
		.in0_empty         (mac_0_rx_st_fifo_out_empty),         //      .empty
		.in0_error         (mac_0_rx_st_fifo_out_error),         //      .error
		.in1_data          (mac_1_rx_st_fifo_out_data),          //   in1.data
		.in1_valid         (mac_1_rx_st_fifo_out_valid),         //      .valid
		.in1_ready         (mac_1_rx_st_fifo_out_ready),         //      .ready
		.in1_startofpacket (mac_1_rx_st_fifo_out_startofpacket), //      .startofpacket
		.in1_endofpacket   (mac_1_rx_st_fifo_out_endofpacket),   //      .endofpacket
		.in1_empty         (mac_1_rx_st_fifo_out_empty),         //      .empty
		.in1_error         (mac_1_rx_st_fifo_out_error),         //      .error
		.in2_data          (mac_2_rx_st_fifo_out_data),          //   in2.data
		.in2_valid         (mac_2_rx_st_fifo_out_valid),         //      .valid
		.in2_ready         (mac_2_rx_st_fifo_out_ready),         //      .ready
		.in2_startofpacket (mac_2_rx_st_fifo_out_startofpacket), //      .startofpacket
		.in2_endofpacket   (mac_2_rx_st_fifo_out_endofpacket),   //      .endofpacket
		.in2_empty         (mac_2_rx_st_fifo_out_empty),         //      .empty
		.in2_error         (mac_2_rx_st_fifo_out_error),         //      .error
		.in3_data          (mac_3_rx_st_fifo_out_data),          //   in3.data
		.in3_valid         (mac_3_rx_st_fifo_out_valid),         //      .valid
		.in3_ready         (mac_3_rx_st_fifo_out_ready),         //      .ready
		.in3_startofpacket (mac_3_rx_st_fifo_out_startofpacket), //      .startofpacket
		.in3_endofpacket   (mac_3_rx_st_fifo_out_endofpacket),   //      .endofpacket
		.in3_empty         (mac_3_rx_st_fifo_out_empty),         //      .empty
		.in3_error         (mac_3_rx_st_fifo_out_error)          //      .error
	);

	eth4to1_pll_0 pll_0 (
		.refclk   (clk_clk),             //  refclk.clk
		.rst      (~reset_reset_n),      //   reset.reset
		.outclk_0 (clk_312_out_clk_clk), // outclk0.clk
		.locked   ()                     // (terminated)
	);

	eth4to1_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (64),
		.inChannelWidth  (2),
		.inErrorWidth    (6),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (64),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (clk_312_out_clk_clk),                   // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),        // in_rst_0.reset
		.in_0_data           (multiplexer_0_out_data),                //     in_0.data
		.in_0_valid          (multiplexer_0_out_valid),               //         .valid
		.in_0_ready          (multiplexer_0_out_ready),               //         .ready
		.in_0_startofpacket  (multiplexer_0_out_startofpacket),       //         .startofpacket
		.in_0_endofpacket    (multiplexer_0_out_endofpacket),         //         .endofpacket
		.in_0_empty          (multiplexer_0_out_empty),               //         .empty
		.in_0_error          (multiplexer_0_out_error),               //         .error
		.in_0_channel        (multiplexer_0_out_channel),             //         .channel
		.out_0_data          (avalon_st_adapter_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket)    //         .endofpacket
	);

	eth4to1_avalon_st_adapter_001 #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (64),
		.inChannelWidth  (2),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (64),
		.outChannelWidth (2),
		.outErrorWidth   (1),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_001 (
		.in_clk_0_clk        (clk_312_out_clk_clk),                       // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),            // in_rst_0.reset
		.in_0_data           (eth_sendstream_data),                       //     in_0.data
		.in_0_valid          (eth_sendstream_valid),                      //         .valid
		.in_0_ready          (eth_sendstream_ready),                      //         .ready
		.in_0_startofpacket  (eth_sendstream_startofpacket),              //         .startofpacket
		.in_0_endofpacket    (eth_sendstream_endofpacket),                //         .endofpacket
		.in_0_channel        (eth_sendstream_channel),                    //         .channel
		.out_0_data          (avalon_st_adapter_001_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_001_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_001_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_001_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_001_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_001_out_0_empty),         //         .empty
		.out_0_error         (avalon_st_adapter_001_out_0_error),         //         .error
		.out_0_channel       (avalon_st_adapter_001_out_0_channel)        //         .channel
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_312_out_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
