// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:34:58 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sdeW8dnNW6NHTiKPYVepTOfWkKFupj6tXoiRSbcUo4fA6KPlxiXc/jVQ1MB4bKee
df/QITFI/WqbSJ43LiYHSnG8rLPefFnchigUOUg825Ne2yAssENNV8TAgCjcQGvS
uoZSoGmkCJQSSpewIcf8OdMx0eMhQL9AUqq5/rIjtm4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28384)
AvcWmKfN8HiRINHSHCg+XGLL18FnM9xDFUAc3hNGXOAf6Ug9g1l+Qvn3XK4rXpG8
efPgpTOjgo2g03CW2YkDIcAvnaimAw9wfo35SShS1G5JRV1Aj5xTdOWM81p8XvRI
FanYd3Yvqe2HD8Pp6Wxtd2FMHMw9KG62MTbeijzLD70AAUoVNFcLBVcgOKVRKYXF
tAjmbjtKGRZ+3IKB72z0OueqBA60f2bf4hSz/TK/8TwJT2DEALsvHEcqaNek2KeT
wfrwPUIIBIDRz7O5I/M3nBy64fBzw8y0GFnZ6YN8O1whaqz1lW1Da1yeZunYYsVb
ZdC2ujtXrDm9eE03B/thKhhFAPiMjNU8lbDUO/Zt/MAyfPzpAKopXxAOv2Wu3L2P
w2m59m3oIdxZZYD1XPzNedjqLm1ruYGXHmfYnhsubZto1pqkhdGLwxI96+LyeMeY
m+qgXBkbawEPUy3UUiRv26E6PSRmxDPYi5JfY3Bdyv47yKCOtwOlQWgn0jf7Fyvb
bB7ft725edEWvPXunLqyfbFyyV0r4dvLLlg3GGiwOHFaL6khwb07uTnkww6EFHAa
QtKH8RwkB3n/RP1tl61ErUy3p/DJ43g7tGytnZb3ZYMYSF0cvvgdiJJGqSK5yWRZ
r/9k6UMWMwgQ5UJ1wTSjeCGVPw2Bu7p6JR8VZz/oMIJ0c/MG5X2RaggWOIY9/IHz
yxa3rs+kfXqhmah5rfguUY0yriGhoaiAe/xoD0SJxSHipQmDBXcaj6zw1mPTKVQC
VLSbI0Yo0ZoBBhExHzn9fJkSCpB5mH6QDT7mv/yWsU5a0FiEsByasrePt5NoyNEJ
OeucIb3s7j8W7GFot+2fJ07fcKg+2VDiUxrx8QWgmxw1MwMoeLnJ4tU3VJh9gVw+
YK37bfhX6nivHk930PbDffsikArA+wPm3sDJQw1Iq4vjQJy6QmXZvtPL0sgVNSvH
xfLHFDDm14SjKChjUozXd9JOiG9+4yyWZ7HIPh4mQwx22L+Db1pnsYo8dQGBmoVN
ogPnFNXn/Feo5acsTlyeF0U0GvLQrgDnOeYVkehHaOFF+eo5+l7QNyzWN6A6NJja
KVB995vRLAkex+q6flNKI5hu1gCdYPTbgFx6Xj2Q0r4QUuXVrxJDZIEz1ybcSqSF
T58a6QlhQKGYDzyblV4tu2SthUyJmIYU0COLAEZOWBHBS6+ItvNrXY8/Oxfga9ou
UZzrnk8GLXkT+VlbkyNhmyrOINfWpLvWk0TQQQq4YmVvkn7sKLMgyzeE5yNR6W5/
4kA/JiezHfXEK8+6RFG49ItCEYzLsLAptLhVQnpicLFeaIK01rR6Pt/tuMWuI+VU
NegICxN6+8VCzFGdKVk7Nio/d0Ak8GgyiDTP53SJtgvp1lIcXDjyiAhfio4KCLbG
bRa5VXC7jsfJfKEwnTINRABJlJqChHCbHYDo3BxS+RHqBsmO+8IcVZijik1aftLr
LQFBMgHuVjWfYYH8douwuz0Do/SxSagP5gHcdbktRcomzxQnP0Vg++HAzYM9hKzs
6AHYvoOlAb3rk9CSAvFi/Sdjc3jBJ1he/UijKb6vc/tR9vq/5o6yTGiExLyAiAeG
L8pn7KbU0uNClsdEnEKysbs8P2T6Mp7w6lFWyxYEi+vA/067KERXByVieajge8TG
BsKFbSzk3khYJljGfstY0s56Tt1AZHS5XTs07toUUPQsyKjVemZSvrhQXaiKD30E
NNbqeh5Ajtu3mUAyuwUTciAk1GWJX2BelrjJq8CAi5Bl6M1lsJCADZz1E41wSDMp
t4BRFXe3+1BbBicpXn4yq3bRCcvhB1emCfgobuIGh+5NsKSq3/tzKE69/kVI18t3
Lw2+8wrp7POiTYFcLzbSe6RUa8VK4RTbodSzfKpfy4DenY0K9T561PMA8moOCOtZ
sXScC2dlxWDa+URQXFzO3Ao6UsSr5SE6cxDGu3EUO53eDNyVLphTINmX/f5MxO4P
4Puo4EgNBtpKBSs0QukVjoCLikdLU3uYCg3zyQ/RUAGgTvL1JX/AVh4hOEJlTgcX
7jDXE9iq3P57gQxV1HaPVHWujPaBFL3X5g0CaeMaO7TthFPznK5nz3CsWWqnBEV3
TnpB4IqBVUalEyyuI00QpGcxpHQd3uPhOO49xnbmpZqPDsyZ+f1S9XJUEGGrS2e3
ke/mXeYlLVEZVxILnjuSOzbTeu8acE25VmFD0AGHwqumwoaRE9N+70Io3C3tAVht
VhndUzcSnrKG3U96imrqxibmJ5SMW5XpkQQ/fctUyT2Ln8b5/n0XqSEm8hfwk1YP
AzJbQZsoC9f+RtOaPGxwQtSQZpj9Z5TWB9GX9fIo0MsRtnFK95qT+RAU8SgF+ug1
iym21ROrS2WtCfOvpVuJXURpH//CXro/Etw06RkrTbfb+BnYH0VWBwiUHrAUbr0E
TypqP1LyTyzSne0XpTTtLaQ56YkwC59zBjDEDIViK7hXit3q1838TNISmfKrNmm7
3vYkunLCold3WKS5hDkZDGy2r29spA4rQT4VTv6IZmwQ0gqbzI5KStgyIcxKXLZ2
Kez9No13/5qFJ22pS17KUj3pwAJAN+4XUGEX/chuN22/BkQ6+GNNszOdHnZC+HME
OaQCMwkQcBTbYJIF1BmrfPzyKEA/u+HQ2+JPRzUbgbdEfDpR9OaAwJHDiUbrN4Qa
zvSkMFdk4YOQbU9z2X019Bw1qrxBtM0gaccdM6NucNJBzwDZv3/jrC+MIUrLyMfP
b4UynT+OAXZSt3MwaNhOr7dexiWaj/tOs7eg1yUgJ1bSkM7bL7XBy+1ir6AjwQCx
fCjcIaHMjVXP6yZXLphJM0vm0+6IAtvNvxJguS7l+1rH37vyi9jQqDsuwKD9Fsgc
MVHQTkJ9LEss6PxxkJjtei9Ugiv2DKW5oxFINWV79dM0lu3V4T5uraII1GqWw0VI
spfYf7eUCnh9avky+0AiGwXWX+wjxVEPGzOCZ+6B+F0iUcHeYjEwXK/hNnnfgu0w
B6DqLJ8DUsdYoReK5O1LDtTFB28n3znYxqiHLx+2AmQdU6Y+SJED/059YuImOHbu
ZKiQEP+4auu5Dd8xwBznrjN8gVjBj0zQJn4w6LNXiZc9B6zbjiWyuzpelsDT5y9X
BZx4Nbwl+fC77+dzFRM+p1SWtGbWR4DoYA/MN+GNt9cDkB+m8Ap0q3gy51UVN4oK
KPTpS3NDEHq2AhurfrZlsoHa0eH2t1y2Iqb2DPbzTOzGgSNshD417WeFd6s63JZk
Mq7ZjCCm6TbZ68/5YuLSpSGPPBYOmlox0l2Dgsr6JUSiEDMgEiLFxaIpBj8iLruK
wHX86P3ns6YZIpx1c4sr7jQHILlAa46Izn0Yqk2YT+IzI91kMYBQuWYP+GCffvZn
j+mIN8KRGjL00ZYFNnZKBJ0DRjHdNy0wcA7QW6XA9pYf8oWMjGZoGJrkNTts0Zsn
lgZApbCkqV2CTSgklpMuw4qOInTe7cBacAALbN8JfpAw9H81B1P1MC7h5/wTct0h
oy0qlt9rs4i4UohnnQi7KOKmwm2omS6ZDlQxK+MCfTG37tOpQVm8326VQnS8EBWg
mzYkrWZF/vjqj2UuHzsIC58yucPcgPHn/KuJR9IkHaPf42kTGqxwhsv+m0w5kRp3
XSXl1O9wByUv36b062M6SpfM81RJznN1jmuIxhu7CIDfD3GuOoG4DjnuiDfAip0p
QCZVckZWJylUcc/1TDwv31Wt36ZqwwtdiQ3Riw4DZEa+beviRI3Wv1kolvfye4nL
fZ+OIf+SoZG14/TaxM/Y64X2EK09E4O/VnKFclRrDx4KrSyqpaQeJ9Vhgr9LaKmg
s0aHJd+Z2oHixTAW31MYsg73iULli4xaBNgF0MqSCwUaXLz531FDjPwTwh1FxyGs
WRIogtAgjDdQJa8IsqD6xZ3U3wQp6jmCRQAlFEP4xhTbsD1jqetxCK019X+mUsZ9
BBuPBO9owXtLmC4rNwPiRs4jGnqhGyVLd96FW0iHsXd8/beEe/0z9XeYcrl69/to
km+XwqG2ro5mnnnJLiMBdX/V7jhCPSMthdvBctNc3oNDAXnjaSLDqPB5sHZ6uhRA
74knKKzp5k6EmdrUucgxAp5qx+bmr0LBv6OaOdS2deHecb6GxlOtSqibKSWJIZX0
e38beAEY3qXAzp7kqeKDouN0hiq6dIMWya6nDS3HHrZmVzi+z1bIadG/zI12iYMa
FDwDbW+drYEj8Syj8qODVmr7DaZWf8RlG5Jcl54jFZTFDUVZBebLy33jdzr0CvJv
gRIQJkeTgQDmf6Q5ROpZpkBcM0LUgHUK5eRdVuni3JNcTbnM7Ep6AO5vJ/0hNM7y
RLTcHAFpc+ZgCTqC8aiakkzlVYV+2qPfslAHhK2WKQmxrs9he62Itx7mvhRWlkIJ
BQLQCYelHzmEk+7ZyWEeI4cGb9Uw+2448yslJwi/paiHdPXWlUOoomIXhhZJuslM
3s97BYj00TORdqStW7+JdpCy8NP0MVSycZ9PvJlKcp5oE6wCI85/0qVMtP6cu+mV
bYeL49CpXm6Bg28N80r7FNUKTSvPrZfjyst7nTnOH2etBp4EHNxDOaAeo2e06yjX
7yrN6rvz+dqllFaSDJcvLymUiepva1H7TO1esLWsz5RovCntfxjGM/2Np9HrKF5y
Xuq27JrZuyFscTXowaVzhwSlpoqBsK/h+f8tyKaInWlI4jv1CH1fYN5Ak38kA5w0
4z9Fk8cIZ3FGhiprKlPc8xoRMP7M8qxZDvJdnYAHL1JwoIAYwYF9S+9epFABRFmv
hCVk1zKo5R/t1+PNFJpFP+iIzUZzNdA/nbcibaZDzEdrgxbJTC2dgANG52Nbg69T
EBAPXgrC/sXUDunpebEOWjMwGFH1Q0uUaXQElnRCUX9Wq5/hfPdP/dAGHALOaSVm
4v0Rr/NvmOsSXqj/VUGQlxfzE3i9VzNNYh+7Yilc2oT3S8m+DfEjIr2xdZWBppwj
CO2ExLEXaRW6PBf4xFn33+Pl4Ksh2pnw90/cwHe+mSOM0S0WyrnBV5qKD8nPEHV/
ZrAn2M4wMD6DTqYcLaZH1qECNqGaJ3tmFEiW109574tytQ1bJhiocJXVb9O4dSMK
Fmg0bOOswccQJD3K6pIYdCuvp/DA6iYhAeEqP3mgMKo9YZGsEYprcxFuYLtWwhSo
tQRZfU5V02USAQhXOHEGORwYR2mDUgISinQqIBo/sh2QwQVEBNhnDOL0r/V2+7oV
LZC6bnYq5XcbteOJPcftVeGao/dNpATb4VesNBv1JzWPxbxWiHmojI7JTokOkKXO
kpId5qPXedWR8WpivTUdWuS08kgsxcu0mSh01A8AGopzPJFry/3fCNDoA0glEr0t
RWvGzs7JluN1fv+TY7ZcdKdqnksoRkBhSuzVVuO8P5fg5RjLkBysngIMDYgNYewv
MLjbo/TiXY2rSU7fSx2R1LZjFJYCWaj0AfTdp5GlcVyukkjihi/Pfwmrx5hl7PrG
QFNdCSfkWi1pUk32a0fCp8Xoxn0keqUH8PstZaD06FYTpZ43owg+NpQAkW5y5IlV
UEzkToMa8L34VmQUMdHj9cecBZ5Pg770xrMIdxu3qEyk52qP0JZUjUWPCCv34R55
wo0kBm37LoEOzz2Qrw8UiXpLYGv7zCRRb/4fvA2kGUcvjIQq+LCN+yJzscRP3v1L
y3YTwS2RrGUjKzhU5R81RrIFjCBn5aWbN3lp8+sPEqT4wyzAuhhPU1pfu7ytEKSm
UYsNQ69Gcn04vLjzicEyuZgsoA8odQlq7WD1b3Kguvq6MJmWBDSqePEzuNrQFDGh
I3b/kSu9am3mnGNvcJObfHCfEbMz8Vd9zifE2lxPprnMQTYXYQwt8AV98hrzc8y7
IMj9RDY2bHhIJhSm2pcvIpIKGJEGF996wAyC6NKh5yPVNa8KGd4alolCilwrcd9G
40LqILUmbg3XH+kk74Pd1TEStygr9ODMCRU4fp9G6m/ezvLKP0+A2uv04wFdPTc3
966dr+5LmRPU10CeD+EPOatn8/qPTrOGZj2OSZQhnmFv3+EpdBa62wKV7+MfBurd
1vd5Ws+vujnSLwv3WB8kXCq1uR0f0zOWGB2F54fFr56bENpXrpiO3dJD3bunergd
lTuSLcXlqD6IjzI5fn4O4mSj44BA0xwtHF7vBj4zB/fSaY3L1qRKTVYZse4Kw+fO
orb0jgr820WnEZ//23Z4r/OTKIhejH/sK9UL4x5BK66Ra107e9iB3w88/tudIQXg
FtzFhheWA4yL6sX92fTSY7B1TIh/PIF59iL5a8mD3fiJy0v2kWe3P2Pj0AGs8+eN
386KLsS25mbPrJY0GfJZ1lRDi9sdJXixHcRUHC2Ee4WRHXcTXol5epL+7LRSLt4Z
0zBvxaJ1U0YfKNrTzCZQXNjkbj1eMHQLCCH8Sd70QfKlNCoQKz12phpX8eS67/mQ
gLkEE5iOk8dqNnceNMRWorcfIqF1DB2i+P3WXpW9o+BKtVZceAaF7+X8jv9NM0wu
nBdeXiMjhYQdz4odlW37QrszzSs09jxWaDoyaqlqihkrhnyj85R/OpWLMHmLnzXL
65Tz/BgG8BMN13yASmzBUn+N0zC7VH2GlqWud61vISrThXnio1lFBTx59jxv0ecT
wPYDKi1oRBSinGVPVxpniPtaNm+piYEQdzQ/4dEvsgdo+9FxOSGcJYEbRyNQkAAO
kpNJdKuSZ/ewmIP6oOPrPY5l8PTTxWDuI+iUehs+zmJbxdS7qSiN89c35Kh3xfHL
e5zskD8/rfM3EFxW/ASH2Ja0Mj7LMuRT81k/1VaFAzOopo4myA4KhCh/71KwfSXl
o03ZWsdjlnDLydVi5FGgRuQ6jjzl+I7ziOYrY8/v7xKcAWD3e+VkY8W6XqjaO0a6
vaIo2KXorCdSriuJOLW3S+fJWObRMl+wmgNFGSmCpkVdw77Ns+zriSN9B7UREoDt
yotN64uvRSCFiE7PPmAScRkF3xKkgDX6gCx20ItIkVMO30ngL6T1iVUDY5ZwlxRb
UQJ4nDOF12UP8WTLDOAnBALM+lM8Z1x54jgkv848RpxuyHDSjF6zEIEnuLkVrcby
eLiNjp7Pb6anjak7ZjuNprtVqSRJ4j5r92bWzCj7ndY4T26YoYgNKvGw1MEBjkF5
RSBM35FhPW389lwQOdi1XXCxx+XISKnCQ1tmjXciyZP4ER5eCMDCXGoyq1kSjXiT
hrkxbhEjzcTzLKJbHGkMrzP9WJ1nVftuJJE5uz2e/XmN9VFI9EnK1OEFD7MnYlCd
5tJzk9d1BZPwjfDJSAMzR00GW8g/39rpbS1PbO9MeKxfTOntJBc8RtBuw652g7p5
lUWX2KtCo1urM62RUWY0s0Q9wLgaTVr1lTTSxcOi5/prtJcA9N442M/OWXe46OzV
TipUXaG+BZLGMfyxmYWJIT5+PdT98Ml5BE0hrNNMfawwtcINyfrMLS1HmQA1hzUm
iRp5eiZecTcAMR7PWKFFapKLs6wB0SBRphlI/ikhwTweahklFJiZ3KYtFv/23NH1
fem4NVbvTXpWFpek58AdJ9u7MH3th9yxi26tWdpsvPrhLH4c3N0h9mwS3mRbl9VO
z7rGSawS/MFdwtZcBD9Q8TpSyQ2OBEh442tvTUaHk3dJXAsLKFthDod4bBAFY9rn
I9VMqdkw0QKWMCGaaMxqJ6UrN9OxOaGpXE7bw89qtA4NTp2pA6oo3JvG01w2voBu
yQ1Zzzb1L9QpEAbMIZWyNHsq4V/VSiQB4SEmmmQaEbdCczE+sF5VUpuPgAvLreQe
EB8GGQ0q0l8hD6E8xgyR+jUOsH+1WwZNqE3+sMaDYR5RIdDs9f7cal0CBfIo+gtA
lUqEszG1JTHzLAaavbT11/bGhi15PX1Vp8m+m1ZTN8MzY8Ej5MIBLgzRkdHrCRVl
QiCiwOgP0yVoF0uQHAzPwm//s/P9IawJoV7FaeUPrx2tT3l5fajH/RenkfB339dL
TmcdzoW5/5WG/QxzsoRygtCuHJ84s3md1vErrZzXLSJFVczYMKw8xW2EsVArZCLP
sfOPo5W6hlAuAdgVfjvfCJrCqWfG9PFFtWq3srswdHXkfbZP0PbqyrPsjfSASYCj
gQTFxpNkEKei8oE14qmc8713aDbfmcOsQWYYcxoTsabjnA9fnJrp6cB/CmkRkJ3X
PLy8uk/SMACS8ODdU/k+V5sL+MNzbLKouQeijX2m2swn+KZWgcPbdYhupOgG0/kG
S1kjmYBGYAhrq7Eki0bbJYcrpolxIf3gmAn0F8LwBm7txfKMeYQPe+gJckRVZ+Hk
AzQLqkgk3PnAs8XqieJVx15ivEu/tZ2SLplny8F0kK9Ex9Zr1eNDjKNACXXGgkNO
LKYiz6dpCB0iJJvacw8/Qq7pAlLaa5+kUTwVzm7PiwbgfXHzA4sfGSVDEJxIKOYK
2+sq6tO5hxhZeycHDknxNHzgpOn2fz9VW21JBwUGOlZ8VinSAWB6N1eVUEQF2Huz
TDczpx6nw+ryOmRLtgbJ2nO8IQBX84X4lOQ6UQQrYvLzw6ftc+99G5+rVtlM6cSc
2z/SIy2lzrUlEhCmRiJjPA9TMXZF+3+OCS6JI/ApXH+fB4F/CqmYfIGNNP3AIQQF
2j4zbro4XzaBLmRksOoq1oy+J7crhB/KjfeK3IM3ioUmiNAkEDpq3F22CkQmMdaG
YEstcHcgdWof3iYNLf7vmxBg1MFHmTFPBZffWnbi74EYZWYJGH7r0F/Ib0VRFMNU
UIiHXXIxQVgr1UUcipidhAkpr5bJH3h60BRzJH1Z6rl4owKoXHQuS7LfC6z3XEtr
/o6YhfvxyVNGhHQyk8Iv0eAlQWouuxdTxdJETtVWFduC8YguBB6HmCFTWlMbM8iy
1PbdQT5QJR1nG5v08Swjc183iLNlKdWWA92YB6TQIuwhePLLwQgaVGRN/9bTZQad
wNA0NSDvyaTPmhOTaGNFV9vlbsDIunme1M9rpaniGuh3dh+wvUS5xXFEl3Ve2y/d
ZI+4EcT+vyzpwjqp+4WK2nezAjI48tfKq378QRdR6WHVUWK52ulR4yX9L1cuwSPo
t+aEBpvqZfU9HbGViE2vLx2akdSrBjsW1sPApaQMoFt/75qxJ4Qd67wpe5YoLqeM
yWZnEc4Gth2HvBanKFsDrmhYAOoUiZiGCxOqVeHIZ4/vrzuUOtXdcAOsfnjDfdFF
pmZrNP8+fS7JEzccp/LQZaIm1T3IzS2e4ErV4lmwcYbqg5zaLcqIYkeuIl1rjOlg
HJ11BuwPaw7YefG+DMlabqRPeGnLSWiDoRt3n+IVUrrIl7ojw9DyxDUc79VQDbeT
xxC/JJQ9mxUcqGoWWexm7QO7J7Ks2xQ35Uzz3c0uknKUMoQs/+m5tdpTM5FitfWm
1u19Rcrki+OKtKMZ2zCzF5aCBsX+xLNkcJJzsnHu9KFPOIEyKgVgPxLvfTkDD0TD
obU0EhNi2FuI9QKOm8QmMBmpbNJrvLBE2YPOG8vaxTN+XkiN98m6XMQH5UfAkRNr
lTVFJAQcNbxeQ8UlH4IhaWP3HvjsDnjOeONDiw33SON0qySvN/ck/CyGXcMv6o4k
3w/yyqgYY9Hme20xipRHmmdo1T2PkJre7VIqS1EQGNLeiD4I+p7V/tFAzssxeGLH
WSOLIKgx/zWV0HyS8ObncYn6X1GceL1EluX0uTWNY7HKpV+QyZaWNBfP+imPGXW0
02ljg1lC1n4RvAw1QDEsn/TtjhU+iyWt9ewFOOCAxmzXpWdeaVUZMH70PX2ASDnn
n4Idl2T/lcN6ZheHj1B9iwtV381/n5SZnCQOmaj005olLJA0B1cf2qd7LBDFKinH
fP/7mR0qjR/cwQRmRLHoM4x9pqK4Fm8C8XhmMEv9lV0FbmqIeScMp8g+Y4+4ZiHu
Qm8PWLlvmHaXa0tjsrhSeo7bx9SW69HuEX8Msggg63OVBXfcBT16CTP35xTMb2EK
9hSRHAXulwOSKlU/Dr7uiTqsza1oP1iKquyggwoQGxWSUuy0LjLomJAdEK8f1Vf7
5HOL9724P7soFs7NeYhtUpVt8NNRvEShak7TG0oK5GAsSBifjpD8iUqviKjevhYU
07oQrWdQHjN+hD9hIXKhcp03ApHXYK1TDUuY6sz3hEEVNN/K0JWqxeEuLvBX2kIy
qS7U8o+yDN4r3vUQCR+/sN/23OrgkE6GrtHq6FWAyekmcj9V0OFfB40EQMMVxIK8
u3iRNV+uk99wnEu1hzRrUGQ9qjg972dF441ZDDENs87OIHJ7zmFRbM8QD3Rtjjek
w6cYyAqS1+j9i0jYQA73XCmeBFm0xGMc2wiOpbHpkW0p7SwPr6XAcIweyO7W/Iqx
mPdaybz5Y4Dm+FLJqWNYPOAUxVstlLo/yusf2E7Mtp11ARMANsdtTIxhCFFPyC4n
uH0UAa/XCyXvpNRgIq3rA14BscjV7ywv1GQ0u4ElMcHNdMAaIcPNSQQaU9iMHJrO
5HIqhHNlSCPGDW7PnoRGDIEMmMuOYhChdz2qT0JptbvfKPQZXT9ZKcQsff3hWNJx
HKXsO072o88iOcYGoWRs1ntM+jMcAPRZTEHmSJzIcyMre4Sa18QkJwHYXMFZmxrr
jDCHwXRO6OZOGinmC2WgJBLIqehHGsrjy5TqT3dymge8NS2YA17O43SBQdMXnNUY
rAYelbw/axdrE9oDZfjxOiB6D/zP9tjz2Uenopn2JNnAKT7RAg88lwum6rlh1FXq
6+cNdblSEpPSxiKm5xaEaB8M1kE5iZAqtMKaAHW1UKPz6gPoLbTlyiAr8KB1S4Am
BN0vGsUfSepjGNb9jNFRCwEo2Z/ORhcnZxiC+HzMux5fqmFnRdOFSZd8lIMRMLww
ekKTaJPacevL3o2yjikaI91gGA7nr07QgzL9XrWey0q9G34yPOtdhNfqBd1aRDYF
lYAyx87osINmoVZcoX8+O88D9tgmC4Ovwn37HF4BfzozV6Y3SJU5Rvq9nkRXrjlb
AH+hMJAh+EEskTebvNghKx3jgYLeLOa4hnt9rqUKYGJrI8qzaIP8kbk209DrIvcq
LdMuezjEDWW5PXVS+Orb4xob59j5PUyKuVEFYcxmF/wTeKmAESt/MR/DHyeCbJyO
Fzp18TAtU3i3V8mspCrcIXYcSP8+dESCsF/qzKWqT6HV9ofw50VXzhfWgpkLcSrv
8Jg5f5vbO7C61SItcbT3fJ3cremW3yjRqmy9si2N1g3RAzvKK0Z9ac+5uwmWf7Wk
rzN5vurGtYRK3Ukiyi2vOT+KchYLutQHH+pQP4jkBrgYvp7mz+m0d/thew3pswtH
uNcIBGp2YYtXx+0kjZzTzzgm0wtuSsOM9mHTlDkSzeipoRxZ2TrU2qtvSrD641Dg
KcsLD0qCBmE7q/pDeBfTMo1SYVL0dfaWBHt5WvkQL71bz/5n//zvJgOlGzJBphzy
P+dlBqaQvRq8rKdrWtX0KZpiOSGJ0EXM+yTCKpyA7OZEb349hwzDfmPYiDzK3TqH
8v+7GYhwB+u0+Pc0qDizpWe2gXeHLa76x7/aJJe0rpbUWiF4TTliA1YrIhsx638Y
yA96LKgxxKED/fHTyMI+3Xxk+7sDYJ6HskbLQBuojEYTtZhiHOj7s8+am6wnUDtp
OHqlvUCKe1T3RXX3E6C2uTD9HdRekdv6BYcn0xFwO9xNNGUeIGh3op3ZnyfoX9KZ
KuN7X9KvT6Bi1PezmGzVZYL6/jyJxwN0WOFBzXakNT+grMPCNzK7wGBt8c5aFwsc
mWYnWyM9nVQRVrK1yzPMkIi7msWXpnIO9XwK5JS5ctNkK6WA9Mi5Ppg6Znm5PYPp
D+35b4g1Lxgvmr5bB1up/yHfMfUYPRSdldQjTnwrWtpFBzyH2DbOXF07pjDrP3OK
68wZzQ08XPUB/dE2EOAbtHNEnKSlnc45YNDrEg97i4ep72xUm2NM2iOKRrMu+LVw
sKBWRwMsNsr9m+50J8JiO1Tz6KFdQfFJJa/k6frTDXrnyrIr7/9XQgzbGJEHvg7d
doDVLBI+RvtMJc+nniAmq8F4klWtwIBDaMLvksbVpjQ3to1Ba5noGIh13uvOZRZa
iV2cY0DblwypZWJqslTw/UMj8D/5eylcJoUcbMMH6UgZNP4KzyZA8VLMAV7F+kHB
9EhJgJrRrr8nRnq6X2Dm4IXXzNFYdI2EttCwZF8XI7CHvFlkVtezsBC2Wfk5IoAQ
I5y2pU9rhQviAFJT7hJOFmo4kw/x+/SRuZmKrOh3/V9P4tw3Ka6f84wHc9c0Og/j
pTBVr3qlMj2pojJHJHuBtZ/VVOUWmkoJFeKQ9Y13w8fhLizX0SbBH9S/FSa4M/ld
vLiyW9YXTLHJAWspZJHok1gG65LfwU/g3jlc4P4yf+dCr5CrVtNtPKNnthTXM+pv
kijrWuGMvKk44vjpJzl+Hie/jVj1WubYwUEcdVaC5K6TFlYzt5VZPLOp8ahx3cFX
o7HPsYOE3J9S12YoVSZ/Ou1NzZJ2oj7j1Oqm74Gb6yyiqVQSYqoLcazydvKXbXlI
lLedtcMEqrSHXus7xNJ+7KVnMq1Qg8pT6gfYNWjgB9YephoEEwn/P4/txvL/0vvr
eqbuFV/riwsBqWcINP1x9rW3ZlmsHhZ0QVheygcTcj8EN/NrE8nYMmmW3Hnhuz3n
hzP6ypAfmTpObPUBxmA4PNoytJhDkeu2W0OnNLvTO4d7DYokcu+c4fO93+OlEGmN
NsNzn3KlDtbMPyrwSECiJBHhGY+txbvJipQ6WakiaJTZRq2gV3pFMtY8PwVw10yl
lWp38Bvjp3bCsPa1YWVxA8SaWTEPnLeI6qeQ412OuHz8R2eY9/mPTL0nWCkHBxV7
ZYwfVYOdpDSBEtUL8Zp6+bOAaYwhqPR7i4YVtDj/ejmA4kKP1TBqINW7IbhRBh1L
cq2JrHIPm0fx498xuknEAWHiJ4P2+62+DkzHIR5crlWRu76emA/Ag+lep7SgVYmq
+M4t1k902wz41EQlMk8wdjTX/pd/13H//1swdoNLCwZnmcBhV7aSNd/hp/23BcI1
DEGAONMuy2qRgtqR5LvsufbJ6XZTIekEmtr0qDUqTMl6wdiK/P4X9x8dtS7A1BX5
pAS0WwbZkJ4+jqL4nuBVckzU/0VnC2JAjszX7uMGFOm68g+De7u0N3s6snIv+6hA
jRPVUsroTDp4yXjzHOyJ5S0YtjOx8CyEPI4YgZ5ENj/n+xq2kftxJAu+yLkIMKKW
HBkDAL2tZ5VGzynSW07WT8N6BLYyK4dzPU9wFQB8cq6Uulej8dJPASKe8z3c2svr
HKaopVE79QXuFS4Us6zFWcJ1PE3TowjeJqC3EL6SDXk6C4s5eg1tE1NHUGPm9IDe
neMKbXK8gOfBXm6xGcp8HVYmAZDWBGaTaQXjMEiwjogUBASxVujyYySVrHDbEMwt
OgyqNqvtRS3pFEhu3LFyrEnpK6t7ouRysN1UjgYzMIQTK1wBhF8ZgP5WfP7mRygT
nql71jpJ0JI14bjZgXsfgHCzfWFw+fYlP1GUc5xf+onPuafcWMeIhDPujDA8keLc
g4TkFLvtvY7y8E/St3t8n8I8ohD4ZdnDw5nzZdvnX2xgiEeiG3rM9hYlLr1lxzeR
2bU9RjtTu1iMT0Kh1hpdLkBwU3BHgNaASgnK4W+5JpYDQ5m7WNZmSpBKHLG40n/b
ZhuQlrXLgt3vd8UFGsnjrodX2LISJuyhC2DKOITWoEecDIa7mxjU7rbiubgnx7MX
hkKKUxdDDxB4aFCeYffvm8/DGkr6v7FzcYrdEI/1pDi7jjjTZFRcznBewiR9ERgM
w5GQjUgFfHnwvdlhbiBVKZKGRZHDxtwr7K5RiWRXSq68PuJS7ECEN8KnDEIbzIz/
rVuQrLzfzUO6zDroTgRG4ZL9qOrRCHfTXH8BdDRS1TCBNdZ5g7ckMG2OOfb0SGdk
eldToJS196lIy58vZbGDshCeAmJZx0ntJ+v7M0QjdYBdDVGtu6tGRVNLGCDNx4NA
MHZcHVWBTPP7feJbcOyAy/H3yN2INT0JPWO4F6dC/SPikfAT2nVvUPOaAQ48/KqW
LnM+ovNUMgEGDsQv+hIRQ2dy4uh3XL0lMVSK7DuPwGFlYXhNoDrDy/3u/Oyr8TS5
l6ftu73LbdD+kjiEHQEIp5AElPhWXjad3Hr2iyUTt2+stZeCALyxSaiOfKYVZc/a
MmIiNg7r4MPbf1W/QOE8ogIjEF3zgSGLryWx+l8qK2ljyKjhBdUgE84/OF/RM9hm
73SGvPuRUMb8q57kkeCv/KB6/T9t97snuc1zAmPZfHM9FmgXaUAX2v/VFSsTAw87
JzsmNleb0AVCXR4/IGdmItbcM76bPCChV7pKq/4bX3jtXnkK3pbItBUbi0K/tx51
xIv9rHbsKNTYcXjbHurjflN7EsPDb+D8Yqi2rKWM3Xmq60RTXJZgIiIJmcifDqvm
4q5lc2nMOOqYbaUMJgWsfNFKm/CrQ8VbY9rdiNpIRGSWL8TEI2CA/nAdhWAV/2l5
p3LUs2BTXF/5fzz9+3oxRyHlmJJ6yD+V/AiSyRibXQlLgRqrGBIxOsXshiRKIkra
OAKwfGAXvkDopx4KFnUoY/j5J9VD1yDkSFhgNAFiJkn0SSfrYFMGNbP0JR80S6al
+xmGTz5DpsIgXU1gbsqLL6qOwBw2DAfPLmYqGQr8rowSYqogaZatGZ3uxebzqvgx
d885IyUA79j0vCqhzjNSUt8l45O4/azKRRCDIp89wIKfHWGIbeEssH+3X6nFOrgi
QgwdC3fH9F4R9o+iVBmlp+hkqxA5eQZmeAJxkXCHrOYPU8OZA48acOCTHW2E/7W7
JzG9Lt7W7V4hF+31jnDdhh3PSdYaw0xi62LZ7rTapslIuaMniJ/iIP6ztqOKJxbZ
zTms0PH5eCjwVZd2rtdzRO+jMbdD/4E0qXwfwcrCFvmd+4897+0aKt6/jo/FforA
Ojh9ZRd51U9c2QxAGLLdTovkSqL5Jwl6hR+Vflyy4kUYH3H9tTKzdJ4Tu60Vd2lG
iOb5oqoI8T5s7aYr+22m/07nHQhcrUXFGYrxqaGsnKfnGz6mMBblCtUxyE0ucalk
vOgv92EIxzhQDzVuUYgykr3rIoPHszfbDTaXvymh/doBg59duDp4xT0uBVdEyULL
v+TIbrTr++fjcqUZaByNTX44KoTOlrLQIv/A1Bqbp4F4kKZJ9KUuFZxf8xfcf7XP
kSnE8HY9W2WNCx71NdHS2Sv0PWxmTDnlfaiUdgWRy+9QbA3lNEs1vEp5uspha9ZV
3rs3ao+u2szLdT5F/qhOVP/tOLag7UYkeMwDkx89RyiWd0FcRQeZkXVVc8EJjbVr
PobuivSXOdNmZFJqmtyoIr2oP8wU/RVgaXoQ9ulckpVjL6tqJcEUtIXHC66zPSiu
qIalmgo+qjMQ0pNcaxsK8lJbLV5GbUFnTTvP83TO0KLTbpzCtOBLEngyZJTbPCz5
nPVS/kRIQClpcd9jZG2e5XYbBJ1SNQAS0+BGEFc3oC/o5bkm7teMOWvedgk1pnFB
IciWy8lMqMYkNnEtXkqlJq5yYSvnO2drn+6yxW319fDBSkkyg6aNfffPiWvCNelk
wVad0a8/1EWeDwc54OvHvuf55rlEOcr3/CVk++BD7eR7A3WzUgHYWCz1fuQEzrhy
JGuCkfR5ELXV8/9jl1g9Yg1I7bWzvn+PQtb6yBRgKKVN8vP4naanLmvJZAnVszJd
0Wv5Fdd4pEKhxcyAXwzBBNZUY2+gbnIj/1TF7Q+XHufkDMjOtL5B1hk2gC+5/Spa
fIw9bF1o5nrRdpyyYbaDWLKNRsGW0xWSkDD+3IR6rs0ZCZzK5IQ7FIKhpVfLn656
Jr0DzO/+/3/CLykZIyWqjVnhEZtIVMIz3VQjHCqKC+xLGsNZN9TEsPcrZ3+YZ6Q/
mUWXY20O7t4Vrz8QfIhAlPJaYW70q1yYFceW8QkZAbk8qCMfM1yW8175vFcgfoxq
6zrJMA8xR/bbORETI4NL3askznbKKSqzcPOq4TKtFp8umInLGZkt3TpD2JPrYOOD
Ih1d7DwJ9CninfV/8eIlDWrikJK/W13IkABEeFtM3VxaXlUxsL1RZD/tSb8O7RY4
E5UUyOX2ai+9cYQWckMIhcoW5YhH9ipnqGc+you6RBTnm6aI/zWLklbih9qNibt1
FunuYtsou49UriFkI5llJgJKa2UES1hSLTcfdKZicLcG6gIOGPywF3BEw6AUhreo
sk9Gt5ACV7ZhD5G9tG3pUrwcoqZIC1Jzmi3eZ9b/1sCaoNDx9PjbDzXAjgXuS7wT
R0fH78Oit9Q3wRAq7FWL/0DXoy0d06q7eRfMf0eyQVE5/KZ7nHVotv3M0Hed+zYu
1TBpx6P+wz8DXdBvVeanT1BcS+npX+4pfmCYKkr6qAwYWT/l3ZI4ACkJ68Kx/TCp
9OdGUSZ0RYfg7ygoYSCvc1exK7Z/h2wZQReT5r6KXxej/qHA1bYtL//Nw9pjwkwb
uO81YP3m31iEbiAeLn2gGm+75ihjI3Uj4lZHxnnMM0Ijp282dG8LyZEVurkqJxXD
51x4FrPEtacO5PkiQSkOn3PCtNLJpQW9Ycv+zzdH0JGCqb1+O2xYT5hu8YTPfzeb
KfrqcoX5OcdLj4Gpf8V5lORcaxHyLDnTZIF9kbbMSPrNE4g3WyPkbSgMkarTgkWL
LCxNgKQRTQ5CYMBiujsxwMPptNqQJ4KF5/USSe+u6VzVF4MM8CBQDiB8i8Gsn7dU
B6H75jxUBaNOMX+DwQpfgnb/IWbJnvU1wv6bFHN5u1Wye6RIbt83iAgL6vrCXbZz
qkHxBmPfCK/ARIQIeKpCNLixwzeBsblhQ6FK/YpA0HReoXV1H3qkSLHsOVwhevcF
+hWpwrr1g+fWUcQYILHRdXl73s72Lr8bfd/LVIntTd5vZDFokHSGLQEWQxhYy9Gg
TrE6RbKy7CUIi9aaeWkwv3svrmWewV8Dnh0+uEk/VbPkWkEdXB08Tp9rVEwF+JsT
kRcZJTyyn5D86wFCLkqnPTF5DZwvS3a83NbFRo7kBB2O7QuhbSQS/s3YqmF2nTYU
LnREDeSxezCI4P8aLOOy6xr+Q48VgTxIJmnbwO9d75c9lJAeRiSHm1Q6xLDzCTt6
pg6+5/lrnDj5N802LPWVRARlyT2d3PwQ9LEScY/rZMtGfyhP1go9ZP5b1N41OOi1
fEpRTaQU3M2nbDBYV8MdQstKB/G4o7ww4wdhGyZL6U4GGsCdRnGwe1b8HPvs3mAb
gEhPbwoUxxfmu1C2pN25gxfqjykaidpSwZRV11wqTezhFd6jA0zOphbIVrq02aSA
BfB6vBj70BIs1HVpDv+tr6XLN9BB3n0IJ9G3vqVlUvMuEWpRHmKwnZGOhhgI+bds
7xSSWlevwSVQzZSA8iupKx6htBngrOuXenG3z9trN0qdMENJU2SUJb9bOXbZV0Iz
70AlYmswXRv5dY5zYBkl1X4ZDH/zo0yGlZlWcVoeGpxE5S2cyITceVYXMVFHyXp8
AZSR9SP7xZKG/XYvvYvIeVrj1817+GlDCrjfvmq2TjZpKR5C+yFJY1xTYZnOuKT8
K0LgIjGqPmFrNjEDOK3Slph+5hty7L6gkQpN4KBgEzP3/0PvomD8lh89IJHlaFVI
F88sZohZP/xb3XgHALv8E1ZfdPCIELNCHXHq/QaWIZWeWEmRAMzrXl3YdE0PRnks
miPT9iQBUahWGHjfWkN6dWjnHp06kqZxopgbJBZaQuPDpUl1UX6PyqmP1YfaORGI
EwowDrTyK3OYtUDwssCcqwcCx0hLtgatcCqbetYyBCTD33krnsu5hhqZWbmrc/RJ
ocuW15DBCeATBf+7yCYIwgk+ZpWFpFYSUNajBprzaUdAdJWAb0y9goltpXR/pgCD
tcG3SoTZ24xETKGKmnZr8/VN5mG4vuM7e4veMwPYvWFzvdnFFHOXLyLMaY7oKmci
V1o1d1+Qet+bgKbNXxO5ewuXTYNtEzb3WO0OHVB3B1AzrvtvlGu1QXeOz7FH30TN
C+tcAUTxDn2EMx4//J2XVsK3YqxzRpVq7BTX0HSiYrnY8Ojdvxat/WMQjmEaeyvH
+5paUG/+d4qfYQEcgiH4D9rIFFmIDIfzHTx/SErj8mDG6g6vsqVs1Nyszq2ZJUBG
dOWqqGf2i39kSzgoL0pxhrZ06eJl0bMF7YfSVcsopIwkY3rgbHDF2rstYeQqn171
7Yk8xwj8Mo9mv6LSjeUGPpJ/93YKQyYB5o1J1TBFGaAgksIIjTzhisYECNyddhc2
GpKshzTSMeMEBGyzaWfvw1xtO+282Zsvdt+gAJEjvxp24OWl0mUNToySyxuyeKxm
k9Wl9xD3Dem0TepDv+HTAHRxs16Z1hcJPcuyYAZuIM049Dm5UxwlpMV1eEaaaSKS
jKEDOLXUOCUchsc+YsfhogPz/Mziwh6EXmTHXXkqVlyGCd8JXTuMzFL2nK6TqfTG
ZQOn+73+gqLRY2YIjByE+ZOko2t4JI3GR9m6NaFVcZCV2yjf1vBtMRPsSiX3+9l+
ztzK68OaMmra24M4o+BDeHIIUMZLzUtJpkMBdae+VlLRSUQ4XL4+PqDQibUBWYmW
ADkEoA/09eTVXOB6+XrKheibT5R4hl41eFu0KwAtvRkMFydIuOrmNbfhrvzHMV5p
T4pLKLpCwhbmPD+aqgefsZed7+smnBClo41ZY2YtGo1GK9BHln9oi+HUW4Y1Xwwh
vU7mYxnkELYHFMR79Kw6gxlOpl3oniXd0saSYrW5QeItXu4OM1HKcH4uoZthFw0j
WAGKSOVkCwdybPpRB3MwU5VLYih1E9Og7G6gfbzSDy+1bljCIPr+GR+aCC1GGvCr
3rCIqMbOmzMCsTJOdxIMENys0p+upG6zeHA8NKA4rsORFp9yec5raxjVZsT4sBBU
HIelXTGd2mBZ1cNx0fqUEml+2UCayemSRoRNqEd6mQa2I58M4d+ZgnJUtA/zHnqd
yROSgbY4U/KHj3WvNoYIiBtOJdXDdftXqTTsRvdsHNkME5ftmXE2Li/+stQs7PZl
pmsJUa+FlPH1Xbm5C6RlMnkHZu5rRTDbtYUnqC7UTpbdbHn8DtPWCdRMIQXi0Ixb
r9/wk1RN2ELgf4uJu0tQNym/2NzvYiwd7Y+CahfC1SFMYI6PN+ndGg1u2MgKMOic
y8FRjJ7BrqgNicd/JN+JNWvoq0qSNd2hItlg1ydzgk88bXauMab2HsAZWUlnA89l
SdZJzTgHqDBG+3L3m/lJ5oV4PhhhCKFQ8HEOg6pGkJl2vGzoa0t3se71b8Mxex4J
rcd/skbPfLIUPyDnQTAD72vK/YclwBuKanQfa5FuxhA3OoMgUmE1t2QaGzhYhPxb
5AtU6/DjD3Nvt/4harvh+tpJcOKtQocQgaZgL5NHeLUQsVj8itNYFURJDPbLr1Zk
ihFHyzV7q5IywmYJEcC8YBUjjRVm39IaafPER9d1EZdZ5G4YtaD7DhbHd94b18YO
HByKeyBaGsh2gGPy2gTF/30TlTb0MX3zBg/FQiEQAiFHH/Ul8NgQddVZoAarNlcW
n2+ysVYekn0/eunCTx8YSd8/8lx7tV5SFIxoGkRwNCKm3fulIre3OA5CY29sU/Hh
U1SS/ykyb7b9ySWdzd7VTlk2lb+ZVZQwmzSmleBzlPMnoqy3C09WAirklzn3dH3n
SGM85/nDnSs4pwzk/KMtyd3ljONdducyV7J8RkL2H42aBEXeHZ5sUCj7VSCmdk7M
9VMJvEq0x8JAZoFvLYpyrrWOYJ5jPEq4EHZY83MTpsADPJxiP9G9Uy9P+c+NCpxm
GkPDRr5bha7EZdYWIgxE+JoCMqGm4GQzCbYReb9olNz99kU7tw5sNeDsqBe+OgIS
6kSVACW1/ZPhlOFZRANY5e2CAynDaZ2sI1QfBMSginh41y+/gmluaK0S67IgYsiH
TpN6vMEQ4r6SGzLmrmkQ33IkW7slLXwonqY0IevFSN03323X8EiPGtICJ6w+QGM1
ftTsrvwPenbZCXJi3pVzIbhfDHBgP68KYm/L72BQ2WOXVnbCdMAU8OARfTI/vr6b
1YK7+5IkXyJTS9DJ4hHHwKEJRyq4jIYXVScBySewnz1C6DXco0OMbmm0pL9mb2fy
cRzvgHVSejDpA1NjVJsPZ8GOG6Cn/76FSoAjWsZBUvDUagPD5U0AslNFZLMuApdY
I4W+5H6BS6Bg/s0n5EhVlcaZuKpnLntMNqzOoO6XXOTgh5+0umdSkkqibaAXb4wE
xtGdx6cid7I+MC3QWHVI33elyZzoBbdu/r9GOxryoHDH38x8TWiMOYAHLnvlBY3/
JGTMQSUk0e2DXXEdV9NTcH3ChJ6tK/ecFd53UTUo6JGjhf1TrcYax3Z0GQfD15mq
LD7rRXvg9dh1HeeM1WYw3LHIhXCKpAxzjp6vt1pVZu9qbxqcGxivDxT6lW/r1Wsf
HfDDnwLJ7Fy5imWXAoZgt15zG76zkmB9070W8DMbs0dR3V+nFyWQICfOdSTXAk2F
OPhSr8Fqvrk6Ro4IAIeKiXe9yrd1eq1U4IJ324ax9lx3cO2n3+q/ZCx88SBzfAn/
sET9aXb8sZiBLLdBsfO1br7nITciLSaSQrMN3/CDuUjTRnUM+ieU6xkop/JbzAxX
/Y9vbnQOZoKqeZJCYsXq7/+I6bC1kJDizWCvbuczepAO5HabO9oUIM0ilp3OZ7tK
6Yi7RJmn8zJW/1pH7Il1PFSN+uBBO5gLQEYyYbez6NXWxTFfmY+IhhOJioZPe7q4
50X3aqTWLyilPB0Z1VKdVtqSHlDQiTiUOH7NjhspNCOHEeHC+0UZbiK0NnpN89sc
ZGnl6VM1llFmwQfB6c631zjrGqyP/s5Pxql6faSD9cgMFP0jGxTdGj2raI234rNX
zSQ5X1i/aGsqs9EFRZLSjuda3ajbGIC06Z58fiF0xr5yeIqnlYwkx2gZ9DQ64gE7
UpbV9pntHvhRozLsmOs4cw+LtZscRP93Kr8bdAfjDcRl5vPqTQlAaiCFcNjRA4i9
Xp5Vb5ULU11LZS00KM6ipBR57L3yKyDZcdpuiEq6E03XeStPv3WBPFxS7yuOxuxF
tIrf6GOrRIFESKgnETfTmuow/gsngoofbTSKa0BB8Y3pJgcX8OucpNaDEm1VXEzg
nd2qnrOxfRvzUizYaIQly3xydaG+xhH9/uOBG8/tekkp+/SlwvyVCSzD/Wek8AVX
lpbKpjJgC2765inChQCqcx0LNctQsqIYr4mKLiuV3pi7dDzGLYML6wEqNqElwGfX
yzSeZJx70CGp6DyemNhSnrnQkmn6fvwtdJa2htHvqPAZv4LARev6jrtM19/K7Pnj
wMYdAONz2qqBvXIl/hMuGOTz7qAZa/xAeE3JxUD1x5E1vbkuL9j6+GAN+Sm7yo7w
35SuGpr/uOgmXIgntftxiyXb+flOXkKMR9znX75bGva9JRfOdCIBWcWRyRHgbvv8
T4DpsqXEl21HeYsgAHdmFg0uPbHzn2/s9gH9PxNIi+oC+oRCbRIDRaVdyWhjGmKR
Y8brOpLJ84iJcHjer1uqovPBcsmmiITvLqCdPmIn4LABumQrn2oY4FAnuNnacwFu
pqD4v05cA2iiwKgHjvQeDXlVtjAVk9YPoJj2VWuB1LTeQ8Mih8xcmrhSCNpy+008
894nQ5qoB4fjI1tiwxuboU3HbEBXcyfS5jgHh0/xqGLHTYLxl+eZViOoZral5A9J
EeZ2m0ng3PLOw+9yM9v7s2aPjpJmJ0DLsHwsW2FbYuLKlvDqZ+wfqv+0YheRNMKq
FEaTYYLSgmaE9PReR9bphIv7bGq2u5wc1L60V7QM6YWccqc2hhvSBFeeyuAiE3t8
gMHMmOi84P5f4Ct/Gv1B1aAtfn7YIhcmEAzLqOv9RA4+CUCfczvHSBMmkX49i5Kd
+CkSTyrpoyRFALAHpAvcCN/c3KA4RSAz6IFWeZ/cQUudPol49gSgLG4ZOEwXfKZm
L4IfPGbDTdPPtYObQwHFq//+9Nhj2u1Ct/EzAPzWq/ifRwlxFFEL8na5obzAAvZ6
kyUrWSq+5VH/ar8YFc/387Nua06cF0+DEvE2eUVc3XHsExCTUn0E1A4wpLWPEZEz
CpU93o0Vi75XdScTT8gn5ulOALu8Bj+1bzemlJ/A9hZIeN+zoOI2cAKeEAlQsajY
aK88sjlctRJIzXAiAETMipmGs70d68QJe6bQnEMlWCVeuspVOwf+3Q0H9+c2HEZX
2iVjnQy+CSWMCEOfCxUM9YRUPR4JWJXB/Q4jZuCg+qHhxyuHa0I6HUzlASlKrmME
afOowHwyrpuQcrpjYZlqW6DCXLXHMalC1lvg/G3wzCvd62WiArcdEMUETOsSN9QQ
giB+LdZvhSDPw0w5uT38I/tiaPIoCqyTiK6sJsLXrnTGkVpprJpIdwQ18HbEvswe
0QrQqbMrKIs8RCxAsLOZ0zYXIGjAAy//YMF4j6sGRTie0ZxQS58X+9GD6Gh8yu5Q
/sGH5CUA43L8uVni78VojMqjJQGePBFewbMzFRTUl3hbBOazjIVgVFtXYOV7dpSM
Gm4wabxyIaC1DTiR6RjozBDmsYRf0f5egeBbNPERT1lASKD6S4SWSugWjCYx/Jhr
3d0pVTx0MeCs7c362xNNL38DFMZUQ55h5gwHpT+kIjfRrX7aXjTqWee64EZf5bTS
nVttm65c8qtdrFyZrCX8A2tgMJ3SBSxDa0EdACwqf16OWurSMyd5V41dDExdOJif
EqarUuh5ZTP7EPtFDXyLX0IziXfiH3jIYhceSFGjjn5o6nMAJjaLVSaQ3HPJ2uQi
R/e24Q3P/jfc3Av7jK8lj3HGOWnmejHMdMObmUq+z8wmKnfwHJwlnkZivV44Jntw
ZaumoKJLNFGkdFWSGnpKvfUgGDDQYxFLvJqdviBIaOzveRDOy2ihXYcuBS/PkKTN
71Kee2MXZMCkivkDmSucEiqr4/rexHzcXfnoasxFMvx5isuveP1tjUCXBS/gBWmM
aMP7TBdedL0NaZssJOUcS6k/6cxdzjSGuLE2YmFyIwQFXPhPjkTXsNQEmVM2xxAv
1tAURwrcTnsKBexgg8bs/Ry8jE7PtfozYKdx7k9W2Wwh5EUCws+Km0C9eeN2d9lW
mxYBi3R+6Q9domNyn5VvGvfh9V0BZ/F97I0lGMb94/3sVEHo9+luvfSTNdsC60xZ
lHaYLKe5JRd5tw+mb4//Ma9RK/rtQ8uuhWDT0c5blnvKCnA8nLYlNwhbExIxSJHu
rfoi+P9iK3DDDYuqnhLPCREcCaQdfTVNi0V1OJejRcRyuc6l/HZ95bLd+qJm5mF+
f6sMWe4K/59MykH9Cum/htd9kiE14gHv7UOEkY4M11weYUjNjSYuFrSvwM3DMh0C
auqleMuDnyeInbCiuoBR4YMGwLqxSChpGJTMnTbxDZRVcd4zd+x+vLvAw07kZRW1
++9WA9abvDX+HYfU/NI5F450Oc1Ay5d3dxjan9r795OPdVUlCyY8u4zYxyG4yNy8
xontm683MwXpRnyS5p7dTKi5Z1oLAFtU5e1r37PIeswRtJbmOaDEAhkgYZ2Ba5Sy
/gyOH5Fffm02Xrs2Lr3rhsQIt0uHC2W0O3kgJQNR6oi5xaToDow5s1CX5IcjCwaW
xEGFFYxKJd6KVBlaSwexxCmsCWhM4VLxccgyFmWIoJ+NtWXwTTrQKigzT1rodAuA
NuoAyIaLb/WCRKrA4f/86knfhAGOngwFEqofJbeVvRKPCRDXKYduMiotdlI8wqKo
uh/5wld42+tSMZBHs++8+FTT9h1xqaZsVpzr6Nj33/zYvnvvv9p543OEeQGpeGpO
qcQwehodZAZ/+WHkbzU3IcSNFW993T8FXlQcG3ElllbhXsyPeYtqIOnDVNUXjZrz
nVWcgnwgtOeKPbKapKeK4Pm2tXWzViooFl0Cqa3X6xbLkO1OLcFCTnPq16OiQkP0
R5iIiecP1gk1lLIpOAd1p02x+hrZPfHHwN6wXUe3nhva/l1207bktJ6kNTbhXwVa
qwLTwsHX/OFcL7Yr7Utv5edy3hJ5oDq6M1yGUHreUIMdkUYC9cOXTxg3KIDQgajc
+Wug6P4he/5SJQi/zOLWRdLgM5+acn45RfwHUhGqE1Dv3eKFLe19mjdPIuy7CjDC
1M3K6YXCUpjMC2nG9zDVZqT5z3HTdj93e7IFNyZXCeZTgf0apMAQ+Jkmuv+T8j8Q
FeLjDKoFQeg7rqx9oKoF0W1ahlagVaEACfRfibnXR+9q0yZ1QWlSfwKqcOWxHNLx
sgEJQpO0CJVRGaDEoFTFoX41Al4+X4bsQfHLxIw5KDN+f73bYFDwfSBFPJ0qfErV
Kef0cw8Y9wLlmGiZlQX5+q9HWeyPqRhGVmZVmLaoAVXUYPaEzMgaT9DxXX3vRFFk
wB+7Cg42lzeC3HiLoy9j7WxbiASYmvKK8ScGR5j8J1ahJfhJJheR+yVRy+YzkLBh
ihR/dbw+yW6qg+cWsFCSCMCDo7Nvi+GRpy5Ubi4uyHyVD7Wnh0aT58W+jASbJE0P
FGpmv600sqDcrFBF9tt4dPz2aOpQbqBNOvYnWzE+0Trxd33k4GpQ2SDkZXvTiw7C
4HJrDqMXtKgiHLTcp2JeKXcTfpKXyW9934/ZV6xtX2ybxWabCbBPdmmrFNXh7E07
rdfLmoTFPOb38rUdeYNWQj8WMj830WYu9VhsLlAHNbnlroyNBpLbJZPCSm4wDu2a
pVm8WmuZBMFNQ55/tsWEiV7Jl4aa8UdzgBWcV9ikGZGApK5ue2VIUxC5UO5F6irX
ftkQm614QuVERTIXCoZiL84q3xI4g0MEkgmW711T4YjeDCrSFs9Fews6ny+061JE
yR68Wh2l8gwRrZp/wfHX918qHl9iHVUZuD06J7VCvj9lG7p9OsylhHY3KFwU2whq
Vu7/F1TNUvn2mQB4aFqY3yV7pGUfgcEskeZRtB7s+kpjX3xCGNWq7A56tdPGpgTd
u9/KWMHWWDRD36rfcEGwLtx5Vi9o2LPGo0LHTyQpE+MH820avV8+8fJTrxoC67Xs
bv9VZKUPI47TdCeLUG5jyOyBBLMkl5bEPRXZp26lKkE8pxRtvJ60/I+BK4X66INL
DqJCCjtd9lMTHco2umzyIowkGe2lSzdqXsomWttgcCx6zpx7HQlh5duv0LSiiNjo
K/N22aY8Er7LCbVefx5+cIir34JXvsJxP70o5Xaj9J4z6nzXidvJ9k3uZWwnim5o
RqlpUhkApOTARQ85ccivDnxEG8kE/8PgXGQMfU5RtNGCxWRBpYzJm9q0NgwLa2P6
r9wmd5mPkJG3VShXVA2mP3XQnWdAbWgTnRfCmBJO91fAQL9GEKkrpMQlfVkLeRk3
UdcrSV7jLLh81YCTMNsLe44drB6UN267qzy5J7+jJlRCim8jzJ/QKjoN61ajxeXy
cHYasDRfOITigvpDCA3s6P5R6DSl972mmjrG8dtub8dHA/F/+oVwXQDJLVhA+1AZ
FzlCqkIN4QuqEmxQhL9RLK5L8dGaMOILgs43iMfbmzIB8KTl3JTSwSx9OBuGya0r
rGYhFUe6SSEKBokuPRuVoIybLg3kbEtK5auLrlsHHuATMm232LgdSXoLVK69rlpk
WxP11YlF2PdXWRDZyluxLssrlDDeCbm7lJV75mGh7MtQ4LZzLpbndi+by/Gsh88b
EhnC8vohXSkz/IG1qg0wpl5DYPpKI/tK0Y/Y33mvzExxz14m/0M2T9/b/+Msel4i
tK9a3DZ2KpWBuptClPpq7HGhDeNNpOHkh6oiSGDhApboHRX1tgKeshD3vxdESa7P
x99PjBjHSC4Asv60Fto9FohKjvSks7Rpps8N1LKbCOAp9uTjwEqP/qpfVTIqgZoF
/ogkCckxD6/ILuY1XcruuZGHxTdW0N71R7rZLzpJkPoQpNkSiXb61VcWISuTr76C
vmcSwKb1u2oCgtKRGXZ2lJ2Ifs2TinNOK1qln1BdssuUm1kjK7rrfUwaZgwqlgQn
oL2I0oM7FUPRH6QwJ2z4EvJNIMRZj+58cQX0X38ys6F1V39LLgoxXjAErfezoFP9
FjOeD/PMV26N+c2nkiOBcqJeke1j+TZ4joIY2XfXMXl3XA8GeKOPlD1YDXpIB3lU
Qs5ck08EROIgK63hEiUIQYuTM44POP0jPBOU4T6q4ITx494may/4d7rJo68TDhO7
PwY9GbE6ctHZGFzsaBmMdoVmmjzDdqSkdi5UgtwLNY1NUyv4vYOyhQ8EY8bq+zPh
z+C9CY8OxvFXsdEKYuPTCBIC1KEWWGsQlY5nPVFPhC1R+MpifZtD8PW6obNRa5Zg
OLEsIjHxLUs0ZxRoTmbhvyfdeZZ6elBjTKWkvk7q0elMyfygcO5PLYtlQxzZhOH+
hMcRArVJTMhMMtCFYaznU2TrCU4lBt1tCGwuWppzO59qisSTBo+jGMLI2ndNF3hJ
teNXOyy9RPF7PogsHTPRNx3AdRc6AuaWytC8nApHsd5fk4+EDwsZ7xjBZVhgOmj1
XC4E2fpGTX02hlBhBQnmQTuG5uHVNoYZXvZU4ym5/TfYpa4s8YplxIdipMjC0OtX
YAk/dk+nFEZMcm5+yv9x/qaa4HkHpgVTpZ3BOcvE4VOM7TZ/m/8Ym070XVmkELWc
ndtCFGesajHUCtYlEz/B534KTdEpLKZEv5AbZOJ2z03ws3MBlENAx21suL+RgV8h
cKMEhAG6fxGGKlKuIKjYNKmgnH6rCT9KI40sd0dXLgelVIIY/2K6bW9WvFOC+Iro
zAym0sgtcN26KdrEqe7/yduguMHE3FPewmrl6DrUfTtc2ISknBtFb3It8QAVTOmN
Orvsb103D9qW+uOrny7vZU8B/2ZawHsCL9uEW5yy56JPHZHAmAado8adp7UxVUIa
BRywO0QTAcRXY0Z1lIC307MWdCzEBImmqBONetKevvQIh9J8lZfvY6JWi2UjNdhV
Lj4YHosVL0UYq2dG/Ue6jcSotXTJ/JZ7+bdfl3q2Vt/yL7lCVm6Y4USKhqEDlt+v
BsnqW36WWnt+bqzCHxjTRbnkU0xS+UCktmwsar3NCwCwXqW6+SvYYIcA18KLTrO2
537lg+XAa6XTSLS0K3SRdjaeV4AndCRZCHpNbwIi8zi7Kbr3T9Hp92nsuSE0Caw2
xEdUhMX8X+jdWAxBjp/sQdX1bzFvmS7zulVECHjGANU9nL1RaroEjQeY68ta4TNz
5L4v9tCUuMfpZJ7ozT+/asRH6yBeQfZCBJJNgMf3LaETuieRMfiNZ8Q76TxzG8i7
PlG09YrWOh2fYNe0SsCRlKdzzoJef93SPjgdUYQ55eRZ54kzdE7wD3HQFneiEeSu
NdzQSMtshJIhJowyEfPhiQKPhakHHlXE2VliW495vnsGuf29+HWGtZ1vCnvfLcxX
sLAb1u7eJZFfQquj7FdItODVhknuKaqCFPHOBO7K1MfIS3TDToJgN0CCVOMw+Ep/
GCDx+PXlBYtpoyzQgszvoba0U1iyRihLJRAP1H0B3dT8E7eYA53D/F6huGDgllBt
Wua1upcASI2hjQuf0SnLjEWs4ZKGTk6EGzG2VbGzT785WHcw7NFT+E5d9iZy/0Kx
rga4z/hDWnjxErvQJH9ykz/GAw8O6i0fXMtE9UwJvG4FwqCet6exCsa0tBESkCPv
dRvfei7Z0abtItpW4cnh7aoh57LXyB1U6d5yKuSPz29+zIrkIRsVqyXcPiF9z2sT
IyQfT/K+fJWS8Pl7UYbsQWwr3zoQ/SlXp7OZyvYNBVfw5mVnbJfi1deDKddFuAhQ
IF/E2e+kANjg66exTINrJNl/rJjhPEGt1vloLP34O0dTZ+ctOmd8XIV4e3mudj4p
zqVahua5jkY4D41tGi4/Au3hQrca33tsYiSgapfUgfalu1J8S7ovtUTbLrs0Wno6
/T3FzLBFbdwxosgJt6+NHRs2LqVCE8Tgiqf3JLUVpoYjr+kZTfMdo75YIB+DRb5z
2lZ8GcVRMmVmwspzT8z8Qx0LItX6a42LwXROFUBG1r2V9+9duLvoPwVuFIM/SPiM
Zb58w/AEWJvevl+fe1kvB/YoV/RG5TLm2JuLNyBFrrYf9mwvSZ7u1MqQRVI5gQDC
UC2wc7GMw78H38KqaQdj5jSbwrV/gUJtjboLVMdddHoVzziajtoNbBrIvBWwfhT0
sItZPHmAg+ms9HEFE3J4LzrPumWKJVCcXvvzgPuAsx6TQBboWbMPDCFZeh1AAmro
MlVgWiT9kWhWBrqhJ6uKmvEE57bNZ73YE4ypAzz+VyeJaMhpNRljUVpUNaqwflQ+
OYxdjyhwFecf+Ul69Va7gVZ+419JD0TB8GPQi2x+RJ8HuJYTz20Se6WpMCCG1XvD
vlL5s/TuBPvwDDCG0ia5UPHhPhYZ+0UqA+R3qLQxyf2lXcSRlKb2slnMr/tkYMbS
bSi8bYvkc/iBFN8mxtdlWOgOx78+tbUue4c31epe3PZbyq7GmAC6hHA+n7+cVPwd
eaQ9nWtUbRC1Iup1HTvJEp4m9+WdA9mvHuj9W7rYhjrUuQs8M7NCaNhKlQhWH10J
qV1Qbzs9TjMixx6BaNOLGSLjER/t6YxuMRnEwx2L1pRWbdePDMHGlbRyUILuWjT6
uBYndxaO2kaw/0jmvxUmi2yvjHQoxWt9TVvPFX36jhMocyU7wW8WEbnszyjdl/I1
Gqv6yJV8hrPoeZCikzrmh5s2znwI2xDIRHN9OiUzoyR/e8wP1uc6wQsFigXHfxQ1
4u5mabs0G/5BHb91mBHjtdkiU35tajndOKJ92P7X8cKfYk44PRbLEdS1iW7ycU09
LHTXrnmG8MahdEZIkdLH/u5b8lGbstJCB4zJLvQ9TyNlBPHzdxJ+vm5AEUhKiCV1
VFD8jxWDZv1/XVGT5d4zrZjbQ4H7e+j5NvLsKWSsAA0dnsJLE8nxSHW8xWKdIOhs
xpW5k5XXapy7av4g7CRRo38toQn4yVClJXkvSwcyaO2Uqcxe+3TcWIzbpP4JmdWk
H2Fnxqh1yilJXxDqqDcSAiVrCsH4GNEH2IWTNd9zyq1dkwPDeILulV9444Zz/O2m
rqm/C1ms6BwTBNhgLWeQ6APXcySIGyQC2rfvwcDGqif8p4KIE+5tr69go6zqt04b
pBvB+SUQHi5c6HydHe7mTFIMnkX/Dhv5COUUjtksUWX04ZTzGxvtrXkDuwhE4bGv
xmfQIcG+HhYI+FLEBgQZgHivlURQyO7k083855XqSPnEffhStEvYGYaOOwcEiGXm
yiBapGE4cDPPlDx7C4gI/MSB0rlP4pSYLhzwJICvWm8830RjL1JoM/vKaiRkLFYC
oPpi5EoN3sPqetIuY4sa3cOSslfI1mCkBEMCRGpwMxWI4Am2cwRSebCs6w2I9nvn
FBMpFrPmOUVZAeB/c+oIT3p11yrdRnXHOpksU2HNfpu5himeB6a4GfyW9i5c/Wdx
j1WiNDVfXBgwiWa1vETXxN8pKS1jOvttiVo+S+t9WHp4utL1jkRtDOvN34fsyHLB
eU6krd4u8SXuVQsc3UM+0xswHY524yHshMZnq5Q31Adi9n3LuzTaVEuNLlG0RVyq
y4Pyxti4vImCMmaeg+eKlUOfmM9Pe1pMfP8bMFLMAgykpGnYxv8yD2oOpfdifsp2
m8NJrSJkMeF/cMQjqD/arlPFp2YfIkfW3E9K1z7NfZecTRZlj9sTfYra9NCYQMVw
j5u3iYodI3reDAUEXCsBQNE26k5OckZ6Y+kn/wYif1uBq3mK6lryOyyWXJ/AjWf8
j8TbK3plZ56npOAKtzWlKXRPQxmZLxR8RFpxr3i7lNR/1LTrJOZYOkgdsoSUiJQt
MdiNL95igBiFWrGSyZKe3pXJog6/jxe+gerDSUG+xCxE/Tkx386zeAh0ecU/hUZG
IrLRqKWHb2ouk/ZNLVYZ4Nzgql/MqCp0gZAbSgoKaNS3F2IU+HrEpAcSa1h7UjNU
99U/ThQiZrhBLB6kbm4mqFBco9ulbtEnibIqmVZ9Mz+rEgbvat+6YfMwUiFqxW/3
kOaY0LdPP837lZq5KlBjUda9VBJq8F4oNpCUrU8a5X+5sPyXTyMQmTRHyqrIFolb
vmSkfVBL7uZWMIyuktgkPcVfpXnBOVjeMkO5bRFdXgyR/WF5t8y6yyWlzM5opg7C
F63R5ZlYdkkBJBdwr1xqI2rNWMUYkH/2QCNaD3GZNVW/6/fe16ehtX9LbU8h6xWb
aaLVy+bqkUVe7FeB0uSJdphqfgxwnXlKXdWXuoL8JKHBqU6yXv7dWM7W/DYUdEQp
9v8tE6YisUxO6CS6cAvhHSwaO9o2S9ZpAFCwpGIyjtsSiQ/EplYKw4KfkRPOyPDM
B/+OMM3kCEEoOpsO5y8aA0wMmQSLfF9d5Ag4fBt1qn7+NbwNV3c61dlS6awRBAGA
zkPcFTC23RGHxQnSqnEwaSIX3kImNNwJIzMOaHn7zSg/bTstsN3v1Qt2w9fKFH8D
GHqnui1A4T4khxx3HTO6zSMfZQfTEDkT+l/gx46hlaVESG65KVPJwlZC6ibkOCBM
fblzE/L+YfG/AzCSSkf45fWJ+UTTFXqctzKrR9/Itpylrl0bWAj/CQdQn9KiNOb6
HISZaSPc45tLe5kg+JiE8vmEjmAXiKhtpo9n1gaHXXYzm67+xuCCBc5doCqk7uyR
Kt+EhcCmVGNgoyGVymTKid90oxS6FZ7L34fRicWqV4fNkV1ZgRmh0NhH/fZbuUBb
NlHUmaV8K9ibQVL3DSnyLi8dqeyX1ANibw5+jJ9/0iveHIH/aWIbjtP+dgMyAeSD
U76e9i5XylmWO3GAjAcbr1VIZ7P8qNHgnuA87evF36zTGvm7TBw2SwtRXgjQocWr
bEzgUJFb+5uVPRIaUNaLMfSdXdmYQw0D80K1/ZL9vjBVXxJE5jDO2kZ+R5HFu01U
W7ASHOi1evBinT8uVucuBYhpbIAvZwUAsmYzCjeDhb4Ts00AlFRvlz8YRpjuAS0H
/dMe89rsYHg1M01akU2/NrngwMSNMDnSGHgW/fZvbKoxvF+657A8/NbbPFGo5LJL
sA6/DM+13HcVBGtPfpPHjoq0tn6kowZd1QhMsQgBm/33JLxG/poBKQ2fyedd2vQz
24jFy6E2h4aETMbUEdjg9AdF4XYfQYeH8MuvSMHAeDuMOxCqwQ8R4WpZPrCspo+Z
A14srwRcJLawIXYe1Lw9W16vidv/bzmukkZyo8yxpECiDt1k/akgsCdYHUPOEXsH
lDbkdrazuXpno+UOLik1HNez4MSSf+SDcLrjZdQkyOn24rdzMA9jZRty6xDLjGo1
/HmjkS6yh421WpiV/iu6quJIgKTPgj0Ex789CkmZ3dx6hfIbXk1/eiAZMseJGl/E
2/61cAK/MGcf34AVo5sklWw/B4k+WudPkHxUW6QBXm7xxOLniDkgYg7Nkuzi/0rs
QduKK5MVpy0WpwglGWAP8HplogsYfGlC6FBdt+yeI33w/qkSS7o/2JgjTps6rJHG
5S79dgi3RmvUslJVFh7mN7Xsxx5B4TB8YFGNlDaZYTPwoc/gZn6BDE4YmlRIQxsd
uJeGOIP19qlU71ITy6JfO6lXRBuREjwkQsRgtAyDIuOrZU8qSKSXXvWb3Safuydb
toy+ViweN85d6HgpqxjeIC9DpDKVK00XKbjaSJ2dA6YncbaW3JDCDULozSl6N6DG
PRSx0SPyd6YsBp0seUNuDCwtmk4uyLDBCndnEYopcbdVjBPIAnEk7SxiSPuovCW/
0nXX5quZ9Nc8emezqyUKRxAwRsyshqO77yjOd5raKDoQxsMIE0wgD8XIxTMz7+Tr
1cqlQR7ddoFPW6SCez61TtFt0hTFnd1uXsO7RYdHYYpVspRoq1qAXicB3t2xW30j
H8xBQKnSZblaVES5ZJKEmGfNrbVx3g0YPkWthrfOoBLxJJh1iYhV57FdoMvTS3Pw
SS5OY+k5QFbSD5sb9IVZhYlZScaCgsXbwBSw1FQRyFaa05V3IUF5JJRfERkUdAPx
gSS73f5SNr6M9K7Me0bZt2v0Zt6vY0Lue4hL9uuy06NKm2RKCtHl97GhUO9lE6Yy
ed1Oiqgb4GVbN9Fpf8SY6YNlxPN2q2+s02vpT31QwqkWFNpaUpK6IYbAEB/SfPaX
j5DsEtAEs8+0AtXNj+OEQPjK13SETYuSmO7JZsaWmF2EAoBZF2opfhYkJDpmpSOP
K7Roq5iRldoynHTCHZ17swK4MnoTJ2DYnGH/5GebTlHdnkTsxnXAMQzWyF65pFag
DJ0JZo2uyK0XDwIglZu7Mi6yZlNAHtyiPvvkLa5aQi9vBu70HLBRN9p0XmUKCTG8
nGaDKE3cn6G1AzpM0PU7pQ+nD6z3QzIY09W4OZCn3S5rmyR3RpRA4SMYTZYjuJ0e
Yt/GxtOz0sG5XNetKXW4TRDOgo1EQ4IMHg4ehlG0tp9GwQXXg174ZFx7oDnVJbj5
GDf957k9aV8KKX3X9NLxBc6J8YHIHPebJRCcsgiotAwkQwKIEN5FsxyZzhD/L9EJ
dugeF6DahXXHbpYumDhEUyYhZw7WaOzU5taAV/Ndtz3MBeYe7KygEEkwH9Pv4Cgz
dTy/CpUV5lZLUb2OzeOmtaTCPHZuvWOkmqjdAou5KCrFfTCJWTnpdhl8fboFOSRp
X/jBfbMgU0mtumazP811bOFit/msLgAHFqv+TXMsT64GvhOSsOGRMRkigoQNPAKp
E+hkjTILAqTzGzqoKFE9Qmq7tPiXPL1YxnauKjgmgsKIoch63ZpdVWAjtFh96B9M
DcaHe6uOZlgP1pYRXPaH3NawaFynpD6W6U/mvxbRt+CucBjHTlzDv891fK25teNj
l8GG3Sxtkv1knkDPlbRJ9UkbJLdJk1eWtxBS0uL1LTFNfT59htGeKqQCCYmFLcuy
3tf9Dwfw3TBbnBwZY6C21uF9ZfiT7Vimd6TX1QHxEX69pdMixvfjr1LGm0+35hoa
fDKeejITZJM7XHMSeVz6qDLgnyV+EQ9k8yQAaE9rmWxZ92ihvsgCxUdMEIWjS7r9
wEqCAQsUzTeItyWKDSk0kv4EzpldT5QGtvMIOXbVdyBdOYYUCsDf3WLbETDD6K3w
+ZkC/syZL++DRkm1giUNXfel8FK9d++92tS8YtI8TA4n1mB0vUDjxvzOZPtiC3Wd
bZwAzY+jdrF/6RNPLgj6VdLHm6gmk7BLIXcMISYKkbqJGkXHDiqb2xOW+kGUm72i
rygedmaSi7I1GCcDLWd2tj0g8dyeGjqdIkshhX9TFB/swWsoU91jLx5kcZdwNDcJ
88vea6gqFLD1AY/Mdn3WdIAUkzx2/Uzsa+obgdOAq8T4rzsfoIJY+rYDdFyfSz3Q
QMK+ZVU0DbAij9mnn9Vwm394xbUZGQT9Zk95wPV27vDcH3Ri0sH1mjY6XplxbFEz
Pwo6kkpcG0Z8Z6JhLuJ4gRFrWNI900+Ul8lYjlXKzqHUPNln13uzjeS8oZr43RlV
/dPSdNJpavAxFaYU4mXQlQ1Pa/t1QVqNKVsRqgAqi2LX/gwPOYDIH0inbAU5L2FL
YjLQp9mExfQYa21fjBZdmTb9MuWwlegZmObnnq6o8nXPkmunvVki9rbbHt2s9aml
7/rEpQVSU/mjlEHqwab7+71NALGxUiJFfIIg/M87Xe6zl7OZJoRZb5Rlot3ZPBKF
6P2s/j5xcbzJabcnQnyS6YuBerd5LvPcF0i2qFM09HwNvxzpGAxHA8IgbkeT0Yc5
QtmPlP7yhoQiEn+pHfd3hrEmwdGp398QyEPK9c0fcErmD6Iuro0YhuGVUA+0OZDD
tB8W3OfApf6W2Vn2jBmztQ77Zpr3wvDa8pw1/663/DWnH7rN+Koq6A/Izb/JzP4w
czJunhy1rm3oP4rfOoNOhZxgiJX7xJt5LuEbhOV4an436D257/CybH7QMHzDjlzH
9tQHU/dzqWJKfOtjm+bMK/ovEeQxR9OB1KDD3zqE+Jhwsq31w7DEdHfiUkUKkb6g
e+h+bNE1qTcSkvaVO4ys131FHoZmIohT9Fd0N3PLRPFGEcS8fy3EyK7w2MnN0Z9+
lApuHLX1rHbdYqB5KIyb/ryqrU4z2E4CD5hcyGVd/CC6X9jI+APhUNuGGMlEVwkz
AbrtKIsDySs5wZYdJ5L24e5aRQKY3PwiHS99JS3mJnttD8g033CC9fP9AodYfpLS
ODVQTGDhExNB8OeLe/o+fwr/MlJpD3ClZPPA0dDTeGdl4680r6jAkOkSwyBl0MML
gxLmrnx8uwVA9+EbGx2KTHQ+jnTr9Qt+F30JV7sP8utbTk/C8auseamfN5ivLMqi
8E0PuatPXPJp0ODGWj20BaLcGBoYtqR139lYkDfmei2g55ehRDhpISSqcinHlmrO
Zz30VewOjYIclwIf+1O93tyL8MpMRkTvNxkT8PRYBtjJh+aIxWKfowKUqoPt8CEe
n/iaWMUgXRSBxMv4KNRe+7Lia1zoc6Quh5G9b1e4N8NWMWupM/fQT3wrKo5tTiGS
lN0IE9TR2oPTSCok4UOwCHmscqtKREJc4XUUjwoAIZfxqXRNvXy1DNITmJf4WZ7L
duTHRPo1ON5Now8TF4aFkcYO9o8w8Ws8Scg4gLMfEW0RZzeyjEezjoMMr5AI9/Er
p0ekUV8YJZrF10HbSVzsBxKS9ol5ukFbT26Bnf/HyX9gRK3jdcQdDXYpSO0JZXW8
8EB2aVUUg23+a3nGWJ10a94vI9cy4Sn200oT0ABdi3EvxeHIgWnzODljs5PpAgwH
s37JknlnnARZjPqxBNZJ+TDHpCFPxymqFR2dz1C1JkKxjEHRlms5tZYVZ+L16HLE
zXGmEWMeZ8Cs75MIQneeSGxxT8h7IhswgCxZLOljeOZit8lgR4OPZTLQWT7KRfg5
c8eu2i1IcqfRND/8kk7nMX8XozlvWSPWhtXFNmhyG030b3kB0YgoCgF05e/u8BkB
GSlsbfcr9i3ACQGibyDJBMNPSaV0ma7qb+v3kb1FNd0HgaI9teCwg9jw0yNFYzAw
SPw0x9eMHF2HllPTKBseW0cZWhnC6XDqBdd3nCk44V0x8+B4WZnlPdRlJiSD0QHD
EEuNTH2kcBdNKVHTUOcIedpM7VfQ7bJX/8E4z6/7vgaM9IUvFjybDReNUmvilCg9
ab+5CRVjCWj9Xqi9XWbD+Y1sGsPWZf8xJvBNqgPwtSazAaUfojoEBdffFd4WXddN
C49rqnLpDE38dtMdDeYH9v55eizoTcMd3OFcdgR/HUNLdUor+Gqwdmm8PS/GUXMK
yX3Xrz1MaF+mveXmev450gTyh2z/f+nxVWHEcyMHqH9qBK3fCibgFXgyQSh+x/6+
z0lESL3yH0J3HgHOlRd6W6IMLcUE3TQNhsYA1T3Pjs/UixwiM1YCEWyvBaALx01O
GuR5TVwb4XfMvRTi/uyfKy5LVkN8JMD+qyVbFORuOdDCSLMMciy3pyNbIO5yyTft
/7T/F5JXIwRz/6ZNF3/JzradpFQ/U5FznJERjNaJurpDT+8JF2b/hYPP3AkufWi+
Tgm+ZZvfBwvm6IRA32OQxz8dnD+5zototDnGsqM9O8Q8Dnp4MgxUIWb2eH6VH6t2
u0JDLkSg/DJ6ll9mpKrcEZiUdunvbNVLUkr3zFY8j6+0JpVcUPEIf/Ze/NyDFihC
kry8slbSP4rjPx8MO10ihJ2/AbJT+2+SXtio4gFLaon0meGlfKNYVqv8j97gJ0rI
hK7gs18SXr2E6R+nruy6eBCeULAdEAGkV/k8KoB2tJ3r8wjy/T6tiBbnIhgzCPub
s4pvJ1+YfoY7T/TgduIO4x8owI3P3klfBpVE0Z2DLEDwc9GoWJyxivWS2B6s4Ats
ZSe7aWl1x+9S392vBQp4aFxAs7COmlExkDtjuISvZf3goIVqoFcexsXhs4V1EpNK
NY5BdQhYfWZ3n0KoNhu8kZz1FFesDa/mtFysa0p6Qh1Q1IrHrGO4Q26Wf3ScVXSJ
Dc4IjvgJqOCdxuLIm4WuRbPXTpcnOBGSzuwnoV1uiUup8oMVMPFDpf+fpXoV50E3
uG4khduaAHlWRbOTvaxTP28pGE10/LzzZAkNFDAJ9eopHdDavJcsf4F5JSjgoGIy
MFYFKB62r3GuZsHRKVG/mpDO/7RON3VtxMScVKb7CU7YIOWTOocB/viUpvcLWrE4
TpLjyjqUpku2cQn7YExA15H13CD5PpiubMA7Zy9wPI3oHnGBEsO9bj0vWUEUrSTE
f1t84es6/lpvddFrk0ypxcPgShkmWLB766cMmrnCkTwoajFkGkrWZPJuaUKhomoO
fU7t9hWJfRN8VijC0IO0oXHEP+9GQzGnxhChR93F6nk1crwiWkhgbEH/pxgPvoi3
rXHIAgiAD3SQsdk3OKPLdpqe3s4qD/HE33TVqZG4Ao3QdCXKNIxqt1VRuM8ueykP
r7h0PKQTHZOALES9kdJ0PaAiv3H8AemerAtg65iVUrmYvR6k1yCDNiYQzue7gPkJ
2bqKWBjaK+rrntnDMzdjEYIXZX7mlyILO2cLFiRvDQeF46cLZR7enzvPmGjTB6EF
+bU8E5Up6mVXN8AqDepW4fR0tkeVzTvcF0IyULDPrQSF9MAaUoT+j/5ryaQgKn7k
lu2HIgG796YF3nLeH2rA/FSA5NgAmVBpiVRLjQzq+MPOrpnBSFAPyXkgMP+4H0Ql
AFP657/Dip9A8FsjHfHz8P5M2b4A7X7xmyGIRI3QwfrE+mS2LY1RDXQX73X/NjIi
WG0utEUm3s0CGqj1qUKuK/6zO4Tc++8pdtXFrBf5t251fff3T+r4nzRAHJXj4eWr
af9oEXbuJ+1OlfpGw1HZac4vTsw9BBm1z0esk6e7otGHu3lisI0ynVNLAqfe+8N+
CTtaoPbhUyVR31puiExCWriaCE/gWHczc0n+tNtgaHu+NCQkTDuocRB8PdtGu3LK
89Spdu8ir3ISzm8hBSiglb4VS6JJC462gKCUVro4qdhMCsyA+bY736AppIoMCyzb
QNV4gxvCRsMyYbW6lbzZMvAxxkuirzU5TTK4okF8r4m75MYvuXk/lYGq9rooQfXY
pS1xmCGQlFot3GkCLDCo3TT8mXX1/EMaZmotX0YgGGS1iDRPcUQ4T2EPEqSAcUu+
gTWT0x9qGYhbR+NSjSqr7hI1mrAqr/9G56bJ3IAK72flJ91Zz681pNBKfgrziNt9
PeJAEk3lNlTh3Ve2FX7UcmMvwSHqWQ3e5ePAXXOSnQ5sYSFXBDPWcuTN6Rjb/0wu
JsZDOFNdpyCL0ET4ebsrkEnAkelOj8IzF+CWf3CGVN80ST0YXY+U7QBBnQdO87WJ
utwYseD06fWV38d9OrmGZi0wWSRzPlT0kFxiGOm/UUOs8XwiAqqAth7mK+JzocG/
1+SKHapbyyOxt4YZYxLt7axgK1SMobEe/vY3+9329xtvu1tHCTv05atFBadmq2Hj
AkyRsh2WQBcYsFwMjyqwyqaq+On4ESVIQHPVIo2FFMtDgIm6GD7Shx4FM4oXaV2y
OfCSyS4IzQm8qCpjJD5O3ea00FRFVa/hkarclUntu8zwI9JUUumk9gngTbFbOATh
13AIizRQ3+I83c+5OZtCiWjXIu1KX1K7KTi/5UacIEUDrkXOV+em9lvUrImnPuwL
UjR467cFXmbjVIN2nywCJhGq4W0Tg2SUF5QY4wmqWfbmfWYAodxv/nmi12dJQJV7
A69NMP6Btpco+znQaP0EX6m9/Ba1DEWV5wO0FdGwIGQcubMLrgR+t8AzUiH1Fvi9
KO6VpIlZWSBZ8OrXDVVFNg==
`pragma protect end_protected
