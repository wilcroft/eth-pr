// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:14 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Y0RPt3cOoUa/I7Aq2UQLMM1DP3kgxSBSd7oEozsP6X5e49XXqmZUPnK6PAWufVd9
8E7DdIfZRpPfRFeFGE5xZ61o7yV/tpZYOBYoJjVdHK0zrctrdjCGMJTvqKK1lIUC
8ZCogMF7z3k75V33OUWl1cwW53FsKT1FcPdrEwRR5cs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8464)
N2/Nwf0mLlzM4Pn1tmaFpvVTK5rJZJxDUUi5KdYevDrMY8uyOQIP8665SWlh/tkU
96FDyl3RanA20Icj5AugoFv++vKREi9BitrxyBzzvlcJI74raywzdaD1g9WyeIN+
8RJ2Tkj4C3vsouwjmsRErznBJ1/0ZIUwmooknjU5ORt7lzF/1OPjh3iyWyVBVNPU
07ZgPvAsevs4GC3L6o/KKwGjAajAXcZvg4ENNrwwmuqA0LUGMkxj5wxmMdx73hf9
F4F2yyy8HQpb5gbNhWOVzNBtr52JbCdxmDbr3d0qTpzUPk122H/L9z914BkYSmhD
iyDKPfV6i+B8IYhFT9uZQJ0GVGEaQKtCYEtJXzS5HmOVAZeXwvzn4NTjyyF1b5Ia
0nnZo++tsD59QJkijhIwUmJKwefuVb/+6/c3lVMGsg5yTSTbdH3f/lxB4jm31DjA
NOjFSPFDmTNMmDDtIhEwDY3hlm5r3+G+zacjbM0Kigqf3xWALpPw3edZ8CHOM7dU
RgB96UtpqEZmJ6tQrWAYPTF9V6yePlqsZF0lTCNUZCSOiLK27RpFXAu2P8N1GhnY
fsdNdlZ/PwhuA1HdKLmHZWXWIYm09X/Egx8y53dZ5dDi2/QzMd31S6xpeRbVxKvA
r/V9dgkuwYK2OpxzKBpKA1/RsklqJeVCab2+4O1ayoHE6lLgwIWiYLL2BPyjCKw2
aUrz7F2hVUF1LbPZFHyl+7xWAjrfNbeD87xMdcqMLcYGyQk/1gNy6ZjoLzZBaiPg
rnz2mHlXfj29AzCTm+TuMmM6qIGuiO4if2eoeCnhZSimyJpi0+82D0U7Yj5jXkkv
YGQnMKacqigAFARRMIHh+oXzZl3sKBc7mGucD43NwUfVH2ZwnelABEUo43BDL+iG
2/Ng9p7s7ZmqsbVbQZ/oydROx50LF1fT22g6J5ngIlv/9Q+bsVOnM4TKGFNySkE4
xpHLWa1TJDM76PcftIG9knlDuAmTuRayhJbzdbJxt+LeXb5Ja9CC0Uyj0uBEydRh
lbfsY5iAfa6q3/rTNYMerl9uSDqBQOmG1peTPcil8V5yd/4EMKSoDciSdJZNceVz
yooj21hVvgAAKCcobhBMxU0Y6p63AZ61fEuOYkN1o1GefLKCGeHVgH3mS7y2R3LO
bbWXpMFBtCXttyIfVLj/dAzniQbuDU0ibEMbT1s/eCnFnW8lH+Ft4kNGKdPFZfvw
cE5/IUoxepV6uy6ha0yO9Fd88e7eeW/4flMYUQHeohtk0T96w0oGKLq/SsJ1ht9E
zEiRwwqzjHJgHaOxo8qaSjdsBcfLwH1TtgG+VrVYmeKNTDZsvs+P6K+94Kb9kt3O
t8SvnNFDkmmcUnE43SDBbW6fTkXwiLrJ5oYgA+u0LECIGPPyi2tLxwNAejGlRidr
0GZoWSmXjefjUH2CgW6xKystQDEOA8QTY6ynS6sfd/nDd3KuXaFUIkMUKsX9pZnp
ZUcTdjg8ATphsMCNRQWywGBAqA/66yzKZeXBEY6IfuApUUpfjUq1VyydJQW40vuj
MZOoCBPnUXia1xII6R57vUhXeQO5rp0DvFdu3/QpAZ1gpl0k+Xpytl9vHPXx50QE
s+Jx/FXNqRBS+AqVVNvFSPBSvbqtPO+kjqilvxGAMVS9HbHnWcU39uXrxhv7RoTd
DOZnMB3bZa5pAgJj/2+w464CB1JJf6cEASkm4bNxnGoSwEd0zXMaoehtJiGsrwpY
HvzGYP8hUI3QZnmybL0NOVjSisL6nzB5DmUg8kUAV/AP9ErA/QD2Z049rgiNckeC
VAOYvtqoM85wDecXemVv2Fdm/MpIbdJhdVN1IGjAI6U8oX4o7kAPX8dkYmup8eTT
lg3P4YDlpD+9PdfaIB8esPELl0s4IFqCkziQxvU3vNK45Q9MgDXIOvBJ4WC53VJ8
qUhJqtgCPriksUjN062YaF2rjLceQPr8XtfEoOtZsOA3o59/mbKpJNK3XucXcwej
46Y3gU94JoTTyJ/tEzIcLoQsl2K5LF1GD4uyrA35tC3b476jyWQeXu0RLoi7TuWM
d/QEk4TsJpLisTY/7kLwCJnvJCTybnr1YNBvjQmpt5DNb3x9Io8t9aFceLx2nc+E
eR+pn1KWkhnM0n/MhLCWtdzU5fhZKKhUojQXFNoPinqZJcT0iqUDYd5SYRz7Ig58
jxXB53YryEaOTaQCJTC+rhOdxMV7bNzI++/ObzOeCpj6w+PAXbzexnQiOsyg1Q/T
p/dcrMtA0z+CAGujqFEL+G6GSi2XZIbITw5x69L0yGoeHaAYAMAe5/fVXo2m1WQQ
ayCoVF1o1aqj0Fp0KTjr0tMCYcmWFfLq0D3KDn+7ii9CJ80e0iKI8Ok5Eq1cGWp3
s3KnO3RdBiRN7vGszeYUHtRSuAcfYMzS1Y9OIgm2KsrG2s7aRG7F4fABuEmcZaCR
aUQcHeOvwXKQovpxSM8PrBb+5G+rVT9RBAEXssJmxsa9rzT1HHadB1QFIjXk2vlR
bDCvbctPV31L1K14EZ1U8JPefQLVCkyuECzUX/dO2I2iDkPwT91lBCUIE8uL9cJi
+8pn88CT93hAQ+V5PjOt63PHbMrg3N7imKFlCsAJaCafpvqw5VVG8R4TnYHZh+Oz
DZ+9E8qYmH7C2EXw/SxreB7ec0Zf48Yc6V1z5dmxWSYHSRt63gtSJ5d5iJAlYrhw
cMWEGZWN7OH3LKz6f2y4jgPYI8Ej/UutCp5T4ZP7U3/+pvvN1agt9AvffjCzt0lp
DeSnz4BNwzm+qpCjZ3M5PntA1VGQ1bAmhDAC5PappMUgGMZWs2Hf1ZCck0win4bj
+ZmW4MzgPJgNL/eW0Vf23tBpmh3h130xmRtZzghBQBYZcQsFd2qLtXCudAPjydSO
TOfCdegdnIWcxsey2DWU374fY8LIzuIC8Qsc8po79ujPjI65reZFXIYoeV46qldO
DYpfOA4df72O5Of8yh6SF9o3xzRiwDccmoYEH2YhR3VSX38ky4AaoLbogAks3PvD
pm5S+x4aPB0HJw+MGQ0yjNrJw09PzV4beO8pTqb5qqwIvOgJhEsUL/i93j0jIHoI
YR7G7PwtsgnoluTsBz3uoapbRH9aaAvG+pv1ERyd5JbK+yDMg1GeH85x7KA7jU0S
8Gog5sufWal85tMQvJnuydXVSKCEK1vPfvA2UpjZ1Mhveqj7c15+RryNQ+7ZlTHb
mns6JEcY+TvRW2R6ADL+BX7xN6XRE6Yh+AJNDH8QnHhSM/uc7ag1Qifnf/INikZQ
vs3YybI9iFlg3gQQ1XTc6rqUEpOrL/1+Z7T3vz/o2EA1HmzygAbKlnYBzlUMQv8g
YWjNlfOWEyNGfEP5RkkO5veJPyUIdXjdm2GR7DJu1rJeaQV8GLBORcEhVHemau3g
JFL8NQijOasfk+f104hV21XLmBqw4tbzHCLm5TNX1+bdvbhejE+O43CbT/PP9bU5
iydwGVqs9jCkSXUbijl9I5oGQFi3OYJmLPBjdzntEucKnQO1fsQQXGHpGDdwyJ3Z
LySym0qY++KRSHE3nD5R/dj82n2vWY5HvbPC3bMldnvD4D+F1S8BstMWXqdju5D6
Q48itiBMhcvu4UixaaSt4UmrL0UqFxORjvC8R+PPUUJ1prG4TxrvZg+0rXIhL7L5
pcGW8wL/Sq4+ejxDd2RcqV3mrOUKO/WcMR3YxTy6s6TL4lpFYgRAhFYmibsOdV3T
ikgraMGagCCy9CeAGgFeco8sVRrw18nguq5xX8tJtwgyUfbN6GhnEPFsGHpu9BEe
HHzG0sVwGMtXVpbXsMbnwViSxFA+YLCDpFbOOK3HekzU3/ZLWvQ7JuPd9qByENjJ
+DNvDm8aJ+4BCAMiyWIenN3MPchfg8NC++PqsNrZAm6vAnZZ5hplN3+XUrB97xGP
oUgTH4QgNEA9owODlUpog24/y5O7wiC+eJZwMgIN/zKLAjPwUF2Gwn0b3JeeuV9m
8l6gK1zPbGlxo7H0GuDtMmckzaYjENLVQFBexOBCzw2WzkXJ6VerQENdv5uZIH75
xHs3g+Omhu54ol0LZHD0o0BIQWNx93VynZtHEt2xidzTXTHbLyjDSQ6ZqVCtv2zD
rf2mx+w/nnGAa17iQ+c31ZbitYLnpsAJDpZCepZVIAMvlZcVvA5jTtu2llkjyMDC
TF6vN1Ye1J/wTRucou4x3+sks8PXPKBOvlXO+aD/l5VFYhtmvB1WTGRJYIfBx0+7
r/WnvkyhYq+YiO0Fw5UQZBK9p04qkpzSnfxHekHpWApzifwJbClSOjyEu3tTG8WH
rgEh7IIh17ok4j1rDylQFxzGQ3b+6W9B5VbgFUhZXM4y+lfY4tmHRjpMaszkvO7p
3Wyn2/KZ86ULYcEo3HRbUrFhYAdxhVJfvpPhpjEoEOExeoMjOHNU9ip6mAzzOGaJ
Ef+d8xTJMVL1DDv7px+fdTAj5pYL+pZfaM8VP1ZtV3Jvka5SG4pMZ5F3Oa05XvsR
UZbuWZAI4nA3/vdzteUjPio+z6oa8SqiBnSdBIYcsR/i/X0e5nTE6aO/0IcxfESJ
tbNpuPHpi70fIUwpsdphZnaR2pmCSF3j5XKehFmDhCdtkc6RENaXN20axMjHRqe7
b56JqGLAIR8PYSADXuAIdB7cAi06yItRPO0cK2rvCz/BFuUG34o/qiu4V3WMIl2W
OrvtxsySQZ94zUhyhEHFSfYNIcvzoLyUltwq6uA41R5rTk6YUXCnZRZp06Wqo1Sm
ILak2kiToobhtN9SqVaQM5Gym6445//QE4D8gi1lZnCv7gRFAwjl5VA5N4e668l1
i4IorxFtj5RiMY3J0BXKcJSDVV5ErgxWo5faqSoeF1NOJiUp+SCcv0QUc4g4Ql+G
SOncTc8JzbWImUTYx+pp3ALyVSR1WgAGD5VX5SSPYD7dNd8exVT82iXJh41AXslW
jdQXoi9RDEK4QwgbpFG8vD8xzqWle9s+z+VItxog/97po56M+YLlgv8qMjn2aksy
9YRSUHkY4J4z2E+eCHvHeTQoHL5N36/7L3yl/0P+mhOY9sWcrZKL6XRiCpTZwo2V
xw6eEebcht4ttO7YzYk3A0WHqFa1dzQIXONDn08ZArFrZpAC0vhZ16iimXt1p/Gq
QxbZsvtuPPYYBONIvHH68k16dR+bVZTMi6WDAfUPJXqUxGK+wWOtWpKye91uIUOV
ZUUuJLBs8pG7uC+KDL5KCCahucQwLOHtT9QZMhLCIL6sOtpjdwPMwwN2NBhqSTgc
yRYeqsJi5KPVJiECG72VPeOavuoZrzQBOhviJIG2Kl2qDy+SobWZjMLuuimRSwP9
gFCzYv5TUrm/keUf46eBUuRSwignGtn4jHywJByShuVaWm4euG+SkaRRgN8NlkSE
bF+VkRsII65mDXDvRlYZsRTF3r3p0i9Yh5y7JiVz/gLwnxZb63XGJsfItm9TcXWM
ZKiL+Vkdcqz2kDKirdlyI01en15cIfDpY01GujXF6agDIOEpibfW0Rk16jNIqbLT
ktPSH5eP9WYdrAGo+4O0S58w1yYxiJQqEvr4VZ+HTsxAinsoekAuS0kqOuzi4wq4
pV56AP9KEmUrLafbWYmz5VUI5TPqSAZTXH3SwVL+20kvNffB4m3MOJf8xnKzBNd9
tMayuIPqPt6lU+5MDNhuQw466MlCkWXPpSP2EB41WGg0n2zCPOXv0QZZR2z8h2o7
/6ej6HLWeJPGJjhpRORanM3p5IvxHPZoSVMm8ziXolTBt19gIdvi1anHgidmelRf
dltIQKo0XW34QsD4mJZq209olkxUjfn0BE1wVtiZPKp08L0uu17hNKQolwoyeEPT
Q7jA80W8qdT5gGcUdSxPNIbNPuh/KuJRhdun8UKJ0FD0ON48zOGwvd9PPPzc8p/D
2EjanjRLwgH7nTI1GjJfGZq8xBiWrSn1lHMBwNTRFvltyYLm+xA1js7mSoME6uYi
tdh3P9fePyyIlL0vV66v1LiOKMThjqb26n0K5767J/ywIV5cPtJSSaRF3FDmqLyL
KQ92u5lnIky9MDNKPPvR22+gebJdHMXlAuHbwebARUqwdjAv9sKQlhBeHVyCxvIU
tREjrZS45o8ezcKA7OZMkd2qHpncf+/fY+uSCOMIObZsK+rKS7j01UKB4G/XT8Qr
etTaXXFwZcnC4lQzimPPQqPM8Fp4QqxMeQNXLVk5lur5+MnJNoiF68wJZLFeNr7Y
R7faf3xM3tPWs3ouok8yph0ClzPT5OR2L4jxOMSLKKzRoMq90iTU8NIMcEVQfk46
9dRPqg8fTXq/+4KoA7LY0obGcwuqOCq6rHeSWKRY5k28o4m3U5R+AZ8TAB3X064+
i6UXd5rD/FNUwk06q2ENgM1oV5JkhER4p18B1Zo6l+hQ3dxe2b1UAakuCOUQepXy
6d8S+7QY1R4yeFcfD5VeMQtVWL7tXboaMT4P1MCDU02M7UrN5WNODNoxsI6zlvo5
vc1fGXihrX5skhpJ9m+3jx/00kFHJG2KJhwIufyFha0oxPkZh5h8u/4NIAszGVY7
dx4HqC0QAupw0yuSn33cOyXlL1VjF54erkhngD1MYPXlx6cRFNhWyHIK2JRicFUS
5MIZo1PeGa31XqB7b1eYiZXiJiDksPkyjisvik+2zGD3CbYBRRnNnC9RjlJ9JBlt
AblVZujwB0M1sjbN1rfmyEc8oEJS4ioTVAF6yM0VbpXEpZHg0wPHX+VHTP3dxQfv
DU8Mlyh9VL4sYdKrzn2nHmuZXMCsq2WCWj5etYqSfZeMhVreg2OG8/Otmx/6r5xe
YbfAizUqg3xq12C5ecAk7YWoDNJjumZb6k+OuNxoY7a5LbrDDnGZndqAKeIDir54
Rm3/QTB+gPJQdmORWDfNgepkThWknSqu4LByrwwIvAic6JxomDWxlfnD+0DIedv4
vgd8qGDu5Ctp2pcckwIcT9Fp30hBFJ1enQNh+AUcI6gtSZTL0CZ+vcN5c5m4Dbpf
MiUtqgsnKqQlmJETU+kfRpCtHFdaV+2ITyaTnmvreosycdFTjvnbaZUOgK2/y8D8
da1wh3cwKqoBP+os4FEwOdshzsJv8zDezblkIL2aV31WYL7jGM5GflCCBJoVcGjs
kfCimpevaBDCR5vDd61PhPfPiyQGewfxK9X9v8KR/W7nIE3lmO28l0+7EEgwEHkH
sHb7Z3p0R6tacnFjjgL5K+5KQPhgnHcGlfNUiT102W7dq7sGgNNayOrGTlql0oyj
f4C6XvcKjiVsKBE29ykG6T8Vaee00/0LlwUGJ2s7fflnbN6YTXAPDuZb7DYyN2R2
/nSB+hF4I4XDeVjAN03lNstyq59j4ATUT+qr+VCA+bbh4Ml3zGHom43xXh/ZyQrd
OFMfs7YgFPh0CajQGzhfXUTMMeIA9mYDT+u6wSOpgqhYSFj2FU4a5rhFPLqQIr26
n2imbni6gOPQPgw0dJLacXXDL8lCN/el9wcntgc3yKXWgk+5qOiLeaHWue8EHXhP
Ii6mxdrsZdyQr/g6i+2gW/LJ/7WiopsIeGHtEW05sFxucotGNV+osmM6SKTvBRVL
x+/4Jcp5dH/7GCfuxnRNEvrER4ir6Pg/Uya9WjtcRnqseKs9mL8JWI6MWCBo+H6V
AjgT0c+LGA3oWVUDue1GS4fywZVzqmE8oUbsk+BtgmLAlUtM+8Q7XU5Q8EfqT2fe
yeIbZal50kpjWbS5d+vVu0SbSE+szI3lys6kwsDaBR4+6baT7cmQKC6uXnUnWGAQ
ryU5+emjdYaA2HvQlurnKpchHGH7Vhf95dsBPnxSUKBZCX3ST6csray4IJ0uPhkN
FptqaHjF8rw4SCi+jns3fLcR35Qb9RaofX0Tf4BqDR1U9QNOJUXCiYCC75XR+gvJ
FBWrwykRoLcpNxBMsULXk2kwaNLCaWwB3KvwG7/TmerAZlyJ2u3lHeD48Uy3ieFj
LdKidoydAU8kzXPY2T3+6CPoBS0BYtvlukFhn9LdGyv2c6Nd5GfVLL5sPOuaXmXd
kZEx6eQ0EHyPn3i/bIxa5SndPEodfp50CcMo0R/Ar1/CPiFyTLz9ZlhZaFfOk8+K
RESrLS30i3VkEPzmwxDizZ4WWE4erUY93km4HZdVFrwbPYkCazZeUCTjSgOPV82x
JpZwwtP8/ARn+9tgRhEnAJBuohHzmL/s+j501r3LdlGs3EIQJsvfEWpfGUO/HA7m
8AYjiLQVJT9ArGbou9PiBV7+HvonHBpZHCJAlyJXtZst0xdIR2DD5DkA8dGFG98L
kyqanz8lJsH3i2ZG9+8tWFShcMNDzzgMcRSA3J0i2rJctjFzuzPpv1uQHQsHsWy6
dnEXyLEsO6Ta/BRpdqoHP6kJqOMJrUkruEPYyd0uMGfHI6RZN4UpK95Jno8vUQF3
o8Df0zxsU4nuBP8HrH5IrHu4pW8yUF000z15TeLJ2H6E9iYV895dJ0EO5nUTl0E6
RThIAaxtk2WdDKtAxxiFoCLv/FCG9OtyrOUzFQbsER5Snxc281fEuWLzzzKj6MOK
/EWcJWZI5+eryIjNxxerYi2sE0mGrOtmdn3ibZtNtcYC4y7NQkY9oK9p71inRics
hzSWEtA0SSwPA+eMBplcV+4edXVfMB0EdPuXgMnhByH4HBmQ65FcUBKGIU/RGHaT
obnleElxd/I8OTrqCoX9H4Geidg0cKud/VvSkCieLQApgOIHF4fCiklX8j9C3qLm
+jTmp0bkKeEXR73FCEB3FK0PgS3pDEVfgLF5q5LKoMuuNvONYEcxdos03Ewfg5Gi
IE11YlEzISrhuFRcpAs5B7CjcRrmGQXEZtuMABbP9VUN4L9cpymeYlsymrjPk1AA
/6cYwE8H4L9aLoLFov06og43jazEdW0FzAsqq3l6rfcowIp4DWoTWGrlqK+C8Xw/
q7VYHFmDyG3RhZSgEHgTpHf6cabjAu0RSmB4r1DTlq300Iu5MpS8YB/fLvOa9KT8
/YpP9Z6qEqmtTqz0LRVFVHD/pjRNHQdGJtE82uBokIkOhkMpe/XRdU15a88ciD7N
hDixAJnGCjOSt58ZNWYAR9GTrtKrAZDqnCbTZT2qN3pIMkmqBy2kygZe3V2kyH+0
NI7t+IiGiuPGxmdJlVOfd4C2gZ+EoqIQfroZqSqDy71IXLeANtTwb0No+fUYuzpg
IyjTCs5vqAugwLAB2gfhFEePW7y0dEFg09dyYoZ8xxpLHmxtC80Gliu4OydbJRBl
h0asTC2icXBCjo5ieRSbZOBvwxly0krrZP0N1eqVVWGGybRHtvAPlv2KrL3vNtNu
hYgNlfeRkOuIx/rijoRGfHWEcVYjd+8lVuPCmZeHYwIsnwm/Yt2LCKbdpxaMGKZZ
PkKufiKobqW9o16BIz3NZ6LE8j+QcJlbGHetlYN0+T8e04ta5GW7hA4vvPBZCmQ3
6Dx9G7yllOOJUXF+BsFfJ7tKkt4qiurBuS9qvjZHjEpv4DKsshBnrz8/15WPkUbr
9AVaTZYOlIMEIMJK/KXgkPWlHr3bD6Jh4CsXG1QZ+QlTRf8GFzJNzw1DwB8Hb6wK
X1k4jEtS2Fz+UfN686ZjuuyZYi4sAESHGX294HnZ4knIJp2GpEP0QRj504g1NRKf
SIhS1t5f+UDxW6SysnS2jLeMI6JC0Os76c5qnB/q9YBTrQFuDZGOrUqoXM/37X+K
GT2l+2iZe+VypO14l2Tlha9qUj930x4e6TzFzZuJpfZ5ZtYwYW6dSfwZ1Oppu7UN
6qA5pkPuX/hqukr+LddavMTdUbbfBPcKFVB7kgefV7CEj5xVmPbANrb+DSbi7XYp
ml8r++RnF2k4w2RALjW2tdyA+Es3w7Ms3YhSqY99LmGB/yxLMznNE0HugDiT7VSf
RRkuvCuL8iLvzncSZuiXVrro2u85We5fwjJbakNWlWMpQHabbCv6DWKA74A/DOG0
bPSWO3ZvgnLzf7AP1EpjXTPEs5DCg7oqO4mbNrkFcC2uue22i60GTOcURy/FBTh1
0usygsY7Tu31+Veb5OMZENHL44mxb5M941Dw1c/upGlBcJ7oziVgozfKGoHJvjlf
hwbzkff6GDdnHeS1LWT5YU7MdMDvDkX5+rPwUpZTv8Hwhnf1cWPJoDcR5+tNRzV7
zUZHyC9Qjuirii34QjqaKKCqkWpChvh6lP7YtgYL35RkPGyLJlbNCUsWdg93bNlC
/yfFCvssH7lSgIYAJayWNIVN0RcePDXyjqH0FPCtvAfxP9VklKw89QgWSXjpRsMH
mdJZPvlUFnqCuKFCCmDIuMlu+rcnlxTpsaG57232U/P8E4luTQIfjedOTOIiVEkw
8pouE5nDBMYcZw01srM2jDTfrrWasI9mpz3RFuLvMmoyrjjW3l2Gx4kLKxN0GkoC
o2iTUPSVV7BMReq3tjw+KzH/ujeqwIwCvvxwVFy3GyLsDYOc7+nHClZV1WTsnGQ+
zSVX3rEw+W08V8vR5uUOgR1CviaFxtlh+mqLBlly0WAxFKNbh0qZ20VxTq6hOP6s
HFy9XW3VyMRV4Inj2c9NHjsQiFel2dwpNxNA7OmKRintCV/q7VAhY3VttvSHa2Oa
PkSkk7fe7ESHjrvTdsIXmlNaB7D1Ooq6z/AfIYAG4l6QQD364pkoVhRpQ2fbGX5k
6pHBhQzv7870ev3qrNE+s8vej24DnJsxIfEtN9q9yZ2x+qFe+7jLTNE1WLlgZ5WO
AlQwgEtVEBAWw9wVgMH9ZDjlXxR1TkFvX58pWepbpmSlGeQZx06pGHKU+uxivh25
ll6Z0sgPgYx/AGwdO0n1T+DMOfRGB9IxmVnwqtLdhMqT8nyQaWrYmz72UrWoqyuV
pPSTcGiGqlzyohTUpNOu2G5L+fKUkQCwuMwFt+P2Hrn4fNTSyesLBhGYO9ZuHJW4
SrUGgP8D3DLkKrVD5Xta3gSLqA03a6u0XonOzmySgVeUu79QbbKJ0MHrojdNFgfN
+1ZhlRniPy67eyLYTfjjbee9E3YawWAeb/BoofBakaM++72hqvNzSz2ETZUKlzeu
mN0VCSPsewKDiQmCo6hzf34gCEUop7F0uAdmmJ88icp+p297OTr9u2nJfRxMUDy4
d6DBep0oTYCpezT/ecztDbkKd2y9hMs4bZvyv+rEoNJVMP82ZpqWz6RRri5/qIdd
q/vf0fC/o+urgF9uAJgMP/rErDfmoD/4LEgAbVpHSEYRqBxAQbwExco/ecT8Xeuk
J+vb8c4okeI4liXkN9dPTzNIL6Y8Xspz1wbTfrpd9wUQLuTm/a6Q1GGGEeoG5Q1E
S4jhbVmReFQh70lwSIuYgg==
`pragma protect end_protected
