// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:14 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PsWrknBQPBFt2r1BId5Vy6zZnpK2POO0pCazhNu5f4ZG5igMPPIcyOORViDVGXES
bwao7igkqhruFPfpxBT4jN7g5TUjIfozZhKmA6KbRzzHj/drl22hwe4xnEhY0tGg
WEn1UiLF6gBUOzCYuOBLN0nnAFxDoeYeX8EBXDSqm9I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 128304)
Mdkqzz4l8Xip++I3o28TbSuA/kz47ilMbosLbb3onuA2ohvvo9ie9VvOe8b+ayca
UlZMNltVuI+vZa816m458khim/a366ZMG374SAl2xpSd8Jqu04lqIuNLFwlC0d3s
2Lt2ayiLsruVnznrKuKgBdTMubpTeOGd56QGlbtol52UmFwqhRZ7VKxnzMHZeCg1
DX13T5dZSa9zt2+8Dlp9WFWB4KFTthGhk3b4g0HZQPZKZbZRpp8sDOOKcLOq3MNx
RrYnuhrIFiy2Zf3wmcqPT6mmG5nqRnyBOpXokohiFZwVzeOEaUmB+3eS06ZkIJY3
8ST/qzf92HEabY6Ilw36dURbfaEN16NFVrLphpZfnNAvSkzoigzz/KUCBe849LCH
V/tjXKcgmU7AiRTZJvE9xD69DZhBX7+S3nQ9WpWGJazZOU+8x70UwT0HRDs36Xoc
mE5aPqb9GJ7rgetKvFkfivsmlR06bof+3xibTub53gVt/7C101us/SrPGkwjtyBm
tY5oLpSuA8CiYOsVUx0h/O1++9Hv3vwlIKkkRIFM5IzmGZQLaefuQiIuuh3/8Acu
orvqoP/KKFu4Sb+Or9L0O2+ILndBbjwAGv/eWKEeB5+ILQzuO2pBVxKQOC2eGmM1
GB/WaXzKYxzu3h2wInf/RAhxcDrVa5eaWsnWfF4VYDCHP/xvNupy0TTjl9+VcQd6
/JDAyLkM97bOMhn0GEn38/5NkkpdA5CbGYyC9FhYEQpvwRw2csUqHqvM+Qy3FNM6
X2gH7jgsVynPbazKfkCv8nyMTd9i5BqyXlscYl7/6Gu+XBRuycPX0s9En5R3SSY3
GlkD/30co3QS6HZ9FF8ZmWeYdzQGogqIViMid7vYqwAkj+oImk6Yi4UnbnyGkb8g
zPZEipotmakszGQpln6hnSrphX5Vat1Pvjw+SZ5Gv1Afyzglq9bVc1HjJO8mmM5w
pOagH888hShxlB1u1eSFwbiYqTbO8KYrKDymrjtG8HxT48WTe0erzo5vNYq/Rd8r
lI1w4OJoRiFduW1XlvPnP9GtZttKkfr5Jv5bx6Rgr/1cORfy1pUjPzAQ5DffEZYF
zJ5mUOnhUfB25ynO2/kc4dXIDiuVo7ydkLDmIGMxyhPzBfvBX0fstX4VOxTeJQUs
bsUbLi6KpEW+cPBZcb/jrZYELDULylqE6TXZJD+lvI2+BQgvNS0Bvbh1HUpVfWwm
A8pSJcLkzm99e4mU0H7yGyicaVUyk4vulpyuWRs8esF9Ou3gdJRoiJ+9DZlNBo3j
kD/Ln/fq+n2JDtky2eXf2tLt+Fv7M7E/E0VtXAA49oYQhK8FndpOQK/LmUdWif48
v0FhtDwxpyp+7kLAgldYJM3zlOuK/k0P0fhjLQmFlFBuzRB3r0p2ffly9Hvk8aD2
2o3FH3MRgt3pt3PzNw1Mh1IBPm7T37rJBLZI4A9uF/XaWL6kmDnqcHQGIWgrA0Fb
kNv7HZvGGw8mZHzRkUQWujI0/CoGu0IMlTp0p36RhJ62w/LvX0g93y37ETKjqqQG
98E4nAbD50w2kTeEIwySExlJCXTmeEbgO2r6ujqbVhPolXCVjwi3MXx41F87WQ7f
2yYW/bAWI12IEeqctFfuzFDKvFC6MIe1GtmUsJMPqudgvqJXpPUTrkYLfwGvDjkq
KdebH86xpyPSXLcUAh5QyV276i8JmJluuJ6rNJ22FKLp3FvZOEViav5f9LpW5Jhk
IIXwYBjbV2k/w/jac7qtVUBgYwXTparQ6lZXXhFG0hHYq/30xp68FTZpHWiheKjd
GFpYdTp+6vclI4rghvP9m5To/40c9fC2COpGjtqyUG/pvyiKvEv249Nt9mr5TIaq
rCA/KSKcBg/RVqFizv/j/O5UmYGZ/rH6tAk/pqzTyO97yYqboiqrCRqzpSn02aQk
dYD1J80kKRkvm7Iuzw2HDvKKbMpnMb4Fg351KtwaLDxtl3zCP/lHcf2jsfsb63jW
PoxOutaELXwCA/4h/Yaf2hgNCmObgReHWDrUlEWSux8u6rNpJhPjgxBOG8MwwfKo
rnXhNSB6UGN5u1PUq7R8yCiCQOL8TDZr844iKCO4Fy7KdgRTN/vVsF5oXiZPybRM
DBb0RSoAJwUVmTQJEHrUXaRy3SFhD4lWFRl13qNGz7gfel7jxhQNw4DkCtQ5FBSs
/c/DCitifozwdUIBCb0IkKwzUZv7KsPIPn5IDHLGb0AXvXQ49+nUJpAwGBuSrjB4
6zztnjEf6e65WG4vmf6v2QR648hn+5GobBlD59I+NfINcUpNSgnHvaaec5gPG9kL
Dcepbp+1dsV1BtfyGb1GF/oDd18HvRe+g6F9G2suvgxw5B9RiHEwIH0A34Hzir3k
JT2FdUrzU534q1X40jCirgQyWcxq3JT1i0lMA9rcli4PeYiK2JmSjZNh6FCuy2jn
eFkpg5AwUkb4RwpRwf4Zg1begb2XeEdoJ2gKqHqMngm8GlKx42C06oWU0hZ6LE8p
Iu03OLwPyPquzZvPK646vG4TH/G5Zi74x804Tf63bwWydSBh3bAd4hzOdzgykgkZ
PsrseMV7n7H8jcgDajT1RYVAhJzDJCfv/AxyoNnwUxpmQvKS2NA1DpEiLYOZYYeD
EA9vC9o7i/Fy99zEmxWpnkiuuaT7QSRD2YKR5otQYP4DVzcYy+UCrYmXSTnJu2o+
qnQK4C0J8nQUk7zfRMN7PjJrdb4rqx1WR3m31pbIKzf4ojGdmTovyz5BdTMhZ+Xp
J3NGFFoDXTESM29WUlkPWfTIJQbBNLPuClRUFdm0KxD/wmamwX50NGJKzCFbgHDz
gKyqrYqhHjwzpD5DnZSzgM+UHEORdXakpPdefaV06ynfaEChrQnXl/KSQqmFewsU
0Or2kNVBVWgDWYcXTqXnuAMniZq60GO3TSswkaTumLebVBWENGPC1vvfuM20aAIm
GeGRQZn6yBzn8cQS0rtsAeXKUv1xdNwP99oI/6BoWERj9q+pX7yMzahdnjsoMUij
USCNRVi9MvK0Bn8qQglz4qYRk/719jF1t7H9ej6+XKTUipWC1CIeVOeHx5tFXpmy
kdUaSfH8j8bvkheYDT20Q+TN5sQRVs9sUZ4IXMAW0Z//tARJWXRSHuOKek7s3GAh
uvpS9ICPYQECLgZdGx1p7TSWjq1l+sA4Yl5Oqj1e4Ot1b8/TyAbyY8vyeUNLdE3w
F/MvOpe3AVZMZ6iUngGELRp8eY2LmMdSM8f6XC7CkGAr+vpb+lNT4VKVkqdpNJLF
cg7kzJdKP5KFQkFSab3kcyDKgeI0OLDsuSNyt1VRdxFaIdhziiVZBu1NvtjJlx8y
14KevNHBNfuLVwHl4Wg+2P+nGW2s0SKluMF/AU5umotd9f5a8VAWiV2W0G9LQp3M
joCwYkLEYnxqATSCdgCCdWlhKEqyzGK45JS4UsmqOTmvSGgzKFb0Sv4z21nbUw9s
EP1jKnF1aVun9j6gp8/aYPSh9+yI/Jk0K6kslwqX2wl36/AuXod2pi8aKGIrz9px
x7R1N7yzZut60d8PuMzwEAy+lDM4nlGaBK2A4sCj/8+GqhmMyJllum1gMS/OMEE+
TBU3igmyah5lskVkkkhJfieRJ939vx8YrdHV66mDfG0kIeWnZXlHfjEdKHZ1LohA
p0kiJ9GbqT0KsSWlyhqYLnnWMJxxVkYoNTLXHIp7acWVrxbYovdCvWkCC5R5oG4C
Us5TB2xm7Oxhbk9aZrvzoKmtLIAxfuHmLZ1VaNvx3/A7BEUBv2AFWtwExm3CluVG
J1pxIq41DpCz6dEYEaxtPfqq/XFssOG7LVy46loryIYjDsmI2XGL1KbLCw9xWHAt
wWxuDjkco6zIoQlWCIv3VbHgxpPzkNb6YFh3BSQdm10MINAzoX905jzQSbzOppS3
lBoFEVqPBBynKsx9AVxqmk7CWLiOPAzxKmCpMGPTM+MvREtuugxTLJ98SVpYJ38N
Gv61YIFk92mXAec1252MPtOGYt7ePbMtTE25QAsoEZbV6fNmRf1vGZ7mFDx7wMqj
E/4/klynPTClVNEoFXHMP+Q+Goe5Ojca1OrubqnQlTE3VreJWbfaWRhNLVoSNPNC
9M5zAnQgMuA8FpKOmuo0ymY9WhKAoirAxhAFUfi1nkVv+o1oL4wLiHah/ApZHRBB
nUhjazg1evfkwxu5RtkfimtwDZqtw+mixW64hLisrA/iVGqfPp0ZKdKb+BJdxSU5
BLvTZY1/SasL0dNxScRWYSDvWwm4VPTFAjMUd/L03MdAA4xiA4+nvrBIOr9p8rh9
h04Fs/yBLFhpPAtA2snML2v3GsHLokxGuqLWrmwKZHBhAo2+HO7X3N7fyXUTxjbe
/OV6onomEiZplCH1BMU3bbHmrnNZfpXjWlnDQWlxtVKw4j9gc4Cx9LVjqzVhsg2g
UUNSfGQgF//W1E3cbYiBqSpFYYtv0r87dZTFjZ95CAjv9J986pDQ/1OUqKh1vi/Y
pd8yiE9vvV3icGrYYaRT9WiE7RC6gfbTwSvDWYrz8zhiAjuc9XcjPCRGxw2OFALB
xwc3R1QBaLUG+NRbPNX3hrhqzKnZrYvSmoJKLzuHXSTnmNorJfFNJq+Dvl2QFmCh
PjZmkLQZGlgYiMQ/O+ix8fQlui+wsOnX3KpgWbA0qFwGWuWLSIqo5MCENMqsPTA1
ONJLomXJmieaUAYoFnFZHxDMk+7xCgmdkrViayGvRbNyNihP69dD2ZSZprQXQU7N
4wzCoqy2UOte8n6ydK2OgQN9zgLeZbW6+OL5mLhr5b51qaIwzq8A1Bmh4my1YtoQ
vTjLvC5auTcI79olzdB7CSSFU9Tbqo2nd400PaY7+hsDrKASjA37AVY6CJ3eyIFz
33ZWbfagGmEDB5TYitL96iNBSbm+fzBSROZi1KU0+rntVSOJ2icXy3x2X5+OGA9f
/VhyaJB7WaQePGjJ+ax6/s1DEUA51XBO1om2j7fModVgHP/Fa0X3WKIGrC8LLHoy
l3bPMZimfl6y7hGdH0Xz6WF5oxT7kOvCOABCD9uO7HQueV/4qFrDkLVVjcCtRMXq
klUGcp6cdddv6UuaycVyaQiVxnB2YcHKNLjCBqVLF1mNI/woPwAQag0VB5E2mkjA
9X2HZgEEylCHX58R9MNWhzXP6hNJ80u41ktKVcBA8gb2O52hURBPWjSZponioafK
nhOAObks8KgtCgq8Q8VNfFtpxE7JvArhgXO4uRDu1DysC67j+FrRciomPYREKL1F
g6/MkioUtTlrvrUAuoJ2Mg6yn0PL5cxLeHCuLoGMUPNO2NAC/T+biZVGnamInEYt
pc6HTT884nbuFiFxAEIGb/hXjpuZEjWf7LNErg2HAzxRT5ZXe6pY4sQ7nM+2li4G
cArfY8kL7ROivVNOXJcP7L4fHS/ciBl82QLba5uJDqvkY783GwjEvR0bocbZmqIn
TaCg7hYfEiQv6BY1ZI9laJQPjX6jxaI1+dBx3bleUQcwnkxK1I3T5xq/VdMKsfwF
2zGEbv3tXX+QXy2GysTkvYfREj7GUkDdYedfgnURQ4XIsj5fPk5zgR68QokHJGqP
7z9veggju+xWNd03RnqgSXiWEnV+wkLQpLCfYVy7VShrjs4s958WWe6IObk3qnpk
NcquS+wCZDJZLi5lmLyjD4N1d7GPJ69d6dzk5ImhO/1BwcqAWNrErddYp8WgpUpE
Z4B5/b+sabjyD+zBAzbMRUTnOJX5/CW/7ZNv74P6tmBeTV6I2rpasgBuHi+Yaq5S
W5KRh+sx53fYnVzC8Jdw+WClq8VpQbnAgn+01SqBe4azaOsieMXFHhTrdhsWfUdK
Zj1yCbSNyRedE3stAb+cbxou1OokIkCxKiPokJ8Mk+R1amCF+ULJM+ABdkNnxAp4
H8/tPqeLkvOeIzFSSp/+ZtWiTbAyvBEQBYuQ3ItHZp6w4Hwk44ARWtoGZHjdpxDX
wNX+KbJs41iQW/9y7Trk/SDr69z387J+eAmWsu/Zyg1H9kl/dhIYM2voW77dOR1t
REglK7UD9FHlK9+tpF2o2azatnQpMsq8/f2liS1Scd2iujufyi0hWqaNYkPFx9WF
2VEq4k/p1KVbNvSLb3RRMUqUD20KyANX26dlCIvNd3KMPeuur11bdsFW3wZcZtRU
4oH6+bcdZLeX2khW35RZvk84SC9OdoqLQurh7RLC96RcozfQl9EQkwndLeqUY/8o
NabB42JkA/Cy8jEZxNDTEIBtPiSEWH5/9bRdSOVFs83yFbeWUUa9y5CTLUffRpKi
NJC9GEcyBd7eicCjG9VbPdkEd2l1/QjGGrpgAT0V0YpV4Q6HTnPvB7LDTLSbwqDn
Cm7RwkUkS3bH5lSDJelSAK1Xxs3T3U0xqgj/eD0TMht9AxTJIJVfsiUjtxqbsQmq
c/1ob7HAiU9PkRVfEBfXVVKNP3YfPJph6S/N1ubYwC7OfB6B/Cp+jnshzvheoSFN
gsf6vwawJRAlIEYv8jDeK11WgCZPIK6JnePkMwlt1VqgdtrqeX86Qg+Ld5TjqMht
48eKiMaYwsoPXErdx0aRUszHW2OJSj23TNXDabvInqXeRsNt7Bdch0go5NYgwwGV
u8v6Zm+BNj9dKLHRQOuU8UdnbzMYEy/KxQeiBYhv7SwNHfUQTkYhrQawJs7skwr8
wKw5nUBMrPMwfzPc+RdqoUHHt8EymhI7YqkUSOaGR+w1B7Uu9cp8SA0Y4XphaFpR
XjvyGQmrZciBTfqrn3PLHP349NxCDuxrkLepnaSmuzNYukYUGj3mrrocC9sbhAaT
Hv2CB9la8lX+c24s9GdgFnt9eeUdL+3men/RZZw1NTuQ3GvJAy+a3kD4sCdI0pJG
204uQRZoN8/0SjvU4Tnb5n8Deuwsl5qaJIZRBZVPDRiTTZjkeObtyDjKI1pZ76D4
Q3/AoImmyY+/PAHw4lkDMA3DvcHCmADebb+ZiozoscEXkcFa6nx98WDtRnJYqMhY
/aMFF+5ZtUY2hwRWgwgL9NpaKE4SFwLvDBLm2WEvzkdqaR0/MVCAkUX4YnXgs28h
2uVtCuT/A3iBaIau2Q0UdhSRblcTXFDPIUuFip8qe/fG/u6zC4yUgXWdb+N4rP2E
5TKhohmm1dsbWvcGYYmSp+Oy9oPRl+ozvB2xmthONn2GDhVRZ7e57SMiM6qCIUOY
tMX46RRAl8jnMUSTysVurkK+9KQQbdrkli4WNBU+qtWeRj5Rz/+Zw9Wc9GSmulaA
fyDXwR3zPkJT7OHOMZAGJg2pXuF3KbT8XFL42E+WyXWmtyU14m/4cQ6WWL7+0hXh
50nzz+5XkI4B1mnn2QQT01SppQ2E7THUU0boEbv9mODq+Pppcl0BsxuAJMcy8l4k
QUOZ1701hECrm4D9wRiaJci+BhIEJxLpd62BOavW/P9oIWgaCbNwY2wzOEF61MFx
VNtauM1mEpkznlwngWsTEjpk9vXSKC8ERQ1hNHPSj9vIexNm0ybwVBPYNlRE3+hg
rCPt4zTLii+CpMnUVDBXudDQ+rTAfCa01RKb2xmU1K8zC5QhK0JCzaAOXG2KwjLt
J2fHNFzcoj8zlNBt0L3/H01B88SOGNNd34iKgZYBJTXHkKmQFM++jeUSpJbZ4/do
BKBdFh0nqyHiw13H1BNQRvHBx5pHNPNO5aGqbPEQcpkoNAFsRxbyPh6fO0JAytGq
/ZMbJ/Up0DizuIB01Irp66hVGLcu+kq8wYxyfyLAB8spym6MkX722ftGvz1SFZWN
ZGBzhNP0APzrS0DVlW6RAgndMjaI78KttZQ4V6L7kc1kye+TmTjEcOC6R1kVCMjw
TFZ3YILNVevMnfFkluieMZLd0I7PLoAyB/SOr/T0JGdPkeGQLYpItHihy9oQ4A5X
Yiji5ss87NA36biA7zHVLANhJuNi+TK5I2TcrEowojol1VBMzX+aofRCy/UBBBHd
I81DBdjuolaTz/bWZvlYNLiZ3GKV8m38W9uEqaB1ZbJP87j2ud7yF0rng7UpZigd
AXRYW62lT1aLDzRZWeRVFFUQvaIz13f7mOASuTQLYi3OzXA5YF6pYz/m36IgHBv8
FRU2hSAWXUGzQ1zYkr+3wGdScmc4cZnrc1V8sA1/gN2NwVjlEACbqzqHxEh6hoNy
rnchBDkGe9vBEJwapGyPaSihOdXyIDPDm3zjhVKV+CWkLoXzfgPDaWxDnhqHkSxv
xFrj32ijiOxDAjL8UyEPuyqgxUJtd/qX+AsR8DUzF7IX2REGunKUNtc5OiExWc4s
KdUquvLUelvcI188X/5qSW1M3ctYHDdlrdj0Lr8J2HzU2zHyw+p+vDOC3Etgc8nY
ucQPdJVWy2mKGn0DnR03UoaxMI0g9W77dS7D9Etr6+YONmaq019rcnhb9cJQHH62
yRjh8eOMOqVoWJHCbANjq4S2JU4gRBbKUQ+z49OLv+R+Z5rGtS399qUzHeFtiWzX
CCTABvmWfkaqQi/AjybLcsXVfilTiKFRXXL/tgmV4PtlyBgfbl0T6EFQLlMj3YK+
fzMdy0/310bZFxYJIT4Qr+g1m5k9AvOeO1lCNfkNsu3Md5iyY00TJlMoHBU/je4a
N2njYBEkBIgBrL7/+CaWNndGYpa+jUkw7tIHwbSwvfl3J0bLot+Dig0DHCiOghiV
vpP2y+YqkX+xQHCc3KxpelsS3LoSljMMyqCG8NwmOKVRWrOFqIP6IXTA43lR9/SD
NQ4lfO9Eb5CrU02ng0+RGqtXkhZqhBV7YtyJnWrvXZtqVzFdaepw1U7qAJepeli/
pz4LXjx5uWQBZWgU96FGQgHrBKBH/B+PcQRWj/MUjiVfglFZcjybbBvmBQjyWPhv
bFXb9MjsmFf3Oj9YRd75woZR1jkmDm7reABD6spbcMNuJDfMlEl45RXAfY0PJmwh
jzkDCJ6AFFUH92XI4f34TujkrfYHV6DoJY++MTM8ZR0d/dC9u9C1R07t8Jm6PWzI
FSMFMsujJe3+sI0EgQREtzqEjtGlj0+pigoZsUlJqN83TQJ7RA1urN1xOrmco1Og
TTlD40BtKjDpVzyE/ieOjZTsRUnkO95kjir6P78nZCI1JlTnLMhoeaqtBbug5Rbc
RmKiv2QPfw20BskQQNqdTVIso/2la7OJbYbkzSZ7spjYb2uLOXz2WHJM9Um0NqaU
hL5/Wdb8tLiiB5JZUebXww2KOWyw782aBAh6wN8kcC/Inet/ANcxLDalC58JHRYg
dRXQtysLJ0hvNHoUl2dyVn3oSNby4I8Vn1qgbXo2qcfgqqE6AU1Bs48tcyqJP0DO
YR4J0uyVuslAaJYmcTvVKmDa5Aq9hqhc+e/iCOUW/u4VMrUlKZvh5pnlJaqjkcC3
G1FEQ5yGleDaOhiNRtD0oRLsvSsdOTvjn1WsjozA/Q0uNDVXPNyPqRAERqw60k1m
KzUGqZfaahFVK6SL7lEr/g0Ghst8HSYSfzQIW1jGjcL2Yb/GRqV0MsDjd631Bt5S
P3/1VXJoZjoP8EQ0Eh9dL8ZRdTILQ1HvRyvIVnyvRfpdfYwfalvv5E5ZUzjGyYu+
PX3Lh7hnMiytmgjebW5DGP2kBwt5uX0KqpTxoxyVka2InUfJZ2a38KZH1kL9lJ6k
rVfTQRRU2XUik0E4KOo0aUP1nT5aKZDyu7LiFxctqrFHpCsMaPsEo7N9unPhu5Pv
vFaIVZCrkgqWjED2mv5Y3sItqAoHaPRJyfoej6F7NBd9xfwirIJcbZczAZTVV8Ul
941R3jFG6xTEDrqRWdfcyda6otfsKOezDRFC3mLQjOorh4OkY+i3PdCZeSVThhK+
/iN+tUzPl6VJ99JjEzJB9uz2lXZHn3JcrsmBuG7fyK+DzwWPKyE+ycsXFko4nTup
W+5PHIUtcomsV6VavlCmpoihpyv+haovmfMd/xS9Ko4Y6/EIDg04deWEHFLg6l2X
Lug9jZuPTX/TVDVQzdrUIcEmr5n2Nr87wUEGZftfYsbDfFr12gCqjpUHJCDdlibG
psH9fIIASKXhwqN3Lyv0/32HMWNEhB6Sj+cPESZAGJwe7tMBKE03VRuonxhD+rXA
j6mzNkOO/NG48BRcUgtrfiDyUYnF0QEmPCJ4qZBFSX3MryPJn+tQBJ3crF8JclYm
qgo1MS0pwz1NHmxK/TYBpqR7zcsW84AlGIpaOy5HTWIwdFZggg7VZ45PxH4RSxwx
Dlvs3lRKTRgyLvfw3wBMqCM6KJ6bk/QHMIuloVKbxvf0iHH0zkNlfkFytjde+1dY
EnUaSvHe8sLMI4Pqo6VnuRxXzOMTq1QAT4rt3lJzxeoAbIlePO7bKHto+jWwL1ob
4zyd8IbcX5qjU3/daPa1yVwktCWZg3uK4v+w3Qyv1xZmjsp7JO52oJ2OW5yz6m28
THCHSbXHRC2bEo5DPTIiCQq3/mlygjPDhPp84gfSOqUOsnc8IiMuP/Bxx4CZ0Yzb
nvjPtnGDhU4VK9X5VMtPo/YD/VvQLYXOI90t9Ogf/5RVyzN3aZdETx1qbvAlXNQW
4S4cPMY5CP0u00+HLTGXdHocaA+6tt7c8EKMGF75qhtrGxFpYjyQ3EJBCZSa/2Gn
jHCCDskDHkHl2uWzuioF7bp4IUZUC20/LoEJHwxyA2ODgNrNGkcArXpdDfMX/L9+
JK0YUlDiNSi+iroRZto/U7hDI86sJbcHazRx+x3oC5OOWS0fMDo5v0js99beYHFo
ljZlK1ByF9HTQP+RJun5S4oxxN99x4Xbw7AbMYPaCk/XMvDNtfyfHGt1m+1Y8xu5
mlYpzuU4/LdRZfU59k2SXbxJQKzciX73dF9T5ZHe6FG/dCEhU7SZL4TaAwrB1dsX
bfs1K84NWaRMp6dQ/c4SBi7Fc6p7WVk9NDmx8tEwR/AbNc0EHcYQEU9Hu/eMddB/
Oxc8Ep6+uijM0Pi3Bi86m4W6CTCkvYvRivQYg4Dft67MMw0zt7zVUaMIViE+Royj
EKUdqS1EFn68pR7+ocrcOm5gQ9nZAhlclKDMIFk/b6ese7yD0iAoUxbLT+lE2Lvd
hFsMjbTkznFuIxFQnRZ14gkJYEL5+P5lnD7esjcWqShJDwrHTRjVSTH95dhy13I9
ynLvCQU968F7ZYB/2921DfstyqFq5jFd4apmb+z4LXkRdl8raEYi3L4BZhbotLdL
5e4NgXAjXW2XprCUk14hvzKaf8xKSeF9RysOTaRnZV32KNDgPrBV60pXNY+YL6V/
U+PKaTxe505k8TIznDzQOTQhC7QT7kyT1V4Ru399jueImuW4w7J6Yd1y8oH9903N
b8FOfzrByRRtGqE+N/NRbH4dz/IJNPOdq4aVfTGG0yOcjULppmk911gePzXwpwrm
4gmgHmHY1otml8i1BbpGkzlJgFxbPuT1TYPcnsup/42sj4p1HdApRIMVEn9Oy8hE
mCHQhPgFe87AwoXYZd+md1p2wIoOsY1Zt7WqJVR5eJjPPTtHCFYGz3xmcvHU0+uD
uKJ6H8VtWfJ68wymDG3nmx7X+cnXUqUKFoTveXU0zlm4bY8Xm2JCuRwQbL946iF+
W5ps6LfsxS/0Z14C3V3ppXoh7K11/snOTUs5fPWTOU4mKtWsJKxn/kexFCdKGFai
XPQGYJBURcBLE+YU20E9jGclxc5qgE1w/9gPiZHU2rrAhi28otQvGAHtnkUcSSu2
30ZlaOm/aj0rhkOg8/yh2N66E7ksFgdgqrw+4MeJlmuKmhjq09d23i2LMMfjDoIc
eCVLM87pohYeenAvAT99fAQlKYSD9a0D5PdMocWM7TFZ3m2JZV3wI0b8pyu2vXY8
19C665ovk1rQBN3yYrs9HLEY+hwt7JLWwqTDfiUtVZUodov89+ITto6DCW3M3j6F
qE6agdpwjnI6E3RgUfqFvr/Gt9ZuR00QwgylR/7rc9PrASAlt/+kXDjv5DghUWjO
//AoKc8VGRdApJ8JFXPc0bublKd223tZGJ+AQESraL+fMUzbgT0nijV/RUUkIux4
3X6WFESmgdDZ/HyT9ZEIPJGejVpJ/GdNX4JPGGQY1H9H5OIc82p5D2LuyVhasa2T
LAtX75ICMfotmQQMklBkP574SYTZCqeRYeIMc1kRy/i1hWXm5ru/E4YZz+c2vNfM
FJ2mZGlPdq0tJnOas6O45uN+ZtbH4hnmTyyNOZ6GnhDRAJYal3IrbSTyB9Y+g/HJ
VsHWpuhydxNPK/FLJElEVYMPltzmhhjoCoxr98WZlytJLj0BkVmRMNQtaFj/Fs+o
ZXiMQHk0H49blx89dW2Qh3EhDNzGL3WZZfbyxDFBhOqMj9VHYgwFCtxyujrBYHum
eEAYfEQnuY+vqkZJxegGV8RGhS9yrpqRbsYBG8aDhV37+FPR0d6ueNLbusR17Y/s
1DTWqVOdzSOHNtYlIm/vNNHY/KeQeikf3jW4Go2RuaA4oHGS3FmsJdZP5cKT3NbQ
wEwG/WAz+pHE0SPZrBonQTI+c1rUQpoxFryIZv5IdxaqPQ68UrIEQ3i4HJNwyIyL
c/qliZ8VOlkKrUzDQpRGtziU9OwxJ9wmIDyHVW0b2//2cWgl2pODipxdEB4zXAAM
6zfRy9UDHAsfZ2TuSqkUiwy0iR+arSuqU/O4qrs2a/MBNnqfxJzwDMJoKfs0s9zf
gZOIDG7N+//+iffsd6+p6NRICynntSVktZ6Bw727L/uP+XYGHwxVzDAnvtrzXceM
QPEp8F98pTC/O2/5x87JXtJE/p1Uqiw286ADJkb78irRm0IDLbrGyKU+LThwI//S
OrdSn4p8JUvTRJoXXgwOgzlRT/zCBl34Vbg5LV7rMkFjh7INTfFYy5nGY7Q+pnKD
gZ0YZZYuCtYQsC2SsOz8jQHfiOxmWDp3vJTcecPk7zLrjzUJ6auZb2j1fW9DHxV8
8GB8j6Qx6/Nc1wlVfrES7GoxaH+ghSdzJvrkFACSw2xCb98JRiyTooG83wUSaVQb
mRzC0/J9TCiqQnXG8NGdzQkJkbeXuIUnCYF/9fmcykyzcDyTtc+86tiv7UkCARxr
rxvyFb3tO1IJKLN/lCU3iRKNYJ+ABIgtaPkmjJDFyWlS/Ay/aKqFZFL1o4DMQUgY
ofa9hu580HsGDE88cmiCyNX4ucUgEkTdQ3kzi6QxeB1iQXM1VGTdnvZ/45RPtibw
E68SUYMiD9gupsNy0smALARxSuFSwNXrOdJQzgL2tGGm/QgaUz5lkEL9nMmYTy0v
DD/Jyleu+/oriXSwjDUziXW01NYKlBT4Og+qJi6JaLmtr80KZ7sJQWtOBQtQ4QTG
vLarGhe6Rr3aSWl4mTaWYSiegmnjXbv/Hy5RgfFq8NfyuloGSEc43aZUHS9NqehG
QtFT1cOXtJprWKWLs819UUWb+h5WxcYTP6N1c59OY5KmjdLBaZJEOvYZre8t6MZt
C9SaErf8RJtk33gOt79GUWgbK5djF4FYoDQMM/BMIud30BQHxmghzSEfIHO2r6c4
WGpFhGCKuTDS3JowGJG50GaQN1Wt1hLtWi3tBmO1e3Gdml4WF353Zz7nefXN3X+6
0Fpv/ctA0cWTmdQhdx2VWHattrcE5++XT44FGs7ufS/XV74TQnHxIfBVI4PBkiYC
JqGkPoZ8Z1PkKbAUuyZqLj72tan7j1BhfyP1XYKhRtpe/4wjoHvYDPwWyYSiuflB
z7UKF9pmZ1CaMAV6BwTrEat5GtKWiXUP3ueSYsgiQBrFT6bHxLZBivvyU79pXmSA
2bqoYJX/FAUKm4xvOPBZYi9dY9fq0Y4hcoJ5shVNCT6jkJYEQciZI8V1YcoC+p17
VJLlzeWU2XBH7zC2O4uto8mwWUfj3ZQdQ/GmCu+whMB9qOGSzevYgt8TNCsTV3AP
sByBLni9y3DMpsVOUfbN9jbfZy/OC8cKuBEJyTMi5m5n6wVZUqShuVXtrt0ztHao
UFMNHA8W58b9OUEVLxYTR9VaLZIw5t2Pk9DXYFu9RFXlRxrrXcSFzxezJ+HtJc3q
gkd6aL2pLsrV2ySPYU06x5uv71C1DCr21lZYCax+9qMfIpRrHpKDyhLB0fNqCH6L
mDou+dtW3m4U7VIAyakl4Ef5MYiJPkh2Y0dfSGl9EAMRMdb5pVx7ni2nWzCbDP5/
EnR2+uCMHDTVvaCEVWwPT07tDxgqcT8aqEyVjEWeMIfhHzddh/bTF098REoNa6Ye
SwchffGhXcD/bJgGRGWOlTRLhYO8yKgF7C3TRaSUH8HSRekddXZ8KLdTj8mCqrT3
LxJep+/XTMiH39BVn2Om5laN37kUYLNN0EyFLEGZhuQlpeRS46b0ykArB2L0HWU/
qhspkvAaweacKbsyuMucSOtJbEF+5v8uK/O+c3W34JI533a5WOGpVlGZVk3ksXdM
Rn6lciKGjYL31ZDkmB4AKrEOUotzdBeJThEzpzA6DRxsc90eWrpvPCZ2fhF5DCml
bnKGsuJwxh7iiPBrA60cW3iQbmlCCLsWAnRRRIdt3Qdu0SuU4WH43i0jWcMIk3Jd
oE/SzurxXGN+hh3S97FG+4p3fs1Ek3dJbmR5YEiPP2qkzSI9milZwDgP2MJz0sIG
tnCQQOQWOo/Py80Sy29p5TFBFZfGDD6U0Q3XYW8/aJPRU1ItYWX6DBjJiihScTzX
Ccg1zC5wDQE6t9YSDhfpIzPp8ibagzjoGMYQZY0ZweveKEjtIPr7ddgiOHVDAtFQ
NKWdkDCu69SY7te/etvN6bpCc0HlbGhWdbHWpFdKHc3CcyBqo82rZ2+TFOLNr9jW
1J9MvLz0udEILni6BOMg7KVauJpoJs1DJTjSHOd58sMEvH+6ztKDWuH1LyWb8ZCs
zKt75bq6nrvKysDLgcSQ7CZfqAYJ5jTg1ZC7vu9/9a5XvxHEdDpb+gmvcp4AHjJU
eO4w9A3hw5AeN+0slChLB0G3Z/cQVptB4/r1mUOqhwroQgRXDLbW39BhnpzvdUR1
46Na+kSsoklnQAlPpNqIKXgb+AsH2kPJthgwrGfMPyAQAmBIF1j3V0XnVZYN1fvv
mpyizO1XFURW/2ltZJXlJVUMFQcwX9wiyCfGdJwHJJyOW0Xo1U4cQWQmVIIW7Oci
x2mF0R2aEMUz4bdLeOy/lxmS1m013C1sbwxF8oZlr03L/sgjQtYpeFB3B5NkJnsg
vjWA+SINj6Lsa/yzh7cS2M88Fy6nN0R8XzG1RvpUq6HGsXDkEnvdECPdAIf20nYe
X0PsS0Lq4XKJ3iJ2R3qziupCVlq8bQ2nyLhfnpxDC+HSgtVFzBa4PlWDXQEdpEMs
/2KDG5NZIBSZPXTVC42kPqGUvCy8oma7Ah6QzD3gIigEM/Rp8YNHpCXMiTZfreQp
S5jNSCael1px45B5kjArikglPsgd0/KGQY1zeJVHlMpUg8s5+BJJlnC5s3RQOZJq
pT/h5yVPmIa8tgDTCM5mkTvvuX7ZPMRuh1l2y+dGSn47MrXML+ks5OBm3akaEFzV
5yOt0WSHH3E7/Pn0ndoKb/i49sIc8ZnEL+rRhwOBXVWf19FTFaaIs1pe5M0znJ7x
kMzSGv4Jh4Zd+CtL6OcijjrBb45gpJuDvTrkinrCmZNnO2nU783aKXC72Ximwask
v2QrZfqZRC/2MriSQ3emf/wAu6Q6gCX4T1WbjHX9wgaFW+B8+CtRUURPSkEbmnRk
TnMDUA5HJUSKZuPMSWsNnaZdpRLvJURnfojiN/Kln/AXOtj6Sz6Z8MK7V+EKMH8m
AcnFJmiToFPzd0X8IsO1XopMVPrEYCxwaWZK//6ZnrHaTq5SJDJ39JExMTiE8Gdc
f3L5Ez7UpK7BJBDFjFlg+v9g+/wQ++V25piOzJrN1E35woL7Mh/kSwUXO4m6SYdL
t9PIlHoEgPN1ZzXkrR5QbPsAIks7emBtANJCFF/Fa5J/wa12lvozswEjvyRlWKrF
ock3fpXFqOFVj7LuEt7nKJFl+QEhapQ6K6G7G85pT1AN/vfK+0YYU+EdbNzNpKBX
8Vu3z93Cqaxo/2Um8Xh5b1kIKrxVtPg81IotYWaIztlk7KpjyuHWSXD3IrM4KZLy
POLP2O6vIbP2ItAlcFQ6JULfCyXdUXoiTqlUe3uW16H4y0zLCod+hxfuSHD7mph4
KnT6K1CSuWM9OalVoLtMqv1aSacXB8YIpal+ELvoGoXWByVPIabRIAfk155vrSZu
1GA1Bql8GyWLxm+VLZs5Io1MWLhr1LI1Ze1gfi1J8w+B95NFgYeo8HcIXTXO41ZR
PeH4IfJS/RszMDlku6EBgdmw9Bea9lVSoucMsXggiGgshviAj/5tutlE5XecOyw4
iKofAXmcyhLfS6ou8AZz2Do1E3kBbRpKgDzB23eBebvKFK7qSSzcNF6wucfbxM4i
F+u1EEcx59vtp/P1NNQ4eM1NVgUZ+btdG6g/LvUVwgiahqbzG0wcolK004UhfxYA
Mv9mRhsZxaPdk37hzMuS47dFgNh4peqA6iUvrW6PTfhx4puivm49GBhf2UN1va2q
QPxT+I003Qb0XWBtYsftXwyHPX+4flu9+6xv+1j+KiADVuGMvdmAZyjUxlIL5aa5
8BSnW4W/imvwUpUHSW9oHRsac/PEjytP0KlorAMvl/hW3iOdEAKnze4VxRgIuEGR
uVTCZtnGjmStu8T+d08np88q9Afks/DFeR6J+OknFEHe3eWmp9fvEnHdvTnqSuOX
cr9lut8Ex0zdhvanMYHPqBvfUTEdzhJYd/q555er/ihp7d5Tvg9gFI/1g5TKbhg9
pqI9loazNqj6B46KcqJHNm2VfHz1C+P4GQWBcpyB0a7C65mCuwSn+hUGeX2e4qUP
SjYRG/Azh+RqFl67EY/topZ76JgSka+0WYulCTsqHwOIpLOLGqimbsauXTlWoP3s
TQIkX0GprSWOq70yOjYZ9QdbO9pikjO/kUmhSg9mp3myCKC7iZVJ8RulRRSbXd9t
Dxu+xb2Bg6svSO5V8wQRqgygV/tnfSoNJtdCuDXMZ9A0XR0aI5JXT5as7KZoW5yz
vQWR2jMaHoI+yoZz6GuIbjuy6LkuUF1MUCf6tUli4YYcWo8dbVdzJuxU4zkd6Aor
UMzs53biqg2PIl0F5+EBtMiST1o0iXrJxRFoCCbQiymURAC6YjiVWJ58GgBs9tgz
oNu5tXsIaSEQdpy3sXR3B7HKkCSFfNtPCJC6SY2nrGt082NkO8MOUj5bs2OpE+AH
5ZMmd53hDgisc4PqRQ90j/CRMb3Hv11Wfi7iIOyMcVQqJjSi/QXJTwO6H+xs9xpA
qXAgaUfowGRjgdg3lfSWJnOW6qeMiaTUWgQQBju6X435Hz4ui+gYl9mMbtuBWnJH
oXnLCMj2LWciGlVGV/8SIC8NBmH/z3sqKGzv5UDJCjF2USG33ucQMeYfKLw0QPoG
SEtw4XQ4MxUaJ98/mdh8r443s9lHKgi8BvWhpzPaqrEi2e5YFcQxEm0KkWvFlMcO
83kqgOho82TeoN2orBkGD1Arlk6GH1BU1FKH38luZV0bpFR2cZ5yUUzQhbJTHFkJ
pF24GFxPjceUC/Dif2honx3QRo2jfnUXWLgfxLfvI9hiF7vfMZCuLONjPmGqWvF4
63SRaOFXq3TtUsJXFmBuCbhM6vcjnVeYg+MnEI21dmyiWxU7IjnoXtVkY9ACrBKk
aiTgzExrufG9z0XusB3ktiewBKL1h9cu+tLMp0sAsZ+XY2nG0wtelzG+1mXhb2tc
NZIbAoJw+11fHxB8hYLX/xbkziNdZ8LZyaMuxPOEQx15q+kFkx2EJLduSGFv95Wn
uZnsPn7C6MSWrJM84nOBMGkuEN8CIDqBMsIA883Detgc8meVTJDy08nB/ooDHhSd
KJEPQBGKkwp73B7gIhOb8etlR9c+PAW5gVM48ywEP4FrRJnISQJLwV4HNTD7VZOF
SehDGdlU+jhA5qfbBO1aS3AUoLFxygSbbDJr27pcSjiirqTbyE3uM60LthjSAzrL
7ubJvAXvz8p49g/fcVHGUxQrQ6W09JqCxpIRza4e8cUb7rPpfMJXgyCa+N4EWlOs
EefqDEmGzXJTC67fP/rbKus5ELckG43rgTotAl8kQ9V5GGkeIzT799blcnLsaUDq
sM+1sI4nLRNe37Enqb6boC34Zs2GXc65Tpkpo6YKARRKTKz+9L4QOJddXP1i/Kk/
63/qcp350AXsNFPO8s82FLtDBS2OJdeon10KOiwhDhFRvv/JDcaWgXC2NehbOTZW
3E2ic8Z2A2Z/n1rS55M5lvNW9GV5GzsyWe4aUThCn7OK6XK2jGw5td65lcszAC4T
HbSo2r8WQzRn4j1CF1PKpAEltukezUIXG5qf1qjHt97P0evUW8so36JZ6rvRrXWG
qjlXBn3kPbdGpNeBWWfykcqbv6quFf+JI3ySHbB5EDt6vNDqIWWl1VQQavH6Pvec
oy/riWAHSgVUopepbF4j2MDQO9nWh9EeXd653aOLu1ELAFX6kFNhT2zuL31fodyJ
Nj0HcGmo0BqPyLfQUzXuwdwV5hjZEkCfMkJpC0vhgMVnknwSvIZuk0nWH/1DbBDJ
dRn485w6wNMY5wsRaxLwDE1xr7lQEJUXd2s/FZqPaRLX0Lal/vMPSwiO2ROZU4Rv
jMO+MDa28ebyCiKBkmCJJGrwDH/GUV2fsWD3oQZQnu9PoehPNTeXa/UFS5eqwwja
FT5flebSOWgqPC1ORKR1zWGy2fjjiIgv9ylq/LYtaTSwREVaZFwDUppu1DnvGrDz
ddeGiFAcSfKtS0dWVAZiQzaZM6GEonoQqDaRJ8l5E9G40aLRnBvcvuP941H4e2Cp
ocjCzwQK3um0Y0kFh2wyap/LckvD3WETYqqXSOJ+vfF04AXVLKuSBtebVdSXLYsJ
jyHxa4z5Z71DvVXyYj4WWAFdQmVFg7s9SNFWjGeqfGUzBw1YGGwp0g+x0huU9gxa
JLzICAW947aCUfDyESyT2Bq6k/pNvXSVldjjj+I076B/oK4ALlM/ge7DWq4TeBjL
o9CNCEgTCpvxUFC9/y90TnVQ7Av6Mp6jKUzZhH95iDwjTQGXf9ZO9uBs8xVrKwrX
jLZinkin3pZ2zKEtETvqZZGSgODzewJ1fdhhWisLYCenqAzFMeCPiiBOMoBAUQ7u
FKaI+QZIoHruNXDsZK4KfMkm02l6v/D61tCpxRA27IpSESrwX3taED7oIzSdeFiV
B9ryqW3GPx2TxE59MkD6E+9nquQMAuoBXC06p8gJgOAMLqx3gaqREZftS/Xc42hA
7c4QC9b/NLK0ExPHj0Ny2HPeQptKXMWDZm7qBWsiU+rJanPQlQHbkiWKliiowI6j
SE5LFn8+UNgl1r9yd8PzBWUiCYmFhMIh/KNFfI5CBF7bWT5XK+wTWcCocdWBSooK
jRLkE3C36hTW4tAJHp/lT98eNbpNhITVszxO/J/hpWzUtI6wZjUoRirYopsxD06n
JQiVneyorIr8x5WrATNlS8ExyU4jBxulj6ZzCtCdZwyMDbc+p0bsgRwvdf2jgjcF
UYstJ0QrxINGPCzmGfrcR0sDjMPu7O9xIS/KxaSp4X8PLYfTDv/kQmRZ1e5GTluU
kDS/4zessGXFndb+dUeHagLTvwGWyMAlR4bZhO/e7Spzlh6szFYUbwD0cOJWYLIW
5Ux8BXY//2ieO2xtAAGCWQF9m9/w8gkT4khn56JbvUm/GZuQ5byCBHfV2SfiPI1O
Cp/KrALKLWEzDMvvRs4e8MoiKfeb+dxFKgq7dfnRKUQVdb8GOupnEDTVDesqnjBk
tTJGYJWNDzHNiZIn5rS/aFbx8B1PQeI6h2SsxsOfmwxs+2k8WCHEIfkF4mCtXFFS
A+Fkwtz0ZS2vxnQ9AeuHqSj5NLIOtp/XYAigaRR65Rg+h1jg458gJKepmjF4Gz4c
TGnkWdO0mdLGadLL9LGPZsTwL9AOsFH+Zp9dGvLzZ+e0GrawvKMPo4gDD+i9T4wr
FwIu+j4JYRV9LLhQhObWqCpOdXc9UDJkAj5alG/J9hY7WrfCx3c6IBm6uYJrgPVG
cA2BmLi/gZv1vabZjpGydyA5xq+O0qs0KzDpuHl29bot0GNVHtZ+BfBup0M+s7Tb
bUMGn+eAA7xzTa1ktdjIHEdPvivMBPjmZMpIgk7lMXAGJCauoHgvN9lVAAJ7Q8ii
l13Nn5IItP9jcwuzjezaoZFA91QgVI7ToBkY1WuQWjLzNHOaFLpm72OOIIUaxk+d
ZRGoHije7TZObdf2hLqMaLSlsUdjSGPSe70krLgMPqDtSmEoP9KA7GPS5tgxKv/X
lb/z3ee4od75j2Qe76SKXR216cqtH1V9eZfGNOYpDTgvr0twXJzplgLS4/CQaXKA
5ojOH6WgyLOBPDfGN4bfXnCiYMqWrL+YTroiaMe6RC/PHDqavig13DAeQwEwgWbD
cD9LlcQSoFEQNLa9y1VBuOUMJiPG1z33s8O++b9YJumEtmTDL12OiQqzuAu9i9Ft
x/dVKjVhwWGUdpfzD13UWYho8a0FTuo/wEOC6UoMHTRzTfZqDZgwuO9VnrFxRhS/
dmAuMAt2TW54TH7nEDug6PkyDdaWX8wCTBg7AerlrWiG2Mcb3M9EiDgNpuOMHMXC
5Om4DtRDUIuBeyFS2Lv+gF83i6rBsbvnOdQNYW9jKGyuEpfICd24tysq6j/2nWJg
zeLf9ShyyS8tFQxed1a7WO4m0U1n9vfMcu1RMNWbreCeCUJt47gOQ3hkvZ16FaUi
NKTjVIt7N6LfDycaZ5bl4HEHzTs3Kj77t19l5ftP0yJmdhL3EQKERn5i3gFt9PYN
CQj5rbycnhJWgD01xG3yi4/BOhNNbVksDGprBb381alMeorYZ3sYIzOpDnu+gA7Q
zMPD5dPAV0LxJpmFKkihrpW9HzGszZflVWJXV3CsteaislbZFuQlyArETnPdrTNK
/tXLwKCAcpHBvm2aYgDSn8S5HenibqzGKgmGRczgEZfpAWe37YsFfsw4ZZ6NlAzs
j+xTixQoUr9//amEd0ZXee67kbDm9ca5Oe5XaXrlcfRkxv9UR3RLRRA1fdA2uCTe
tGNV5DVT7+YgpnFpTuuLeAFLcQMXr/hLWl97uMbzvkYnGIBzUU6kPRSacKKZUOnp
li2HSnt4l4hrToZhYM09els+zr4cgviI7LCD00yIb3u3PQyV6ASHA8yK+GokqeUC
1xV3FRaaWCMMIn4XjbAIbr1NgIVW4m3FnyF8IJulr8sdxunwIxdfdf5xaslIQmcq
0AlclY2OP/05+7PlzoVMh5FBM2e5jVUeXr1q95n1F9L9m08Kl7/huBaOeB+1G2AC
JkVdAMfmQgtralQgM9FaRhwbjQRZLzfWBy1Kp/i8e9Aikaz65hEmnk3EiMaHjlcu
UaftP7bpy58EwPxLsgVGk/BQt0xmR6ZIL5oGurnL7gBq9PMQsX54TVhfjcDXPj0b
Ep9K+u/lSSrUrb0mLE4SoSqU9mb4NUhhDLzVvd5HK2Zk+PjviR6+FoDWZZfmZDMU
Jyq63aHp8qxdrv+o8khfynNg+quK0Cn984thoO55ohOOcT3+/DtMcjyxxtyJiP6w
WF01W1sUmSPa6YmnFIwNZgDvJ9Wzpj4WT74s+sORPBL9w8UmDgR7EkXSjc9z/7ZI
4V8qMMSqyzSWZNHJjC91D+gTuB/cYDA5jUNrMNy6xFYDKA+xXiUpr8VlS0GN70O3
VO1vXE9BXjVCYiV2chAyyeBM2vlvJmbbk2rpN8nfYkQEmzNwOMmpYe4gL10y9/Lk
o78rBpoFZJCxI2anMfWZbK+wmhyDHRb6YY/NrhCHIn9TFgQX+LWONKplee3zNw2K
tKR/fC3k++xCZBwr/aE+mcoftOpGuM+hopqN44RcAx8qQ5Y8OXxrszNibkJ7Nnd3
t5xBPuavMVctZii1PbZOTdIWnTzihOpNuowN3bt4Qn3e7VrjzhEkQ5aZ6v+Zj2ze
gOC45rc9rfjt93Wmx04mIKfEHIorU2YDDA0PrjyWGUXCyqx83fDQ9PiD+Uj/N6UG
Q61ZOi2kPhkpCOMIdvZCWnD8vVJjSLfKMqezOMkJo9NKzuxLFTPzFl2aAi286osO
TESRZo35nouqtA5uMp1h04c/QK7gbfivC9kuEIp1iHf/FR3a3XhL2L71oLKhD/cr
S6Esu0Nz46u69gw4LjGxF+VWG8Bb4505x7Jk04hUySNiTMpVr5C0DGmQoXi73NDV
wTr+r6bL0I5erT6nBT2/uMGLL76O+QlWVZ7pC5cVmNGMzR3+W8+Op5OAc7tQoYZV
fdHuIXBsrfUU+fels+JBSdY4NkDUOBa3WpCuUOHqSF90uEeS0+GFJ7MisSyy6q05
D/bRI4+/pmHP9D04XdlgeNgn4+lg0S31XzE/pmaCKwxAGgzDmAPe0iN8hbLanZho
uAjDd2Pv9LlN6GASDp70hjN4EsvP1RatL4mcIaN3rSDaDOit3WtYOMhmcHjOtBep
/GRsgK1UlqXKCN4nrvVD+FeDwIRppuXudGDa7fzoTT8nrKY4pOmuriu32hewAOXt
jjr8cFi8pSZcjT0gvz0Xwv1CyE7+IoctQD8SCy7+BkbxIeXBo1WUPqzDwu/6gg7F
KJw5CafxsZKxIqoja1RDoOowNtNOslTWWEbgNT858Fzlp+lFt8pDzNDImL0GrITn
rqHInCN5Aap0bYKnq5imEpnwK0OruA2niRofb5gjHNuo7yKurvqtOJBZ7dZH/HU3
zQejcVZDdglCKfrhPXiI1vgWRgGSSOTeq7Ilh4c0Bj0OX/bga3ps2x7MIlCTT82f
AxarVudjmqvClyuGEELwApdr+MJY3tlGvBwbXAJ7b8eH6I5RVPjplzbJlzKCd40C
VwkzFaTT6Nu5Ad9dVljZUygFPG8gzlQHm03SFuCctJcF4qfw4vKEZWrI1j+/1GSA
S4x3/OE2oAwZTyXOhd66v4+pOsK2kHHSKwOBDYcWqR3+LOcOXgR/2DnXWwB+DbkZ
rdWTX7v/n6zhS/Fpnr7K335u9yWBB3e5ZYzqGjIce0tfCkXylCNxYM8KKxD/ThSK
dybdMAjbHrh/VlpyTCdJN+0FVQeDz91QC6FfFivi7wgvHJAKoAE3YGImw/Zove8L
bkpaQKstVhGLZ0S3EGEVPCmaZB/APUctK8xv5b0qzvvnqA+TL9gJg/f+yZYpF6/Q
l7qaFrz9uJAkvLK6tuz/0ko5jPQLUssmVTbttkSIeGohAEX+NATuW/mdAbYVuCAV
zVplpOs6AL6UydsuYrt1JoGgdAFIoMzvbBoHLZaS0mu6I3o6atu3jdqw2m7f+bLR
WELBDcRZE+BBK4+O7f9PwsJwozcak1Im5alGS1VsIfZ5BNboigG0qWVR/s+WLU4R
zAAVgr5EDIU8uXLI2tYHXT58cXm9Tf2WpAsogGjFQzczSASGA5sBQtCJMtyurdcD
XaWvDGrU5v799hYHLwj+2E0avAYXBZFMlIKZuv6aCo1AMKssgB05CXLmqSfrTLMb
ApHE7vK7tBLVfDv4JouFnPUsGsgfbU4AhdVf6/L3mJ4qDgrMM++69TOyjryAAQZk
hcQFxaxUPGPVWRJROn5fOL0HbC01g1KfjQ9FON4Dc0NI5jY97zYVPtGcKlLFttHu
jOhG7zLHTRcw6gehg6i+E32ueMLAm7KXJB5tmOjje9+nLSqrhKktDCZdRD84ZuiI
Uv6rhi3aPO7qO7+VDMcF5ZztGtMeS6qkgzsB2J3PO7aILsASD1QNV9rQ826+mv5k
jkxuFWQwYkMXFXYyK57Xp/XKJYctBUaSmSvI3F1gCD1+IsclEYqAEhEn1gs09x28
9NVQBd0U/qf2CZYhHHrAxKgClISOM3FbggUkBkCnJPaLAjqGlqojZFRYv9yCV48I
YkXmBj1d1TYLAst80r6IUHOJux0X555Cj6XGAwamrj3Ar3VFYDez70ntXodeWpT9
5WFkdofHgkwrD0/j1s2NcMU7AYyg2W2Z9DhWg1TF6l9eM+cW3VovhTYVGgLWvGOC
nJskb1RyBKptieqsGTZ4D4brRwcfwTQuXQFeVfcbG0GdY81LTNYWiMr0GJJuyEM0
QlX5JP7PJXa4rBcVkgvv2eYlL+oOGIs4KZWCkWZ8utNfm17qL0WSruHjE8JVkg8a
cevZeLuEg2211htfNQLyVo6rWttaCrFUItbgJ9ms+2GCucm96ohsgZmYI1LhPzd3
wJ/QrEhUmZDGkWwUuo7C0NZ3WMZ+A3ozUR/yOu0JSyk1XOWSAllcbqykCpArr3IZ
XP6qH8FERbLRP++LS9DkUqtZvUwoCgeLq3YkUiKzm4qFSxN/sUgWPzAteRVY062d
1Jv7PFYk9Le3nbztdFtWwcII4zVD/c8nBkHf2uDM3iQCe2K6UpHup6V4fFHL0KK9
7KR952a9Cvktp792sSSpINlCUTRNDSSeUKgFlK5HWKQUlQyACeuYscpd1w/bEa8i
tyP+KgOM3MaCmUkwILQrHKmnfUPw5KwB0PjyEoqyfWI5hMxsOuQBAfbJswCeOOMg
1Tix/q/7evbDiIptUWL/vsKvConDHGJRcOHZ6qhnwE6uiL3K93uK0hMOw5TMcXYz
Z9ZasEBPZg4q5TQ14RLO8yyd3EhcXaaIo/H/caZUhVmWxIdipkP25ua3KKBLbWww
ys6qUhmiTX9nm4JWh7EpGgvSFqKu/EvuzRrC4ZiDaEmxHTjRE7RlTbiqEuC3jSmj
VbHzQ8P0YSFdGffZwu6QBMySUsOWLCH5+FhEBL8v830cXk19eoUiNZLaee0qt913
i0WUJ0BX4l90x6BF0XqHbpm60OIODrhL16TthWiP/en0iWsM/xksMdu5CmcQgxUy
LD7ul7fW9ni+7IEfxkJ/rnYW6wNYd73kRrc78dzoeLt6Ld8S5VNl6bpbFOcaYNvy
8nfvvZdpKOc+4qfPiYuuIQ0BfPSBOprvPwoIWtBtKYLn6nN5cf3UyzmhsjM0MiDn
lhg5TbRFXnFVrM9sBR2iknPr/6pphYN3VvGI0yGb8IcionbVd9irU4h6JmJLmS73
1viX+vyCGEEYHA4vwp0OmN5hlFK6d3308I2XG3cFxek3H2Q8IGqryjBj/1holD5o
ixPAdwN+SJdb20dWJv8FD67T5GHbR9qLDd0razcpoUI/uV5lcMmSOqIgEJ4CHuDz
ljlWE4PjfJRtu4ua0kX/SD5qV5ObsDfjf5izAgv1CpN0oorhrnBzQNQ5bp//aFpP
kld0jV9HObzURnqx3y5NwRO7zjzmrfSzTngmrHg56Yc2fWDq5EyTLrPsHBVuxE2j
VG1q1fLVxOIGZE6qPoMJ3wa7Be5pZNXJ3eeRGk44Mlmwf51vlPH1eHC+G4Sl9W3o
HO1ee/do4nvdivGDaPCs7/If5VbwVnpuYrOy87HD6DyXMWhkPNT58Wdspr4hA0x0
rx5zLcqD0YlBzU1bFev6iJHSInDFzUXSfQJ6NF7P9uPlnAwEQmA6ZqiNUvEx1r7o
2s5Grh0Ni3rvl2jLA3qgIkK0SntXALy2uIgTBFHDVnwpY7FNLpdEkgYvb7tsHp7j
5ZR7Ve4fZznb1vrRzDWC0hBYcTtBjYpDu9Psoeo8n4xMyfzVslDVkL/kXzhpnr6b
EW4jXu6gnuRtNyGjvQQCItUn/ouCvoOzplkiJbV15S3S6y/iLz52lNtr/SQxHfxl
O8leXe88EECqDiM2RFRWMv+BOQ0Yv8y1VjbPA6bex4XD9TSwRDr9NDR4xnkmTTR8
1kaqkSYeCwfvc2kvugdnLwzmIQUZ8Ca/GvsbyYATFHFXyosxWjlU/pHnqWIgL8fs
BfFY8uM6wcHyJ3vjBlmZr8W2QAdfppJggxQgnI3PbZ6Mzp9DbcnxM3X3QR4q+Tzp
wZ+3uv90dAFKCE0Ajq/iwLYSV3JsIWlBScjzJuTtBIzB8gVjWq8q5Sc0bj50Yy+f
mRHNhw/edy5tCUWngdVMZkygpTWNmGfr89OxrRHYnN0BTUUiRX8F/SoOKLaHL0Cj
rs74vzsDtRLn427OM9KpmhtKDq/3X/l7ULqIXs6tgYux5cg/qVsTQeL/cldFNUuW
59EUIiF70ZOYNZUscs6EYsEvoSvKOhn+N9KnwHNyZ8Mfl/hTcXXJuGzj+Mpk1POQ
n0DlkBMkMUmr7uWFyWkaWgW94Z5KeXmoWyv6FDn1gI5pEGvDMQr38Tj2N0U6kuIs
Grt7kIocFNjAMHu0d3Skqp9Oip2x+KzyMJVZRsD/3wJD4Qk/yDA/DATJE5Blensp
S77d9/KKhuWjEH2EkXhK1LmtzCZ6aOQNnYFR+/GFqQDzHqSx09HGIZ6zPGj0le5f
6il6/D5HD8UONaO9b8pBWlNil85cXFpS6Y55cVFUPbpVOJ96nQR7MLZ9LjwCYGkY
gbNzvBzpkUvHHHc1Co+zQLOPhxn/Ap9VCF+L/J5+rILMeZxX7rKYKPjsm1PKETDC
S3TiLtlRd1m0lShK+p1F4xBJqRFdQgi+WEx8YilVBWTdB7OXLSOim9V2TX2lilSz
yD5ABERANhf208ZNlMdvbHxLmpJGO4z1C7+zMKal+CwedC6dpWK+jgFlvZYEmpGv
wNNWA1pVKiZAiMPM7ceXJJxahjQKJGWEGw789XKccWfBPZoVfn+6ACg1FJvJ0KgH
WgySAWNGOdGSvKMVDOgxGZaaAkD74gehyDl9oIzeLWYaoD4oZIS/OrUbwgd7j2yD
+wrmsXxmf9dpmhZrmdHjkLJmy7zCvd8QnDjWvmersLKbbj5lxe/GlZg/pXRRc2F6
w/pSUyXmG+MZjbpGaE8/wopDrKnLdhhUD7IU6zoQ1zwVpUbDXC3dKsupwBYIbKRz
pmo66PZyZBwXdj2lO/hoMiY8n/XRKt7jye+scf1UYIkqIDBtgy8frYbF72kNJfL4
dXK/Dr6jp25qYqAVhZ7jhr0jQ1RDLfkYIUFutVDw3BkJSX81ubcHg85jd19UOW2g
NZRIdplaH3iXicjbxmgyUxs/5dgSvjItTe4WpULSoJRrQVWZbgmHSMWHlnq7uV7e
O9MD4Ez4fTCl/eLqf6U37kgz+nyOFI9FTGP1jfYwq+l/sDfKRhQnroC8jTPq+uhG
ZeL3vdRQSvDv7ZYPDrtW9Zw4Ad0gTXKqpKKrm/YcM+4yiq77qdQ0EkADcDUpQydf
Zxw2h03uGqZk+PgiJEVP4yRW9hFazLE3TpF/LBF50aPChOxJgXgFFaj8hGoDAcJF
VvnQq7vkzhyYDOoMDThcMVCqIHSnV60y/RO84spVVhmoNon+jwhPvwxceH8bkDnV
UA6c65DtfTznbatTPjt/nXO6LOcXq81RiCAiLUbqpaMJtlp6PtXcvWIPijLHhVld
X/ZXvwlkF2K14ZuBQfIqlYlYRtpzUEmJGc8JEryAUgC2YQZSx98HZJjucYoI3yo2
oK9GAOOzqcFj5SNhrd6Xi4sTmodHtow044G+5uGk1BaCegWWWt0epyFedIz68e+m
ZgRnfHg5+wYgFOkBAO7xvZKmFb1LccFpRMqHytu1Oo9PZ07SQZx4qX1ICHoWL4G4
sVwBs0IQsfumlLmHGRIWXYJiOiERejv0CyVLVBtle1eHSAgkAVc/5pj55CD1BVRj
8OKvIrecmXaC57hxB5lkQYEnBdypDPAm+RMqeb85G/WcFp1YPrCsY+9pytI/6/Yq
kETJxfqp7su4TsK3MWUZm1NCQ/DGB1DU0yXmr7+g8oIySYnEHYttaOGGhdW7FiBb
KzsSzz4+tHJN+OtGiLQs99pRzCwBEjc43kZWnigAjT/Nfbc80FjH2zWVy6Qm7es6
pccmawUgpidW3rqV105+DsHvSkIMU7DRxboj2GgX/1f+thG4szSEVnIZz3LNKiRo
3EXIzxutXAL4GUWub/4i60HRm0ZNx9q5xfNonbPCpbIUTD852OhrfTVOAuQaMwnf
vJKmnpo1fVijjK7y+JianEzNoUiKiYbmPUoN0b83xmBqdVHcA56U1iOq+kCyZZoH
E6wAYeVSMa7kNiJP3RkgnXqoXBxCvE1YF9YCeAuUYMPTar4AxN/yXhiHuerCMkFk
k+YU3woMAwOyzhyvVmc7QPwy+82sd1nimQAhTCrZoeZc+uhvghLGHH5QqaW6/dXf
Jal0B5nL+K9j31lKGaIdWkxNh+p8HErmqd195yXtkPlmun9akA89eH7fO0ovqrB4
Ej2+PayM4mkLQQZ1WntR8Y7oM+DvjNDhlCXjuOtHP/lZWDuFZOoIstMQ86qSAXBT
N3OdOkJ2Z1Ur/CKVCa101bc7kfupnp1397qVPwzIDsSGZQXGYJNZzHHV0G939R25
S2T4p/KWUQwgrOS+IOUD1DTnhfIcwkCxvzgsE1wU3coIr/NCOTfTB4YzU6zZaRTJ
Lxle/ZziE8zDHCS6nxMu1pP8kCSSrQWlywAeIQugPX6RXTebQhJqarRA8jvbmUkt
ggYgsskC0BWNyeQO8juWIUcQDbXEx8knF1IQ4wcK1UGeM7BGbspGID/bY5KfEpvk
V/EOFx/V+4DB0z7zp30kIh0o7DMLRzBHfb/72Ij+ERq2efINwCkWJhIFnX03+P4h
Y9lfiANd6+tuB8zQdVKo6H49uwHQS8ZFNGNHr0ilb9OdLRjC9cRRz7oxGvLEtgye
b0i2mP8y6VUk6toDgZEMolfHvf9rL1BVKivVEAK2EmcfSnLl067tdtR5vw6/o0e7
Wp2T1fMEC2vFifxUHjxsYipKannyI3IH8+y/Yk6ghkEbIiHNetCRsmCoXcq0S8NL
kuVkwZ2PfA7A/lxkxaXdEimoA/r6JQgxAI0680GxHYdeoTdBAYGbYJNJMZOmmLb2
1L3ePSkOQU7vllVGX1ErSwtCLbattoyzshVMzxHe6y+eGaPyampTZj0Grfbfj8mb
QHJNbdF9otlsDmY6jvTVuxvfKEV9ijECZwTkEv6F5m2rjNbuojejEmnga/4wSIE9
QUxnBwjWQieHAs2R5m3bAoQHRp63UYvjZWks1sVaxorNyNQBJUE+6jgtqsOeFVpd
v/WBGKWOnYVMUNm+WfWEU2iWjVvXeLS2fAlXmGUZHhIQP0JQLgTLyYu5O+4CHxnQ
pBGfffuIDzpfAzcNuytLit/pegyXVvY5jXSW4nkvtyH75htl19vZydUYHvbYD+7E
X+zVODq1ycdkNb+HHHhRTyds9v3H+gOKEAU3PCSnrJg6JI9p3nEDyOvkvtel8yuC
/XP9hQS7uCTi9uLpngeCgQZ+iWq2G7/APmFlUWe3KfmozDM41EcU63SJDV7kjAC5
Zp8SDSg/8gsH/d6WG05AzVLj428gHAb6mEsRCS3H8tTfMv/nO3H0o7x6/MR+IT/o
uNe9Co5kBz8wDYmFMLFqJnS/FZUJuIH25JFSyicqJO1xDWWb475DYjHiZVmHTd4q
luE2IDycGDKU0MzKwP4Mg241WuomzJkFdb1kXZplCfmbB3xQQMrWvI2F85/1GH2+
ERoqLjc2Pw1pRomCpI+sONsWdUXMvXqnpNoZo0g8G0MhV1M7quVzEtcqJdYWuk6N
VxHA0RMPeF4wZG0hLpz6Y/xDJQTRjiEBYva+wrFRsWWmjA4OAx87JpCGiWsopxqC
eKu9rzCSvnwn/yNRdMXXCfI6Weh/IRzFNsq7iw1R0/SnFRe+5QqYVbBEuWP4Piz5
qNgAEnw3HaakelJioPFfWiC0loGw0vGKm+Gsoti8K/Yu9VozaGfM8G0NdXaeX7v/
PyAQloizGGE4U9HWqG283TEPLbHDWxBeneIQIZtixfPD3TRMlFX94VRLfjanwYRl
d/Ac17HO5RR38+bTpefx/up/gPjiicN1zcPByxWyr6kPfsScZlDxn8p4gmouV8/g
UmZ5w5GxXxv5pS7Qcc6h0Z2JD52OiMzJq7LV2dD+gH7Em+w4iJ54symeIF3Vw6B3
Hh0wnn+xvXOwsAIFaloLgkCU1N2+D6upke3bUBemjwH+bJ7WrBkdhplZeq8Oj6kx
AGFkU+YyowbItFSWtlwvBTQ6uxCz8D8K6aP5YFE1OuqKIHMmrJB6tjcz6plgcWAM
q6MbQkXxuipnEYiRDucxTi7n5XuzgszVSGi8Yr2kFIJ1wKaoE/JureIeWQcbtzxY
lUbpEGMnb/GkN3t3PuRuXuCtsGWHTbMBu5CI7q1sLWbo5L+qupkD8RscyYicvZJL
2ad69CKFHNsh7wRJMQMSY0eOtivw2KXZOxzzGh7aU7ZJpk0Sz0pftz4911sCSQ8x
ih/caqo5+IUdDzjFaRIaYYYILiFBKquDCOmWpoS/3vo+5fn9N/sqK3/+0+tNcggs
e3QeGlpFTsiZhCWf3tkm1JIl2fyqSjog3ylueaRi/zKZKem5eeOlbGQDClNShVx8
X7cyiIj52WLbJeJiRYhY8lmc58+Sv/l4weyeCUpZX2AbxO6PpLX9MkdmWy5BX0tr
maIkZ5zaon9RhnpZE2wO7C5jjcKFuAwaV2VWNJUY49O6GfEM2/EK67RYTTlie29Q
YjmF9Qd6ftYz7TOkexzlUy3zUuNF6mRzhBKfh4EJ0ScK07B+4SLlF7OACSpE2ieI
uYo/15e1pMUd8MLvHDcO4m0V3YOc00+p8W4FW6aH3riuEZd58FYj+idpbLdpSAOv
spX+c5qExnu0INs1XMrvSuspyEqTFvd98uCalccJ9ic3/1N3njDdMQICI8lH2Y0e
addU1kazivYWhfNtx/m8xwwwqivDeMbN4WRjvZrJ20jNtEhS0/kuefZRXY7nMOzs
UF9AaGOvnKadICwlo2r0K1Wb2qX0ay+ULIijp/NigIxdUQ9MOHjB+ZSdgkj1TURC
kR9A10YOdDJGSk0l4WJ1E9IKnT0MI+QzULJ7GKmiFElorh/KpM8viwXzn/ijK6H1
5VYoogBRCORyM8vCiJyEBECW7tZNN+1C/c5A2BIC4yEZKJ7fgldiFv0jSSsnU6wQ
ZyvQHkbYzMyXTlwnztrMS5VCb4+9RaNT8/iADdWEIRln2tqTA/gSASDrdZjyywPp
wniMp/V5REMfKfl7gPXuPP3szFtYCQZ9HGIGsEVu6C7wa7OKsk6WazGxIoSV3wb2
d037ZKTTcxSKga69Dq0w5RKTf2CKgBor0NnYZOzp6P8rlU/DuQ2zIadenclILY1W
WDoUpKXWN1pcOlmC1InQUxrPyN8GNcRyAVJe+YUZFUKosTmq1RPz2XEafdaqaXJ+
JW3oBJz2GagzpZaEXp+lASRobnFp/yDFWohFrCjNpat0FIGiHEgaYfZOR9X6YCET
UC8tkyk2HAgenaSbu4QhLIjajvvNGyP2AN7IM52T5J0NlwZgM3Zi+lgGs6iohZ54
3yFrEW3oC/2uT9jiCtbM0Czwwd2bc0J4uq6Djkep57C1Hk0uYmpnKq34FudW1yD0
xhDPdnRDvw8hxZhZsK1OK1C9g3V8nPsqIvmVUI4k/zjlEuX4T6UVvBtLHDbmFbUN
aUPOIUSMZawEDrOFSC5+EgaALC4lWDalT6Uirh+Zqx6jx7AohGbVc39wQmuKwLYA
WZYwU0nqd6N2XM4OvEBoc0xi5xqogTaOhQcAvIhLOBeKnNOyEXjoVL4TKOaG141A
BAaIAuOvawUofN2SCbvxfQXunldh1kUq925TRdPzZLcKx/2VBEEhFnTGtW2Xwhoz
YI0l8QDJlPPVVWkeL1QGrknpryFnQV8UnMHZhdI6ofrcVXmVZYNYNxj1N9wdEb90
v5d7bWDKtqcZQ4TSaRg/okezXvwmGAnR3LXFiU/ezfuElWu8vunkzmZ0IVypG4wH
lrIRueaW1FUDlBGx0QiRvjXA+QH4mxT97S6W/ub2HLx4ZSK3HGtmulyLVn41ke+5
t3gufW2pPD6TPbChJ4KA4dIhtATZfA1Q8P9mUg6aESi655eN+RReoqXMMVKZzchz
Zejpol+ltG2/zIGyVUD2MnMWQEVbxLPPNWxGkQUCL54KzQI5X8j8OUpASTVfKwsw
BBPBSquQY0IEfrHSjkPh9EjxgLHaRSe++b+V663pBhc6w8qYM5+qrF4Q5kczoXKq
o3BJ1Rs1qfJRHfN6Jd7wZtwmAWscgK3ogxdJMMDgg9vAHpt4RP/I+ttfCUTAHDPe
UlBb0vax9YYngnlyK+IPQ7azUwJLbO6IWeLKgK4z6/HRrV6nAIWcmiiwL2e8HKCS
uFTFWeSwovRSXOMfUnDnDNSLHaZ9S+Nf+/fk5xCnb/79w+OBOcHtE1NdQfoKh73A
UO+InT7Jqa4k3yE4VH803E7q/YFDP2PNRJwRf1zfvRNvQPVtDM9OYN2qOIHl26OM
oW9H7g0x7FaNpKtOUtPQEao4xCm7QarbqZviKNghhVOBA7HHCscUZfZgVBepZmyt
uqUy+n7TYvRu66ErvwE7ioSvGdTh0rP28DQf83iFethwP01S8IIo6TfGVxEcINp4
a+6xedk+Ng8jCeHliQ6vuLRCnXmvQT1iXZuou/N8ayN+sz9YXSXMjx5Uyfpjr0g8
882EEhXEPQRc5Gk+z27mf7kfETpm8IlkRA9UwYuZGY96Sgb8IA74ZoD7YpSPYQdF
SFIx3yGrz9zn6j94DwOov+/jCiSvNW3YJhx1osOaGbS7OgX+y0CoFhogVC5zCa//
Nh/03+ruSbL3M+bGGvOJ86sA35JmaTwnU+dz7MucJ6N3PiunVDRLQ7oXPG38fKY8
B/m7GKfVsaPfKtp0tVY9qdtn/wMS/nNYtx8XREU+Uu0h9zDlLV6GiajSEbRZ++8O
Ffl/ruFpBZo+1Mfnw5WEA+zmk3mBei+D1Sfdr8ppDah5u0GbSaKdvocfr5ZEWuPm
6jommLQ5J4NW72NawxVbOQMERSIllPkWtNhwp/ko9iGPdWG+98pLuGJ83/YKIrQJ
4KSoKcFG7WkzeRHSqgVtzEhUfO3jEOgZk1ePqRqqw6gTM6Aysbaj6GwZNriVPOfi
MNPR7q4EZM2VBVV/OoIt03hhRZWdaKtA2MfZ/EG8+lnBckbn2Ip9RpTlcExpCX3t
Cf/7AfiPOVaVqTOXsTOr0yoSoGOic+p5YzpPjRMewJF7ZjqlEyIQ3K+1Au3gDHn8
KFjg5nXoreOZ8hZu0AFwbz27P/rF+0P4PwiY4K4Gmn2uNpny95tO8291011uPcKk
NR8RVHdK8p6NV6jeC1jol3WbuBvQpEJsmiM42T3P81Uc/f0tp+qdtWEI98q2TYvn
8y03xjEJ5zzaW6hjIdSZh3txS2bhQYs3WoYJHOqbpeD3KXETTlQ0jZuuKRgagtOT
EijdbiZwHydz8Aoozlacrcta3518daiTgFn6FuyOBDXGqeQ+jyfogWVIxRoKVi4u
ES7pfu38nmIpFOy1avUe3NNkWwfOzuUW+yuqZoYfWSQHkt6qYYpfxsf1UYLnKwaP
lTXZG7zjCLPPbEfrW8L1wpgPF2O0NvM9uLbe/WJfGcADpEHzP3aOmUzSeumPO3Y1
A1ObEaRfXqwp3jUok74vzoOR55e0hFOLx4HojBX/UQ0Xe8nJJfNr48WTPkd5p0vX
HuWHIizIk1i3YCxmJQB8Ml01wGcyZeamnxhuownNfG6jWaAc1tQ61YxdbXX234E1
JcwCj1CrKGuuHn0VWtNOJTYZuoJImtDywm4IskScJy7xtCXnjrOcoFCniG0KnDHN
Eqe5mQUJumy6WhmkzL9H3UoP9wQtcPHI8WgwU6BFKGCKUc+123/omdr0DyMXg/nZ
flJhn+bx3ihyeSV1t+2o0oTXD2jUa7mO3+KA46iO2yBewl7Vig4E0JeJyJiOqHLj
lVUShe8IGi8mwCFAPx9KVef+XZaDYk3vmCgcQVAtWdh2gWpFouPN7UggWgmtcib5
F+8Hl9SKn3c/uvpMQYRZIZqpy7edQoQbKAhiLt7Qu1KD7ednmyuHrzGyjbCWiZXz
mwFc54ljOqbKf1vs8lt7fSrTkmBdk6PAU7b1pgIesWNyE7esGeIGXGt9hZjd4zDD
ZXcGxQvAZU3wpZ5x/k29/mhcp1uEHwrEy4Zi5fsQpESthsySmMo6IZgVAXYukL5T
MGWzUiM5vh8wVV/xr/FBugyVy05gadZaeXlGXv7zGvipq8AifFi9CDka3OJQAl9j
XeN7ON+VNESJkZi42uwrH+kzssJL2BEnir1+3Tcdb9+OG+0hnxOEOJzKzoxD4D7b
GWoPiGEXTwVEFTOK5zKNLrgB4ke7ZFKWVqmCMWF+R6vRMCCbF/pkEEun7PWRfRO6
0fJXjosdr5lEermReQdvVds73LwFDq6t/nb/qPVH9KlfaXi92LwIXd8MH1SNB4h+
IDpgKwfuukw7wardoSHYBrbe7X/NDeg3qaTl0NXru+9uVr3iBSe7lildDU76nX9p
IJnRKMjj1BCkqAKvcm8nHAYvlNZU4nxsLc6/X5Y2/58KBNzGwFmQwTn8q+bIeI54
qftzdZ/YMTpMeTTGTcg2FgU/YoyUEfbKga9fIJeQ+hMu1sYrDELnuouqanjDB38w
TF3y0loZlxPy5+NRJsmnLzHFkfG3OftSjnpNB8ry+M22xICGh5aAmQBDD4941QR2
vaLoBgmJKwqSJ4bGHIJyAXF4x6qMfw3Q9PXP7Sb1OsMB6knvwSKpT7XG3nsEhL0C
Rg108yiFXLIPkcgAyf3PueoKWoQ4OEXyqJ9t/4L1Dc+0a9G0Ze/fN86Tfs+bjiEJ
RRD5qkCbhyYxpQZ/XXpDMQ0HqFAZVx6muV68getyhTvMXHDt7HTwJq69BnvvFm1i
qS3uojrnKBO61G41qTKFlFTNsojYCBwqdy46nQBdfOhGti3vh+dMTKOFjy04s+Lj
tgzKVURkjZY9q6ymdd3Gh+WG9b743vFdmZjXPUK7CVvs7egWF2vAxysgO7X7dV/f
VWFxDc5Dq6ip9RAJOlhg+1c+wMJGjUiKNWhQBQUDik84Bk1HIuj2ZJuSgkgruroe
2Duw7MuV40iHdYwblnRNy41nAbcOaxNWWslIPjULgcNPnd4sFFj+c6lw4oXSAXra
pxd5sV1zLBRBfziSQJx7wTwk1aKVdzol09xVJuiwxlN1/cVjEnUb0kRK6vwZJS5J
GFElD6yNBMvTHAGnd4gAkRWQSmPDoUayZ2AZTQOf8FJGawMNK53VHiw5aSzN/r9A
bmR+wSNm/PlVUxUNNS8qnjearNGZRitsr2e183fw6O7xK3p+BQwMihiLGsH3Ebhv
PB8DzDEV80OLWs9+IZia0hr5fbi2kl4NYF5lCEc+kxBFbMN4xSGDpE9Kk2HEuM2H
OSAuafemOWjFH8ckrYsvsTesJGpK3gD9AzWa5pbMqwhQYxvEBXd3F0UZvYSFK4zI
Lx7ELmTlQEO2po7gabCN21PLfSC1XfKQaU5Vi2aem126/ifRuApgH0GTpZi64JHH
bhHOMjZR3t5xYSIS8cUEpYn/PY8Lfn9P7Y4duUuImZl9Z0Y784eU9P5mb4YiO67V
TguI2ZFxIa/xQZNHlZn0j3HbwVbsP1piYr6vgTFWPZj5O7DNHJxn7Zjk8VcTwNUT
6sajmnIRW7KPGq+w30EEAYtUBVwZggqb4P0Vu6OEjjiC/+gGZ4D1nymWiXZKsm2Q
zVb9cmX1L2tbPXDGiwieB+9pY0IL7/8kDrR84iXoe9MjqJIlZ6mVpS4S/wCm+gmp
Y9OXVkkNFtIn8rCWQJ6KRZBdgZmzmyGGBbYmQNz8UpTxR1GkS9FF0DFOVQ/pZJg0
edEOsz++tWkVMv3ZkuuIlosK6EmK6uEQBlYRD63gdZOSVeJkBzjbWId3ZHtrfaes
LA6m2kfMnGf66MmGr0/faSzyfJBE48PcJi78I3tWAiKsn1rDM3MLF0BVwH6e+W08
3/gR0sl4qBGg8niwUTK1nX253JY8jEP7FmU0bFPEQdhdWyIfvD61Q+ZAvBr1husA
c7QVN0yHapicIXa7bTmzD7nhQ/5xxLmpam2aXOVSJS+gv9g/ecPVInu/LoQUU6gS
0hY/7PsxzN++QxgkUgwRJFML/o/Fb8+WpmSnNZyaZVT82sx4F48+o+KJnodZT/Lr
QIYAHMHXsMmpDBiX5gziNUknWnOONsWcienjFOOql66OLggXfVz/Z+CJUrufkLP+
Gsvwd4IuIh48sNp0d1yov6ZlG3tBSR766O+iT8iUfCdfi4AMK9xzM5eOfYBhbxPv
Io633ddmFH5gdqhSm4q4EfUmybBMBbTH44/i3JQcvTwTg+XqSoV5gUiaBWCru+02
uUOq03WxLs9EAwGNQhkUVro8/+Vsgj9HnzQLWSqjn02TnEbF5AX3yboQiLXREq8G
V5o56BBwGlNNs3pOwpUqFYKz8BwSUn12BFJl/3vsYu/hD8/HnmSdr23htKTScCOc
+t3CduuulelhJjcUX/sK7rBCzb3gtOsbTeSGjFARDPZ0ZMZ/6fbC/QptJt8QbIyJ
4PW44do7Ro2KNzg+G9GwqACdklqGNIVLMj2TFZQJ6CqOlMdSs+zAUPyvnkWTqllw
PJYsCG8f7v9YyGqIJSTdgpCyUqMSZxCZsu/UFoNV1p1T3snPzyy99ecV2M62M5MN
C5W939xtDLZcSmolHSPax2nbrnhllzXoDyCwyAviKJPhvbHppxEn47NzA8vCxa7H
p0mLy+YYGou89RWKwsy9XnKLBcsoiiXQ9iZmkZ0NLae63MS/86LPFK0sI2gcCIbl
/GlwMB4+8riCCPDBvVn5dzk/pjxVwMRn6oAla0rQZlRj5XVwnz+GIjvN4vqJCGwi
zvC2be0eTwaUxc98+4yCSt7/FLRR9jNgZGv7rFCTOP3LARPmn2sfxNkg0JNc7FB5
+zP/W8UDzNpAJ4RyP0pbkxXqFnGo0IC1oApGwx52ihByUHpgzHHMIsH+BuCyBW5X
V2WbSIE/34FriQTAROMLZc+oSVsg08dJkO8BdvMd/5au4OwAL8G9t9aQxSIk8cTJ
6heQx6fYOmw1amrmoaPIphVzhmLCO70WfNEnaN6H4I66gkzamb5rGPGuZzG27GxY
a0LUi1rdoVua55Z0nxsUTpIPYV9/dG/n+g02c4Q25uMsQ/MpeDtAn2aFRMPdRiHR
jQzOFWMNcG+Gcebrnqw2ikxLyV7xBQJOud8dndIKoed9xpqVfRrZGh+FweXm8JiS
Mvy/aNaeZlaf+fvML1gEA5dBJ0mh92v6DOHAW6xexX/i19S69cgkHqXU+KTrKwkC
2WERiK8ruOGwZF6tLPzNM0pVBip5nf6hmHwdfm67EqVwU2KJ6oPhW77tm538dGEY
FqaPIQFCjymMxtSfTuyyi1oKeWqBCD4Z3hR1/Tta2vqwI02ggYkyj9ZjZmgSuAHr
v28GuPJ5RNHi+08rzLrucUcrwU1upZ7yGJOb+rY63cHLmdl+ER/7GEKUtUuGNnI4
c+kHzsM6sqLZ3yGPLlc2QMC44KzyveGgiv7VElHMGEnQAcW4LcDCmNRqQhZYqR8e
wDXSRaa3U7iZ6vv6sQUzAmfd5ZjAimgebwh7Bluhrdwl1xRvusGDf3GHMEY8pi0n
v3Ql68Sxlu0oTvAwTuy+BpZHlQvvVZXcTvv0tbl56c/VrvwZlOFMAoppB74nOKJ8
KJVxuyyYEGCA1uoMgv1Kb12tBJJJo2ibrB/tUx/5mZ7uo92x1yceJZvZS5BfvDTL
OnFomhjL4TWP5L5iAlkZV7c5b0LDq9CbgfZKPFZ1DvVduLvj5q5tBuDUPBjq1FPw
h+en6WObEQ6LiMcPJRBVwqlt54o6kFX3b6hBD9HqmV1eH0TQf1t+r/Fr+agR3WeN
zMZzGXXwq/dgbxzdeleY5lL1/gs3Yv5Bt+u7HCXMIt2lGT5GAMa9ofMahoTRjA7b
LxS7b2bb5JDkvfiIB8BSexg7tY/cVGTd1x9zaKo6wA39s2dJgDEzOFImfFN9HPJE
GTjeh3TyRqH0vH1Po8Y17nK6IBEFUBoo5hSeSEVTTuPOugE89GR7YHqKGF/kvFQ4
GkF56Z0pIHDrK2aDsJg9Umw52g4s5tCJ1SunnGeyh7U/lreAsJu63wOIIak6SvQW
woidpKmCbRK79ooasINd2C1aIzh4fMQft2iH9XKiEThsVMhGFaPiRW8uiLmfBeHT
27g0VVQqpPOiQF/Rmw6J979OCDC1QPbBA5g6Q+JEHRvyA4hqNM8w1KydTP2Hyhlu
/2wmGiSMKbsK+s7sIxp6muEVDwl2I5dfm1F+fO7EjJnCrB2j4ZmYn2yvY0j2HIRJ
2dLlb+LxSnWmE74OPh9+BgBTDd37ovAtUMJqHmhDWdH0jJnJgEqxYwzXK7zkCh2Q
8aWQg8bmmVoDplRHi3xcD902NIX/4ElQXswpKj/qUPuxIPoXIzn68yJdXPJCNrUW
iD5okv9ZRyH5blLdHo5t179V5KbPr6XzY6zlRFEDKRFMB1QmjM6JTZWSuoCk+Kg2
wwgK43ZHsscXCzicoZ5624ztmBlagNCd2B1m4gjfRVoqmly45PcEE2drzZcVCUU1
fjs7uVY4Sbb2oB2Q22GT2gMAUPxfax+FOi+dcLox34qWGeeMlMrP38cutIUiwfMM
z3sxm2CpjninJZNnGq9XF/eCVV4qd6O+nVbeBbrUZ8LkrBt79TXlkMLMld+q0vPr
huziGsSWl3X5OMorrQCwIsokkT2khSWSmPeHEryTA6q0fJ/Mvd+i90PiiNg9sXcW
Th4mRuf+4+vaNYIZ87pAWlPmJEw+mnmmEptAhF6CWZanHCC2WSF2tjXEtMy+Fsw0
9bXfa9MQP+T68i+lGcPDnrBODWwUq+jYxBEKwzbJpG31pzS4QPOHLh4asoX/V7L+
UUOy6B58r3UlhnDGjJu4gZHMuMkn51DxHkdRNxjZLcFEXA37g73vG7Rwkyr6RffX
oDch7LpjECpy7tG5PjFbpllKqDnO4dC/W211VdF6WaY5YrWOUbjyJcOl0+pnlBHr
TUCiisEUaHy+x+u+g5QQ+BjO7ZgswQgb/U5Iz4PkrJro8tGPqb5MJXwHqFniBIJM
RK/93nKO1uxwk3nd8QIJelXcdTkT2j/dSk+Xor5OXvIdGubBuQoAJd0w22b1v4OD
M2Sl5GDrn6ioNaCS4eSxGpBv1MfEiF0IHKtGq5Tk69IW1SDh6YBh+uge+mOOHuqG
WXSFYVTnHnxGcLyxMkkodK9wtC0lafhaFU72uyODYLpkU51Ny5e2hTsQNL7ub0Pa
xa3G78BBXWKODuZjDYFpLjkTF7Zq8nE3y/ztU2iwpbD285XlQiosk9hRFgQlSlXp
mpu/1T2h/4XJMsjm1TiEVgWfupedNL7OU+eK94mGpdDpmHOluGmue+hVVGONgFc0
2PzxZUpERh3RwK0n1CUaoQ0P5zy2MneEKSonxa2oomncBd8/fgKGX1fV0EY8yYK7
JFpKig/SLp+IX8uGZfbie5Z2Pqvxyv24b/CLp3WaT7Gcr47J2Ooy1xUmt9UD63p2
EiBqARqTZW5nl72dj+R8P/MWuef/WgOXqMbSnXz5bQ+M+r0TkdOJqlQH71o+krNg
vmg/H1ePkbdoG9MJQKIOXvhgu7wsu0773yNBrgnphGBakQsX3Na50caVhT6gOeZv
O9M6kWaQAz3uM5h2F4x6OfSvEivXrnGacX75NmQd6Knqpl58ZivPINqtDs+YaWRx
vYpo4iXMeMZcmLCakxDPgJGio+/bnvYZv9POArKOZfcNnUiucalaMqqY09GFlo4a
n54RcEZi+uJ21kZjl7JYympG0IoFVqXvdjFTmfiIONBk1HLMIrI407QZGyZkGpf0
ZSIiwOM0J9krgF/WQPemT0vv+6Tsr/kDwNJtb9dIOKznArT6cacoXgpiZr8jSLE5
vqj68S9Nyw7kDP88zCr+FM87MhIafgnFNo/szbqr2r3csK14l1cD6zMAy5UuzsUe
oALfEw/r2Q/AnU6TXP2xmKS+Hq1awIcpoRnQg5wOCu2ITUgmBNdn/9URZ73jiHBZ
8/SIUDWgW7D5kfN3IHzBNx/T/q1AGemsZ8xF/iZMSn9wyk4PnzzLgZRubUPB8ypK
Qh6S1a2l1CSda5AQTCbU+RFro9eWWGYzx9SLjMi5ARaWQQ0V0vi1Ubh5llpeLibv
MCvILjQoYMGRbxq7n8bcTTGNgck/ACsOpTvctDlRDVqyh5qPq8h3I1K1G+jyC98m
fAOjQQ5mlYva4IL9GUyHS+Rc/GTeROdh5ejpK0ddEG/AZv3gfYWblWoDZ0QxPyb0
sj9rw2RZSMJFJNVdaxABuS/LtplVHhVXECdGICpha42CgrtAbjvO/e/HKc1kPlD8
MQky+a591gHE4yPbRpd0UQ4tmD+gfNfmwZoaw1FcvClCOFqmBUJTq065necznXme
ZEH66/PzCHdBFzzsVmKskCS6uOevOIWfuYvbH9Ky05tEhy5eNaDbx1m3Lv2WTTF9
/BVIjm4xkLzYr0ylDcbFIYcMLzIFXuM16eQ0+4C93nskxEMYjW0aTmexs7Q+TfRa
50+FtlZmIvLulOmmQgsGFVe4gqwRQ3DvJpBpS53yBxRHiAIAjj/VlqwpoTJnJK6B
psv7USusSFs6CkEWe8piulZpj8AEPJoLjXaFo0hMOl9KKKQIMlBPsqcOSNM3Eqxe
qWxk8BQz+/u3ybGN5dPHu2ULOLswbwK65b9VBzM8C76syE1/gol5ZAkCTxqSLLiM
Sr1m7U9cByhn65YjR6X3jfGidmk5XqfJfW8FyZ4WjGFVITz2o0YFZcv1JUi2bSRH
S2CeNE6xsHbWG+zQveoOCq52SvTXHDIKVgCKdGZxNrnexj0391VhPHrtOmEd5gXc
tUPj64sp7vkmRgYKaO5u+bgOfPj/XMTBxAGx5/6va7kUq7NjRGGIKOpHNqgqVzRg
PdkSbehnZcdZe04QoYNmJstap+aivUttSer2FFHBf9aWIziARxKmRaHNmhA2wkdD
TwglibrEJjP80uPWksP/xIvpEkZV1uzVfMoOdQPyKLbB0XCg+FOjeAHeMW+y13m+
hPkck98lWZ61jM2Fdo1265auS8ZIBZ1Tx7zoRzff67lWsxJiASf+ogSA2jOjvwLz
t4EtfqzjRtVAQhzoAfLefMaHYedjnQ8p2LvLdNSrAcUqKJvfHWFWJzPY05boNb4K
vBl/B/cpksL2VN/1JHkTtNggUi0Prq84C6mD5v0eklYDhzw8VQxBLQMDRXYnYsKp
bJ9ejCOvDI5GONdwnGIWfLPnxg42LunzOmYWZ+o4BsRe9h2nnzXWxHmiDZxFKtKy
A+OI3JpMEdmkvTpxXDAxBMjWJMBaZ6SkbARKe7Pch5Mvcmi/dL1IoDznfXgTGm5P
5SaqewoU+0qwRMIhknHL/jNsQDVDK6Da7lPutTwyCBIibe1YADnPfe2KshTezXQS
L1XGl526GSfGbxzZtUZ7w1kyAkGNP246ZdPME/nBolxGz+l0i1Ktqvbqjjh8vf9R
DP6ZA8Td8XM2Xb4F3fpgqrU5Z3C0WfI4jzxuFuK5kh/pOxyb8/s4HD8/SlM2Cuec
pWqu2UDCpcVbWsHcK74MYiiIK4jQGgDz6kTl+kt5PHu47XMwaGaD9P8BEm7YVChg
VO/gzO3nKW2KMHRP/xJc9whCE5mYCW9oQU6SvWVuLnKKedY8eu/freUMglT6/Kon
midN5pe72Ihu7OZqET5rerG9MnFDImz2lOWShXAH6IwXYeF5P73A39A/xoGIiN+s
qZno74Bz2cas8sr7/5OCXC/bFLxZkHXY2o24jFcYiLvOsITsZvZKyAlXs/W6TmNj
7b6IX102ll1ybovtd21OFNTuNKjj1h9gH7fSMwdY5xcJxiPwSP2NAoz4pxmokgGZ
Yi91Ug64gaYlaNqvs6xAoV+89wQ5Ohh/gT+YBrAO+LBeKhTmcn+LEsL/ojtoA7AT
3h5U8XjJZV9+Ab8Pu0fIunR9/t7yA9qkA+3RcZ1biqE4/XtNeV31gOTMGORmsFLv
8YTmpoKdwWMpgP5Lgw6DNRQFD09oaMhAsvqk/ho7B0ZaXoegSz4FiB+Cqmz7j6yH
vKRk6InHNptFqqvVBUTfKvqQj8lfOTVQ0XrrM2dgJrFNTjLRWovAaddCYMFlVlwY
WKDU5lhUBRywkr8VnBUOLqHB+n8GoguiLEHEcNkKz2eibc4PzvkJccoW1NrzLkSM
lr057ulLrkal1Zzg/8ATa0j8wvAr2+MPm3R7aLL81D/UaPczMshP8QZ8X7q4BIbG
oLBFa3V4rZMQQymNGwFHVo7akuFBwvMKbFYNVfLQsrOWuaTLoWCNm4XGty0eeLWu
0zx13+yr23pJkRajmiQ5yZknkaBuGhO6R/6grxVOzXjufy2/US9ECztMb9zWXSgZ
ie+USiD11yDd7VyYCA37rsep4NQ5l+QqzN56/E0anf59Y/m4qvPHyDlJRVqzAK/+
J3R0DG7kmITArWcACpdwFVoAfVxD6Gpwixrofm+AHV2g6Nx3otbIC67PeAjlJSfe
0iE8Qy1yg1k0LohofuCTnWBOpX0NBR8eG6sX3xqCGpsT7CuXlQpa5ZcQCzG0AA6j
M007s6zZn80HJ2RRpsE9HOFycN+SgRLa9oXUCgYLKy7YGCtsp0zxP+stuHmyofUe
Sn/Qn/ci+cK/nnwNr7/Gov6MrkrItbmLL3614bHdh/d/ztUs0DZGxOG3N2Cvw5qN
1k6hUNs/5vt4zzFDut9GfYvc+tVBhfVjm48Xtwiiu532WHndMpzEJ0bBI3GqffX4
LxSmK/s+rh8jGYXVDsKDmnOOQaVc8DrUm2jdFlAp/fdJ4P5xXTm5gJ+5BjaLEQ0M
Nxlo2zxNoDK6UZu6AsyTh1joME8Pq2wWK5+V26Ur2LbsJdhu/bwkwzX3gMbAg1ME
vGfkyt4ZWcYAeP2Toxb2AX7191IeG8WjOunxr5OHfsMWKNSrFn7863pRnjrT2Dlx
THJGRVRlqFex+gplrwUPqqswwlB25xXmFYiLNDx5JnpJMSgW4R4DI5I9nfX3C/XG
iRr/D8gYBdU3WHwDAW/s+TckVBl+TghzDhH/ItEkFV07xFMp0RO3e818wiGBWKNm
deSojNpJwvvo7KxbnIjF7M/HB5O7mjdarAG+VY8HpdTC1tDrLTChk+EPUhJKb0nZ
FfPT1pHLFz6/Lb3VeHC12zpc7gwPcxTFtqyRSHjQZPtEWmiHhBJqQ/7Du4gU5rJx
gNLLCCPfrNeJmxsTnjD3i/ZX70uZqjK0aadF6qP2KjsZzcznoxwa9Ov3CvHBhli7
f9YiM9h88E4xDJyWt8NHxAZyopBI9cQJtI+UDHBpYyKN8MEHDO8wCdvxBRSQm/cD
1EGf3pR1SLpg0TOWcOUtX3wZAWbeENxXHlo3h+BbmY0x+S0DnLfVgHh2rcBHle77
xl4PwIxIq0rOhQS6l24sdASXdqPzmwNR9LePUdf6D8N0nmv5NJs8NPzW4Vss7f+Z
TU2k1WcfUo3bsOow1JATYRKJSaSnrGbrzjtmgJ9nxyN3mkJvbQ0q6EbPqZjn5nOt
fkXOOolHoE4MlqvV/lz6qeWq9aYRdLyXif6GmHFkK1gzBWSM+WvXis1v5WydyC2V
hTWtwffCvP9eLg07EGK4PfvX2Db5jHCRUENir5B7Udh/IKR7AAHyD0rkyvBKbjlY
0yPkoZBMx1R+r+xxbYXg1tfXIUSqupc4OwN0H5zFWxKvEtTwVD3yBAEDtxiynvqj
cxDR72S1cv0u4TfgjpTw8GDhN3iom9xoGzkbUl9P8zrmll/1tIEB9mVU/DA31JR0
3yCUWH8Osum71DfysApRzj+JhRIOSsqNccwAOPSic3cp+7n6KoYVc2iIzwvf32DU
ZNeouPF7jgcjpipalxjzSemlyf+CezNO9BTBQP7Y3nwzWlRK0iKyKfX5HV7NAaNG
3iNYesD2SGiizNzbw/ldoXnSIz7PBM19iMIHWRbjRrAUUZ72XjJjoRUe5U4sXNAg
pO8sh4ncfAmXeOLjJndTGnVCU5+RjE0bIn09guFF8nSt9rbh09iDPgnOyGeJQ9tg
uPBxQeHuKorx+Ja+Gj7KVivhbwdTb4xg57qFO3gM5ZvomVsUZ10m0JlNqigFSkha
cHtLTFHJkJzir/5qdEZiO5e2rQrfR8+K65mWdQal1m8bhx1dSXKmKLUWlONUEkT/
27ds/45KMeMtP37ux+9bn6EmaoEjlGqU6ej+NMDd6tQor+jRy7zhCIMzEdnXen/r
whMeJn0AsLqEw/p92/3SFy05Xcy1rFXqSX8mOmrr7n16HKCIYxXCRS9/5xCRykjr
TK9Vws5j9tHStsI0FFLqES7TK1+SQiBAeQN3Sfck3shYJkSxhNseZ1Gkp1gz1bRL
KzH19XalY2OzZuTXrjFlUyq6JZJ5ytZ+WMa87ueXLJXxni7s4giCszz6P1jIILal
28l4RxSSCAUFNp5mVCoRT3WtktAJ/OkQzdo6qpAvsNxxVmrUK/Rxd5KvrT8/5wWR
quHaPmaRXXLYmOPOIlj7W5mDFqmXBEHdEKR7Y60r0YgWit12CzJUomJGRQ5MxUfw
Ac0m9Ouc+6MdCOxz+xY5vATyi/59/WXj3b//NCvPwfTdSU3ItNaPUYbwfgFuMxHf
5EN2EtCqIh9J+8aHce7wVWVSaBOH+gHJZtJdUZ+FP7UncZWu3HHhcumT0GAS6QOP
ASRd175/K7s7xdTdwtCQ4fHJ+dH4I1KnD8gAXlcYOkk9s0fBSihvQ7HqWmBxelVO
9GyFELM663dDrcB+FbRas2D64mg6+wSGMao4QuSKgggQytr9f8dWKUwUywlO4IkJ
RJHWlDYuCqTIYxKhlulinhA7L9ORth9zUSzar4qJvBn9Yj2ccA2Ay0gShTEXM5ZC
4e1nLnXuI6wYN9dgAHbpZhG2mgG9RtaaQtJU+1UTmwbH0sALz4fd3hl1bBcjiWSa
HMLUD67IohJMtjEveZ0eTPguzpJRekG6ABgObA0f6JG4QR1AK485+SudvsLgbW2F
c35Is4akSc1yzyd6LACEWKrOrtvTE3Ar35MG7maZmemr8lQx1nUjuOdoEJUtWvsd
ou7/TuvL2kk+vYPuUhqagXEb/ZqlQFg0iS7ew8DzY/48irUvfw+NSU11+ui05bdP
lhnhc1VY4VDoeUxdH02wnG378FpOYcbk1C9hbUVw1ZEPdGUgRI4Vu3zBb2hjXGhV
IRtmY036zHuVEl8918JuArgBi3UlZSgWgxqBnGfvZNb1lP6wv2Pm3Kv7FoLBBK+l
Vg/kFBkjb+LSA4XzG2bfb3TYzf79H2nooeTL+weRqPNkB/h7AF+RTf3fsvglNZO6
qX/f/jxPByCZxJRHzClkQj77tdp/CNGJejPTiXDRzBUa2MF1Xmh02oKJRGYs/kW6
vfpMEDPISWZrWDG081luOqmbQzlnaTaG0cwbFBbbqq+oXeEXH5EdN2GiobR3UzIZ
QAJQmNcf30ArMWVwyq+FysaYmoUzAJWyswxhk3IZaEkVKyQqU929ZhFlniY+VFnq
oEDsLepZlBfd6amajbCKqlOiDFfL+EQv3U+d4p8QOy3kRYwdzQv2LieYdV/NQDV/
3VYKsjvGKnWppa2qil5YIqFlupZDhLmWs4dj8MTz0N/wOo4YUi5WbXjC2GP0hHek
fHHPnYL8esm4M9p+BOX1L9axBiV8O6yt7eRgR0lOkvVMEYfrwXXa07rDdPb3vEtY
6sxcql1PmKqVTMQpYOJusDYyzNaxxshhfABGLkUBCMYXedocxevLCPMOnhYXpxsL
ykU4bPEJdgjQ8EiIn4jAo3T9/9hIozKYa8VeDESs67WLfjznU5FCGeTDoaQzBZjA
3goabPuCAvV8csBF5qMreKNJ8S4Bc91E3rVfqdmu3GPPUqZC+ymSSxokVFs87T8d
aT7p1A9PjoRZ/jqSMD4qZtX8sDIuluoNRrNt1zwkVOXjKbjCc4DAD3sXSPAoTArY
twjXAZxB/Y19h98owQOAxAoEhFFp9cpmSH92lDZbFJLsH75Qba1UH1iLweX1slUc
ryQHU1SKJUsNb/hMK88dQMxrudxsFhEuo/uaLDr5Yo185VddQJqAMXzWgdkwoEDx
gJWnvwcMw0qrcHQ2eo3oGueHAf3cj0zgm11fzr5OTMr0vNNjjWeOHzr/Kx8g69xU
x+ArAZ/w8bwCEdD1Ttp3YFQs63WUjTREooMhunROOL2WVcz4Pcb8CMKNOLJtzmL7
xOBxcYFzAxHKCrYy77WwWUVUHYmg7Cyp+URwMJKvuHe9nVCMxkzqPwY2lcq2bYqP
ux235FU9XliCwvLUFbX4pFE7mdQFHBFYjeGk+/3dw2M3qwaFvXus6DpMXvlZH4Di
0qsNyu4cKTXTPQYGQKYUMt9go9ea6F0jbEC/xlU9y3V/LZbTgKadUbLkP7UFbG1Y
bhKy14QKuw39LQ5+uEfJIeiqn7GP6CX5nUR/1e1XiNZMSsNDE3Oco7ANFCxyjkv+
lKV1LIdr/1hEauePAptCHXlhzHoSxKKd4U8qVrcVQEQrlwGeeTxMS6MjeH6v0+ut
vrTzfjBi+cBKSiYhE4qTRdGIZyVCIjQJNde0ntDrG1cNgUUHn852+KklfCujRECu
7Al7FIFIGS5Bdo4DAsvkrBOm3bkimYy/xCxfqbtSV9Nl6uq86U3+Hc5OAZhS/a3G
mHwWZHKTf1OYxwHCiIR2xHuUL7VvJ2iY8GHrnQfyZG9UgX827ukzJ1G8PLh5rqX+
hWImEyN5ytehfYwn4vPp//qVjtxdwWzv8aoA+gIoAP5MtKWBQtTsMtPqLtzegT4/
flrXMl3vUJxM3kuTu0YonRXQvMgJo/Tnk5pOsi38vAsSjKAFIFgaROJBex5ClHwJ
hwwdhDhUGoomZy6qC8EvLLLIqgh/JSpNxXD0J6t+6OIXoMcBlJYRsFxCWrdQ/Qx2
MTYBET0F9fben2mbklRqNS8QvXPxk+DBL8z1si2o+bsqm4NBKPRHqeaU2Mgl+YZ1
llsDLO6QoGs8+j6ezsCcH+AyHIfATxDPvssj4ixs//Ur5XMQJGt84N8j9G83ZBDP
tekJgWnroEyOrGidW7p/e0IJ2xh1vgiWuZlgKNcS6uyJYHhcRdIvFFkPYTcgYEyI
f8pBMKY0DEcnl209qfOdWxMy66Jm4w51Hn/5Hd3h13L2TzOEmBvgQLZVR01OehrS
iITWnLbr97IIgKmpBYm5KA2zl68tmC8s03U7wWfa9ufIHTXn5pB/BFIhGvlKJuZZ
kc9mKEx99jsIug+cjnWtrgQPrpWP+BT8IcOQBAMIMj3K248LYmm30/XQYgkPra8M
taFtVHvDkbdXENKq1O+SiBF3VyTJz9DFQP27vQkFGHJ/tWpH+nlXRM7/HJnfq3s+
QQjqK+x51CnoW9qECWo6IGy//XyxnHbSIpujhWkQmxEIOBvtfl4hQWrwYYPuaAoX
OdaxTykLJitX0gi8vP9Z4X7s5o5qndj3fRoriInWlAzBdbctIrgPcBCidsDar8Y0
z7VK1K4tS8bYwq/eAqx7BFNQtqI9qgx+8G4DmOpScxGH3wcKadFEJUipRhAcPl+Q
msMnV97rBece/XNOH+lkDbQCg8s6gEsiZZttnv4v95RlXcAijrqbUq2cT7G2dIUi
FC5eoJzHPZ8d9sq8hEzaF+FQKLJQO1w/u6BB5Db5omLNbr3FeOEaXpg+Uh3Ob7aU
GEeIM/CnSJmjr59s7lNwgIbV/nphrNtVTDGMXttZVwAejA/cXfz+cRhSK31wSqy0
YpQre/W4HiDpVvxbloZFmXraevl4quO/dx3W9U7ct4pNvQp4XH9wbTcqyS5nK6BR
HOA1yC2yLz/MPgSiHeIwt5meXTiAZ+EnApaKsqcHZCMpsEk1M/uRfT9vLHCMsTLU
EkYmt7v8iAB9JQa4RKUeUOZnptWyWuJMufe5SSsg5Ir1NFjALsrKIxLe6CNAGLXT
89bq+CYHaYpJK/USuFc81DtMueRSOOioiAgdBu/huJynggo+leEsmYBu0fNfd6bP
/6Vl4WUGSfSfyMNgszVXTEIpEjSG8r2lhqkQM0awD6bc34XzSQ8zdwvJaeXoCmjm
7JFjbRfF0LtbGkWEpEGj/KnGChHdD+Qi/Vl+g0vN3ySZPlEkOjnXldtBTnpytBLl
IVmjYaTZU0pulQlSJqfkf+9CrmYObMJz1AeQPFpuk+bu5EIVY3kA33NAoGDEEPEo
i071+pf283S8TxlQv+yIQs1DtjPh8fJ7h0NZopF+zPO4qghQp0+GwAib/chOcNMN
Vi+23RU5m5ITWKvkrqWtRf+jzNhhCY7PCh5+NLdtF7F2QePQk3SkIzq4UPeSvB4j
HsJwDgfRyfwvdlP/ND2lLS4wsY/4aB/TIopYkS5EPJO4AhEA6UQf+Qea9FmsznWQ
hPJPEk9ikIwjtR7AwlL4RRfxVD//1tZWakk3pOY3nnPV3ezRuwo4Pi1ZA1PhNME3
vayphcqv/zxqe4kqWmIIOxUI6AmIIQTPn2h3duXw0d6oZSWBw3+QzeA7aSfdAAUR
LjaV5TIGd4pq5eMZNrjmubTbKbD/873++oVe4IfyC2jrH+m3c7AEieibP92Z4T+j
PXp7w9W08fQ/IwsXtBVDMiFzKX2Dx+qfOhKSwotBjteoz5a8jlqAWsFLyOXP/fhf
lS1dGkA+LDI/r8haOvDwhHNfA3hpwOUMmZhM3PFX56jUpK35VP7YtADwQfYjTpQT
zCkfSkCxZRzWke06iC4bpqeZOpzWtcPU04CxEqMBdrqPThxSIwa3k0yNuuXeeCIP
tGsnHCcM9x3Tp9UP3u3U0egliWE4FTIkZCLgT5s3BLUvUsQGJEBTHUB0vGOxI28F
wISqc6hf78zLfHR+RS4TMUHUJbvdrHAg4hroDKWc4/qgPmYL2C/hbWsH8ulu3lOS
F9raWuCmpH1eXyMHvuziZkpGguvKOhMYBqdmgIZqw5R5ySyqT5oeikp/Hiojinbz
iF1ecP8oVYEhAy7VFfdg+aLjS0zQ1z7NyZO8G6YeFx1j0+RGHqs6iFyDljwzxX6m
jhBfFN2oDZauMR8sSvXamdAzamvmgktxMWoCpnmqkBziIZnONX9x9aGq4hMdkAZ0
hU8yckV5z63LoAQNJAybUpyLzsuLhtZgU/fzJNZadNvOf/qmYf76fX8YYM+OuZ60
QRKtfLLZMmQDXWSx9hpqmTuASsSfFqzXk2LvvAS/brbCb0fFioXbW8IifkKO/aO5
osBbdAS/cH8rB8gCMnMBeK3UDl2FXQIP9KIkxS16JdxSaH19aTyS4k/VRe31/IMR
GgBTxxwFDA56VgYpBvHfmfsTy3vGjAxJOBxwm3P+ygyCXtMlEXBcz2lgFFg4vltP
tN9keYJzLwOHHe5z6zYq4Jz983CW7QUIKaQ+niMJHSUXx36iwWyab7PF8PZ4I+Pc
TSqNnu5b62Z8ejLSIs9H78hFb6wqKfOZt7HrJOiWRmTgsrPtRLykN7X6NnpipbGq
oNq4pA7rdoyd8AsY7uIsDhO5uqAdOTDwCBHJN8VVxp/4C/F0EDrRIm1VlBZ8H7Eu
lqDmMXJ7OTTqdo/FOPznjEl0vkZdX1eGJCbqDce9SvD6pPst6kfj/K5Y+/wttprN
OuSDtZtVG7HAutkSRMtjRrjFKIPmmAdBi1lNMWBlyiDTKemxbUzExajM3PHv+nqE
bsw4TdL/CcPf2xOr9CeZWdW9b22csvl+79zhgQBEAS+Gb9I78Y3mfBaO3w5EGtMl
3kUh/c5U5yNb+vxv0SMlZ4ReVj0xzgm5oTwZycXorJHsU7Il30EIls8Aymf3cOZY
WWBRwLOdUDiokwIwm6gCegnNC8IdMoq87J/7sDszmaG7xcfnXWmEEJPwC6Qp9S5v
UplxxzC/3UtyNK/QKhx54PfE4hwKl4jMkQc6/66XHulQMfP9sP+TJbpeDPqPAYvM
A5XHLY4kVMKdgH6KhBdq6enaLP9PrlodRiS/o+ftpXnb1D64kQP/TtR9nwXgFs/a
O5TLWR7LcYTLKMmn81qLToa/e/YRC66vMbFIkZ4VaTRDYSAjcAkq40lpAxd3hByf
hCQFT92GGEaL1qCsWXV4Nkh5PfCxeDtZihKvxbxBqLYG2XAm4IZYuohmURluegI0
0L1SPRWzrTmRv6pcA0cZ6QTKXHodLUb7zb/aeRU8PsHUNYH2m+CsM+dmt3eSlAjH
5x5Ph8h6gkOo2nhOCSGTQS6JS4fSnFS5MeCwMLF5f6C885jFEz49G+Y9cqMC22uD
6+N1ea8t8CGdDpwTkmTSEtYaMIgeR6vuLUo/GtW4bN4Jov/5IXGQ1iN/+1dzcOoO
FhKJDeK86aG/Xop6l5cw9afUuZaLAhzo3dUw+zH1M7pOJNUUuDhQmexnLWqAFe7o
59I78i/KDfLYTUIxayezqrERE16ocUbYhC6iQ9PdJ/VT1aUzIiPWJvXr3YAV25tg
YDiAEJOEypcbxjek2GjW9XUlBDS8hM5YKzT0yAo+QID2HomcvaqYPbU9xr/18KmZ
CZtRgvxWig3/5qYAdlhehmZf4CI1O7DJRIi+ulIlZTHrTJtdWKsRfq9zDaS5/8WP
FP8cm0WRBrsyVMTU4jwfQvRj6YuJqeYOFpu0ZStS83HWm4E+IgqC9eIihHC1ifJK
4djrQq7AusLETZkfw7Mxt8PbLyE6hLzl/kJ9q1NjbnEP4vmvJA9Y/p0vYpUExq9u
JLmC8OCrgl41H7fvU8e93y3H20ilx2b8btk8+0am+votJRTPoz8AoKXt66cYNwg8
js8XllHdULrFRKW1/DWTToX65lRoXTi/pIOSK5HqNdo3gNZCj2DzZZeFknPiTnN2
54S3UNt61JqVl4mscEEFlb81nJKsEsnjR5QjUoXI2gJgpH9XhuTD8cIHRh2UpCrJ
kQbS0rpwGzKBar8GBAFr5CvTTstkteZ9LXmCYM7aGg2ZjnAgnw+KqvU1qtHf8153
1Bw2QPk6ft905cO/rpY5iZDG+qYgRF5bIVW2vcxHPueub1ZP+uPZn2Jn3nJTVysd
W+5IsLBETD6TnYT0KtK3joF0xab5wJqAbts+kPU9B0FsqmLpeXzJ6ywpXtnD3/cP
7DpI9E1NWLxH6vqLeX2knk0BuJZbCmGuun1aCbbdylGAkutCTuphxbiyn6tySIb9
YcpCm+szOwIKOC4/+YC1SIitFSGnyDRYZnB3NKvXHLqX9AHmj7ThC2YRBLtMKc/C
wCH8767snZzOEDg3sO8Da+Am0boxR1tugk4v2ewrtAswdK6ZvE3Ydp23yqJt9ZlZ
8Rt3ut7EeCgbK8Mr4NdikLff29bzBSt4fcMqmrWSpqknLR09wbhIyeWmb7CFpVLv
UbXwsmZVzZPZjLDvhQqo3gDFjQArxFy78BUjdhj9kRwxrMx1DYcSG2H5et1Kc5zr
dl7CSGt1MKB9YCrl2NSr4BiYU3+kWXIUYOhcPXMvGWjRvjewbSH2cQvofiF9PKlT
KGkKzSY8Bzrpj1ZNIMIriXMlU2ySuQEI4r75PY+Tqt3Zirm7/uLWcA75og4ss/Fi
JExva7dZL6UPbY4tV20agiUPKaiCPz9tuc5bZ92O5o3CriRmH0tEAwp78DyK+Z0M
Aocrroh227851wDGClhz3zHf5w8XD72HkIxcLICTqnc1MRKcICrbIvMvA43kac9g
WQMloyTHezfLIBWCNZEUVyj+DqYcOL3pi+lk8M3C3L5ubYHHME9/W4b3dfoUk3xk
vcFWgIDjHTts+V6AUWNRWLPATkzEyljh6/pYpi/vBSs7WB4wqN01xL2hUKAP+xDg
gy4lOESUUFktvaY8PLQvKP9YZGeqty5yvttRPXWzFV9h7mu0vuD9NwSb9MeLJQrs
ulLMRH+qrvGVqTUKsCT8SpwjMNyKWEs2v3VYic24OhZOnzva8fgSg3XvqzwzpL6g
JO7QNkzIiKQkhHALqT6iCShB8/sfmL47s5chC5BcFjHz+8KC+ukbY0HNKIpzk1rB
4d0kAQgtQ5KYpV2yysV37+AJUnCVsCvOQDC2A3NiwZBpa5PlEGF7sfIF1I322U2s
QS0mPoSAcBk+1SNpusnTSyoz+iw8BCnhCo+sZsEnYTUzX1CRIR9cnYclvUrjoFe8
Bf+bkqiGEdZyMQ+zjWlI20sGDrzVZNAhCGqQeJsAp7dJPNbBv+1dpH8EYgqgmcdu
9eQ1U7nr/7XENT+bzfWIo2vZZsqLshArweYJ6n8v014RnkWEOtfriswH+Vx1WrR/
CtVK8Le5BDvPEP6OHK+1VAasPaQvIptjOXO21zPZym5ipUZoIf40mnA8gn3aCyAd
hwunvc373oXJacWHIU+my39DNdRJMq7iV8Iyzqbg0DbDG0Gb/urEIHLlBst15KxR
Qml33+BEq0gBKxYN4T8zTGpC55qKqxuUNu5Uos9H1XlpxH1lZk3ckoDvpxMKP+Kc
Ev9MDg/IQWu5XQcdBOIDiuJtO0TP/3gkHXYtPsYCL6NuR6Bh4gy3Bwi/mes7KYaI
VxzwEa2+wjUI/n3uLGg5rnnZxxM9eubPJj/9ZLBzOVnQAOdK549PPlojXm8awQCm
mL2Mnzai6ZkFuJx+KBaVYvz26IkACQ0uptH8+YcOAfi6tifwN+kkKZManuaieH7h
QxfR8ODh8YQjQzD0M+4Z4zJ6fCsjIR80WmXBiHavUGp5ogcEbWRXLmWDUcZtY6HG
+QAz1M/v6tpz/E9L7lMlung5o9z8N8gdPrg5Hg5gLMzaC/lD0tTtyjDGas1d+CUa
71n7qxa9omAhOHQTa/gSgS2Iu3j/hqVsvwRvPUQKUAzL9k9qJ43YRHPYUXlmUqft
oJEI8ZSQEhPmO8kw4g7LvW+J+RZRKvX7P5aT1AIwpxn8qS6blpWnV8lzPqr1mmke
WtcojlNTNzuEct1MjePC3tVsiJIeuEndOtNVJNpdTLkv1LIxOxGMc6XYg0lLPiuU
mthHLVr3+EAJmrj/TbAzUy7crDnpjGphpfoSSKCUoBsraNebYNM3qQm4akfk8ZWq
8yrqIRqg3WWS4CiNa/iYwMDpmzSN0HbLMcHnF1TiKWKhtTAh67SDMGNfxZNP57yt
6WpPJjj8Kj2pR2SFwF97tVhNPxQ7awC0+Ov/ND8j8puQqxDVRg4QCQF487kQdrS2
mOaJTTPY3TWrKf8cz42M09ktXwvEKARqc+coXd1JU3+LzhS5mgsJwnQ2iJaUHIVu
St+3ZygPBIWfxwz+YF05wVXsMu1oLboJIMbVk0vaL12vtjYQWi6+iB+m5j0oU7lk
HiEjIR21w+lJe2tgPcEiZLHgEa9JMp3KmLM0SwUsb7I94Qu8iuXmdGij695d1ufq
jEWjISNrn7expfItkQUPoghl8qJ2ZxgXnv+bBShRPNfbJHPo/1/jDP881GGzy6+K
7qD7vug8UkT/8Am4aNo5mqEqJSLck5a0zllsgQKHs4wqTDu1si3u9SZDkQuLijYv
jo5jCiKUgeWdQDQX7tspYY9NcqND5mg3FJmTwMGO6BJ2JSQu2v2CkOn5pIa/BaXt
MgnqDIVruQ2vuspcQDyjMweqbqYJlEECMFICESF8ICu9LEz7G+KOgRXDMuqpXQi5
IQibR58nYXAfceiGOZIVvfqK8WmMOIzyj1HfJr3nCTbz/P0sXZK2BLgXxNuS3bzo
y3deDcTmu8KGnwEfMg5If9ViMo0SqDplobwbfAfYMffhjWGs7b6lBfI1jCiiBpH5
ddA0n5RH8sWOHMB8ygAGm9FAH2UTqIlYyOiGOL7opGrtDU5D/CFNDfjvL1td/ift
UIDp7GwvGdvk9iCR43FYS6FY28+S38Yj1pbfsfb95QkudeUr+dukFOanjx15KgKL
m2jgQEyOtmfUbSE6729Dchc2VQNgwyI1FJQ8okdj0MlZAheDKJ+UN5IKjWC05kRU
Hk/C5aNV+lP/V4rALqhW1BhvWwNuVcur8AUvNcpb6dYthn8VSMdn88yUU6N/33Ee
vSv8zzVTDEPVF8DbN287Z9xwUGvU7qlPiLWtRszj+jvj7QfZ3XtOob7VCufGmEsa
9Viao2ZDrGmR1CWrUSoTx4lE5abzz2DQ4JBBMvXcTejmJlT52JVyP0Z4nauL4hwH
m+iiCNW3MoN3JHhPLCKaH29do2Q7PM+bPk9u+NDa4scfdB+s0AJwuv/JNnzn6zeA
Ovm4wcb5OCBDoBeCXXzaTvp4AB2KWxQNiLscGfL6XMhoXEQ8hHJ4rTpfQuJCah4v
JRwBon1rh22+unm5YyYAKyVQS2bzKnjsdvWQy7AuNMTBa0opDfuVQ2pVZuI1G5qh
b/o+2La8519vBNxJMsn+qHaT3yeu4RDIQkcO61eANm6Svqv1Vl83cM0/cme9v/qE
d7Fs0JWcBY5CWrpeNUYM1QlMxeoPB4LjAFZcWQ8hsRGJg2Y1MLNm7uINFfBGTnWM
iJgEQL4C2it2Sp+Yd03DDCvoqlI07OLzAMOweOgbcLeIZ6sORY2V4gJgrCmgyxgj
cC3itiJe3RaNftvSuEOuDc9YkgaIgrI5ePJ+MC9ZWoP3dU41WTLgxSjIL+EvUCeo
IyBdIPGqH5aV5sbO3OjL72/TIxsaTUuh3cxAe6KeqbBVyWMpsgTGFAHVk4rULgKn
0ux3IFKIVarjNaREDjKMQt0caHpu3ffI7mbV8F5dqbl0C55TcSFgsmzV6hXx6RgU
hM9D+vS5dxex3Jd1g0IVaZmoMq81cfotMPZJOWmuKv3+nGnByxzA09Hf484ZDSXq
RkV7m7I+uVGsUftBP6OH3x6+LV5llEq3zOZn8Ppq4AFwchU+Mkddw09ualB/uWEo
M2tgHrJVe82Ej2ZViUokJunbkQAgZx2GquxUf4Va3cmXnuC2eDYC17pYj0KtkhPM
WAF/eSOqhE/LSm2x6s/tEIImwBcqbLJDyODuoH2w5V+3uk6HdYdBRYndds2hxSGP
+q5htYeX0GytJ8SKRuV5/JDpWbzOl9r4yEfzyVengaX5/+c236MWQyhhfUfg5YHn
hDquZqcR6/k/fxmY8mYXS6acJgy93OvvVCtgvT5+UuF2n4GfK6x1W1VIZuoVqlg5
r+9D+mgSY4qOPUd7avHEpcfPWSYN9N/nxh4CHexMwK6BCdhpBtClPu5+gNpY8+h4
Fl6cNtAgUkuv/DvL4ebMqaNmAYSqpdH7wpj3EJWW6Pw7L1LUqx6zObEhxmULFphX
je12hmDM2aDppXbIz1OCwqT5eb3EGnoTb6Yfs3Lo4pOBVISe2gUh60Lz26FQcY4f
bHZjiMIJRthW2OycqRW9c1dj97xnFKtP4CnyI5I10rUTNcKy697wFTN5iLao0Z8i
/a/h8XwMvBXvk840y2wq2bV0dnI37OFjFrH51Qo19qCH+sAkr0LxaV5SI5aeYs9e
3dw8c9zmx4Yk1KlRWzHXnbdf7p+LZdYtxsMWfDJlAl1efoqcgi7JzFAUBxNBtTpR
uqoFJCeu10YJZnYLGA3s3b6vcyuprndNzEqdyJc+PdnB81jk5XjHuprGAwgz5agp
OyQAcanmAvi1zWN7ew0/66qtsmT7jVsQLjLt9LAOX4XVYPI/Uy2moEbgwyUDqVVV
p4xFNU8B2QggcHYZurUBSOr22iFMBlubc7UAkFkYhToPOozAAokE4wsKJvP9fBLm
eaq2XKEI7BQbP96k6TrEUo8ODoIfMipXhQp9dtBhqAB9RmdsicPz5z6iobi2WL+W
WSGKbv6Av0/Y6GyuYi1FlzTqSj40P3EH53Q6rHM2N11ZfNj6ItCWwLtS/nTxvVAs
8p+D4+mdJhI9QFHTMuidGnBX30Bj8t832kWwZERIGrpuR4P0L+uIPdfDDlhuY0gY
BdNuxcqy3EIYBWJSOpWD9OkqFLYA/4Yt0iy2MTZ3uxojIEZz+B8wpBEVs9kSytov
P3q5enxF0cmGED7xQtz+VFylVTSzbLZqCPPzW80g6U43Zl8OIbT8WEz5npbIb0lR
gdlfCHG2FOgSJjmtdGbo5t0Sf15cPLCSLuUxE2KjQgicDWYX6il+PKfEwhpVnokr
FZzEzrWJ532rzjfAK1/Kobk0PsTtK9GbsgbwJ5F4gfC5ZBrjg3B6Lf7BMulc8K0y
44m73jR73BK8xXNjzmoZBWV3c9enLejjSd0s9M/bWLLK7MPWoK0SZPDsydZwTEGM
AUyAn+J6HHeVrb1Xih49MDu43RPoyyfGmudqKzXJcVAkR5EOh1X3L5Prmdq1R8IN
J8Gh6ylUXTVridj7WkAIpJbXW6mUYi+z8j+HfNCyVGRfc7uM1whVNH2tdAAwDeB7
2m9esPV1SWu8S2JHOUftEiB+D6tM2MSatR3G0N9i1GAZiX/Dp2t0EHIr/2OcZ6PA
lOf3AhX4/4LRpL2ysZdQ0e3jtXGfBSESizXlidk2tVl2jfPMee8sK6qiOxJLGsRt
1V8u7xWL9YQZA9KtrTxJdCWd2/neVo502ap7k4uQzEdb1mfe8C6Mby5NA+XmDh88
CVGTVnVfxXzW+JkH0I94unoHo6dk4KsmFa79PFifkpuyKuftw7+0Wixibty1yUo/
Ms4a9d19eYPF/h51F1eRgc7L7c07bJktz1ZeR2+6ax41yp2c3gyBGwkpKqho7co6
Unzj8G0I7ePEiNAQfl/hU/rBuMXwcEzEIpIdS3z6R4Wb++8IQ8M/Z+1+4UXXQ10V
5Af+d6+Ke3aCVQ3uvHf2BnyoMzoccZHU62ZtMyNLUIBZEe1sM1R5p8oc3leRMloB
UBSbS5PSwsZ+Cvm3d03R025NUfSm0qAy3/kpFAFH/MEUMtTxUb7pV2wADuIzsEhW
DVSTgiSIHjLctVlo2G2cTEhITIIn+FLCwceKcoOGhcfBVVEjAVwJlLdEFqZfQt1n
m5w4lH00IDAxMAs/EokBwn2oM8nVM7/TA55+ouVktiEXuGkn7TOrGiNS0m336GOq
TG9H6hf5o0wMQdf55Jh29br8NLCRGM5tWC9oIWsSPZ+J1KU4hgSp4F5mfJKSZ9Ay
6tKi/3Oot9W24X9rTiPHARi1CCGOxSDSMibEdXVWXsGfa0xxkjHzu4XVa/na3Ods
75QgiIq2hd53zzgPyh5JoF0hkAMXu+vVcFagmcnMkpQq2mX1iW5HgQnn8dfk1HGt
kfDdUmZtpjqV6dc0CSOoaroVgI5kxzamk15awxlMfjBjyqOmBOJ0pbl/Az01HfYd
SPj0hzfr7DvD0X3lqNELOQMMg5DjCU9aXytt7PwyvfzQU3To8+UCTdiLxDIXuW4Q
MSGQep7poKkT8yImWZbLa+VhaTvTC/i/TNhqfzLkcwsvm/OzfDO1Cmfxxi4g4Auu
tgaEc8DS0f0oH6bjUxsQZlCbUQW0/nxdavJrJpbGIaJqUdT9v2z3MrjOAxo4zV1T
ozd49nhEh3pE/BqNZ6LX3QjoVwXDcSHlT/hYfktIX5/gNTGZEdKyygh5galnaUUd
1HrdW4i3GMznLtJW9z70VzSvIkfv/nWfPQQngJme5aZBp6zlYDEracMFC6k6QZVi
OUsKGKAJwSmYQsrR8z2PGtqTSgFXSl0RhRexxcA8xTIC1B7RRaLL9/aELpwgQXbH
amATOY+3ev4t8ewKhWWaksS+lMV1g1gBj1cQ/1CbyEy4iIyl12agRw/iuUGcoQRl
aMR0E3+gtu57qCfZ9wn1L5RX1XysQk4aebw4mYrr3U8qPayLp8tdi2VqGcnzeo3g
G8ZehWDtPO5hvFt8J14IJeoUzaYouobdo1cb40fnBF1VGfy86bLuboNv9szX+EMx
FtU9L0aMoD7KvAe/IBdtYhJUdhXFHdW28tHHw31SyugGbPmmq6f5kzB6NzFKEmxJ
Q61aUokp4OkJWTTkMHMolVzh46AwmV3URwH8lpIXHosxsIPs2epcgencVOUjuFbZ
TVRPGIVyvnUa9ByPSh+5/k8gYMrTn23J2PeKT0LZLsFlvUNJ2nHNrJ5yujg+Eln4
eAwlnfb7voiJtUWqgddTHyVDyO8MnzqvdhqN5m3vIu7GXuwOP3L80kES9CtAJD0j
pvTAwHlEjqaUWyt+A8PRGJ+zQlF7OEc6ckh4FYE+JoRKgCMYgkn4HPVrD4qTTzp7
XfJTcemK6lI7+960obTRU4mjv6neCr8z6BPbDI+DASDYoHb+Ie4LxcbyLCVFI2EU
uuCsUbLlEXAOLF/BD8HIqY4R4F6v/8KdeK0desfXBtXSf1tosZ2iLRmpIQPC3gpc
AAajlCrl5L84y+0BVDi+EOU+j3DbTfGNgSeRvt/n/q/gNKIoCrfcRXkzBYHXLTkr
9m94I3PNzNb5i8rs4WhTMS1m9dHsMS6E7R4J1bWqy0EAx1WBZF43Dastxhs2vcwL
aX127fX7afZT6PGmY49hQXUQQOXvQTifsfPXwE+9A0cwrgGozS2i3mQpznhxkfAW
CzkkBCEKrduIEwGomjjn8SmZL/jRxbp1U3/CtJWZvrfac+9IXaMBS28upPJB6wK5
lCvSU06fCGhTBL7e6a4KBts+pRIWV7k9XxlZBoUWhhzGUbW8MJcmVe5UZkIYtYCl
U0FbI/JsWqKa3ugPSQrnucHpKqj3sZx8Np66bVxinO3mh/rN7BWu8NNfJxTqorea
sCqgpSn6kbhxdhCFWirSyQ6woHeZCctwrx8z0M9SCgD95ScZxS3QzpUD7t2kKvdF
p+/BAFCmzzP4jfQH9DRACMAH16DbNdo1bnF8kgngCXDGseMA0DOK5rH88Mw4pzi5
tz6BsGr/Vm5Uv91uuDgUXOsawnv5inVZhz68fv65Q/f0+B2junAp+91XTYMJl2Gz
LMheDcfYU+18wvdepkzzh62woAYF7rb/+NXu9gHqUPdPmX6b2UBX2PdTElvS55bW
dp9COP+kac6vaBlbsihD2vStC8SzvAXUG/fFpKbsZ0WtVUAQNExeYSKZVRx7KN6P
qOiVKID7jvSovRlZ4bR47oJv3kIgMPx4dJ3XMeDZv5eXMwpWI76dHqUGo98dJctL
m5N3Z/NX/66tqgl5+BP0iQIyLF4vLW/G3s29hXwMecgs0bZPEnQw+6JbEUSzA10o
xE1pir9evNQ7bZiquE3S+1taT+JBTn4iyyT0Byi7j3jSuEHWQg8jN0/Yrg0W2mDy
Lb9KBXagwQLGpYsk3CxKnvtLnJDx7MmcrlERkZ75GSFCRWBlu0TJr7x7X+bMSg3p
qKIkVQ7qLZypYZGexf9UOpxkoEmyMZJnJVCbxHoR7jXz0goxbiIQkrOjLAfhaY3M
lfHT5BcuvmBongqqSfbTIA/4uvhXM4CZoV2d997v8/GmhPTNKtQJ7zYQGFuyzUHN
gEf3zTuKzVe8R5e1Vjiz7/Djz7Ux6FSwpBSPCAdAXDt1cpfUkAKJRrQ1Noonr2D3
3e56WbNAG1T2vpMoXFXR7fngGmu/QIojs+s9se+uZlDrv3xJx66JZeZOFZXaIXsT
O7KOfpLTXwij6mNqAbtfcCiuoBMzCbBs1X6+0SKvClqGo8NngHc2fJ8EPFJCxKTM
chjMC7fey6dnh2CPGldUHOU8ve8srIZD1s5FtlzNTePgCQ/UqCuLrDD0QLI73WYc
+q9p9ynZ2GVHzuYW9VCiGGlmyv3CMPfv07DvzkY8+q0HSgDNvAA2O02rwQxmback
1SsJNep3fYxddbIVdDCpMXQfp5uSiHl7QBmHamOhuOx5XBSb20UD69zN536Sszh2
yvNCegmxfBNxIov+xVJay9b0Vu0sBERpI/mYiPZ0uIHr2PdHgiC/tyIMIbQ0IYSB
66oQsrtFHE1hE4Kq864y9aPuebVrOojfTIYwJ5wN5UrUOWVQEUCVpbje8E372lZe
9zrfOhCNM3JZc441bywp4OaT4ks4AR6yPQCLEUGEVRJBASOyVHztyvALw1ranrEQ
qFKz8tondG5pAQryYnEXczMGaPtGUfuLdNYEMifLPzEL+5yr8ceOXCARH5npFJSW
jaLuBKrrH3DtJSPnZ9W03FrOAxvZm5TBY03/AkJkf6ISPVkewUtVrUDe9VOkNPSZ
O2a7re6HslIey7xFATI4sUsQTjZXJzLdpVkhlGAcUV9UkAYwTcywUvE1j27a0Z4p
yzqK+E0EZufoygvJ9QWrpm2Xi01eOByVuOn8R1enCIuu+Rg7PijWFNhVW+P2sNqb
MNJb6J3+V4hbgOvz487k0jKbt0y9dfdTCwJuIEXnHzf10X+QRF3yL+LmagrkR2LU
FKQYdoA3rwo2/jHdmEg2BC/E6zrtELFG7xXdAqmLcBJuXPBMtNxqGRlEXmMW1nKP
QGkBghnbolFXZxTar8f0tddSCWWSQ5iLOaNNwctP2OEa+1PgnSy1vfu/N6VQDfYc
dp16yKkdhi8joMPBLhKJseduMeawgJoGyxTqQHYSvOI2kE0IlyfIrNxiE4JMAjCr
GIhYqih2JYLN95HHY7R8R5Kbq2/8+mYDUtBypzcCywCDry6SKkoVgjahB2rgcfsc
3Y2i0xOcAEyXDEiBY0Df2zF0Fho17vPksSImvLxCzu82aksgz00OjwirQpaq+d//
XQIbeGPHPe5WNwnsl805czZWoPQcXASa5hau0LwPow+twGbd5m+vjxOfT+L1v6YR
6Z1wyFS/qqu/21x3bc6IuURQOucXBfVf4sCK6+h//0imGh28G6kp6E4b655WKeUQ
B49RKe+hyxxRazp24sTWc0S4hTTIabaqBv/u9NOqzP5X9EZeDi2wdOgNJR8BRIhl
4wu5SNmO4heMGQqJ3la8IsqFf7I5ioWAVaCFLkzmvnYHLDVTsE7QUKzZ82s1NAPv
NOlHIWHRfuoEeJribcAmIICLuZkHBkPYGNaSI+pRGGWBicVEnYq4IwGHMTwN5a5R
gQThVxfn0NKhGWCpwgudBaiOZmCkfoi2IQZfy598KLcDdc6aJaAkQjisp+Hq1FWk
bfPlmxZwlzcxmgsCmUbUmr7rJQ8dHLZAd3XvsPURoHtt2ZkcaPrZilPf3pE7lCNM
+eMzLKOhOkahv65U3BcIxaySikHB7Z1qbmbLhfm1lr5qmYx5jNKDQuXuhXt2Jbjb
fajWH5dxc/XxoukLfIZvaMgdzEPvacOngih/JhGNIHcjbMihkODEQAqJ1Xgay16C
kNefPjm77AwSln7rCYKIlh+1Lv8xhu+LkIV/WV/UxnzSMEltaOKiMzwXUje+6JCb
4Zt+dLMPBuEDFVBRIgI7vni8cK3U2AwuBEuP/JIn5zaPEa6w/g1GgPqQdQBoCffV
CIYgWt0/hTI5xW8cLjhUDzx3/N53LBd6VbfNgeksg90SHXnYBspQQQJc7G7E8zpQ
U7tIqNAws/BeBTNjXqsXb64t49IdxCF0MY/kXA56RADyA4TrsAc3kwJlLQrMs35u
lp2hJZ7PM313uEsfMDJ6cLZzeCJvFYdw5eAaRPM+ieSQdKWg+IpJPU2XCJv//6Wy
FB2FrEGT33Le+uxD1FdKf24BBKQm+0Ypi4rgYj1QrTEykZPdrZy5tOLm3oq2v9q3
1rAANsZs3irw3xW68ItPfGUCAo8ClnR222zuabxGqMvbZX8hKOkttkl+ExZc6eXf
+D/GKV+RrdGKzmWOW6nMmRh4T+gWammB2T/mGHbw9FRRSzeDN+5fMiWqTEBCe9i6
qU2hX7kzgQo5stqYgwH5u7dPBJarGhbJoq7KxbHdrb9Jt3lWTIMPrCOL7nbA5rLh
QyVBTrpLIQcQKYWToUo+Wm7oznv8xwvHwAxB1P21Mo31+JW2KeX2jzc+zMrn1ksY
g3Shi1JWM/yBookS4p8IFJLVTiz0QJMg3vkvGJ8wQUSJYWiyAPUmnLayFdq3tWGe
31GgSTNgpbh0SPUwrPKhGGecrR21y0/ydlzTqBlOCLy06irhEjAd41pSnCJAcd7F
i4x2knv9xhfU/FtEI7ApMvhhbI5Ao+eNLM5Y17NukxTrL4w73JePVi6VgUruu2Fb
EWnVsaf7eQIbApX7Z06F2Y/mD70jFmPn01v4ngRfOdy2/Lk0oF/E6nx8QTpPBgjy
urUEHrvurdy6pgZp3Y3IMFP4HE56HhE89886IodBZumAmC5OoF3U7RhO5Y3mPPx4
g3r0yMGTxdnBzFRqazvdjkC4VRUnCH1XFGI0gBnRnbpLDEehjJO/Pa8mBhqX+OgZ
fbtwsSM0n+zQ7lM6+zHeF7+PpDHgvK87bKL/hnZBSCULXJ2ZTkheJx54ZsGYehPG
evEU3FvTlOWhdkHiG05/75cCrUuCIokA79VPfTjiJCm0eH2ivooaT4zV7wPyPqLA
KxCKhWADzrGVszO1JCloWajXqxFjUGH0ZkOD4kgkLvDoxzjDxtQz/x42tqjhFb5Z
n80lcal2khG8hDJbAxUUKRvigJBwK1Ga0v8v0iuy7UTRV7Nji/amcATt2vezSsjh
2aP3BonFknNjtExGE1fDzQVKGWln23B1fqzydVIC+SYkUNx8zx3+3hu6XdjrXdYA
lBUEY+ITf/wdrx+HvWcnWSTEYruI887YWal5N8AsqqoMSBtzrA/uZu/F/koTmTmt
EwSUQt9bgqIMH7M2SdqTdQx4JrxWhMGuZUCvD4XZ4vqCCPjzKhtxhGDS3Q0B0DGf
EjPfJBbLzm9DlvKWZob+jHXOCuvA68bLMRKml71AgwiBP0s5KpaBarm8RVyILq5a
ZZXSZ5leIpeic5X7laD75ABt8W2Y8xgnsrM2wQ+KvJGLVCICTi7CCCZhzS9/HOlF
0WOmpxu54kEbP+/hKwtlEzP9Ewx+/2TrQqcmBQEB1OjqbAPI6qTQ6KshTYSn1m4C
iBFXPjsQ+qIHEbgS65rMsPLOvzo1J+BlGA16PaIHKTFLSkPEeTh3ljXAqDFpjnQb
VxhEON6X2FvWV+U5OqNnWw9CEn+fthl2I3bGmhySWIoTqETLcPpfGcLDMeVKvbiA
3BTLJzVZMqrc1Wx7YUNoQ4IGiA2CEgwTQpztA408lvw229IqtKcXccrrQlW5jH5b
sr2RQtd+/ED0HoI143WJCSifuofxRlckKz6igRg2CAqtzBSGgAlGOiO9FiOcqEhh
BqLGa7nvvkC5BthB+cO1XVDub/u8su2SlXdqqvCm6ARHgkEf59+VGHgaBuuLqY0E
CRSfgVyQFRTRvi8F84GLHXJI+VVe4nKsY0HC8rx5yB6JB7nZaEI2C4UxCv/iXSgu
Rcv415O/F/S1AGYmHtUFXcmQm4B+4ZZvfTjxaZQImzm2M/XrXlVbP+ElqxUF1CDK
vStZkGIHBeA6DI0IIYqiQ3qtVzkL+gWvXygyONIGF+7NLjgZdmuHhQC36fQBmrx7
KF+/fP+iOxUp0T5eF9KDGVPfp7UEUww8sJvzORrLuvv99NeSbzSlrNjgmh9FDtGR
u7kIReWz3WxTMERVYj4+WvMos3z6Zrz4YtPOMNgtfk2uOE5+lZozeW7p7zC8vDex
ecfJv0GfNq2oPyc+HoA+HEc4ESkYv2y1Z8tVx9F8nYgJs9VZ5pHqNBpZZKiGGOmf
OXriHxoFpPODwjdVaJpl6FaxiLZQgG3yAyGC8z5LH/sOGDlALOFva6U1dNtz+Ad+
Tz6p+V3JQupMoE8eTtyRDIp+mh9VZmjYtopv01HZJL2p4fJquAdCY+euXEGONd5C
HzniDEl6ALF2g+5d5jAuqhijlZH8vWWxnIVVhloDs+XsHEGVlqZGBkQQvMrDapLZ
Vam0+hB2DiT6zMUOR+zCJP4zbaWwMsiJNaTUUuQhqAy7cfotYpbG12TPWqL0bRHF
hrVlhDCEPui8s+HYk9HtwA9LNZHWB/sRBMfdtG2m5W9CIpVw2YQLxn8rt+L/Lbf7
FiyEKWMpVSVcVtWj2zF0LxLcUoKaiTurD7SOr77MVwVAq32H7Nb8/UIbxG03QgnJ
7NszGDIDWeCE7volc/5eVk/0kX6mLcggwrbhPlWZDtFOHDa4OdoXeBQV2UuXfQav
fbsh81eyvxo7WHTKppsDsWgyRasKjdFezY5j8PPk/uczcbMum6/sXyVtXj0ZUhQx
xuACgjQv1SGVtv1mtMJW/Y/Gw0YGafEPxgY9ZtiNkkLO7wHAhf0WS1o63IUrglnq
8bvEaV0TjRAN1qJSmn0Pw2IDRBHOskEAZtxZrXsvXva2OnhF8HvC6wdRCwHgbhwf
cz+Ke7cYronPsFOEsm53AiT+iZjboKMC+cVWcymrvQMY7Ecd8hWoQnB7Xu8qz3Ah
fzTyheMUTI5lL2P172RYZpbKeNfwiEwsFtL30lM018fhp4C+bnBRDK2P0CHgCum+
6Rr/dGGpyrrNqWeOpXECxObf52tMNiFHp3RzsLVc1Avs07DVmKjkQNV73pzbuadj
vbJxOkogyvbB3WsdKTNtNR+3ZUCefyHVOrfJ96d+XuQqyViOlUacMtbQE83SEpi3
isfDcuCP79DdK+xvKqCMbhzinqWszjY1X6sRPm2/Sj6GyHvoPLaETRZ95msjWEhn
CpTo99XWDsCGvGvE5I+XBnWZoNSOJF3Cuyw2gQUQ9VGGSIvsc65CJmI8WWz/pqhn
RjM5YXzXmaTyWFQ6B5aSftnk9X52jTecKLhvqFLAEzOO3dHWdm0f6ffIK95vICx+
Pdh/pcVVb+mBNae67TNs29QGuD9cmHkymaFWtQNpWVhu79oXgqKnMk4PDTAHXq2U
XHFl82sLjaiMKcsyjgf3kOMXixEAR4NVcQh9UY3icalIpowWHgCi4IOETL7mfs1A
wyVX4myjOeQeUoRmXOu4ed/b7sRRSGclW077D6GktGBnQxB+kC3hOF2iyCqazmz6
qYWtB0TDb3Vk/lGIKRD6ZPZClkpNdT7L+EgymlLwhzQ1hhBAByrqULMxPuFwjuRg
1PZfTVJhgfA379dkhkkOdlcxBJ/zEAw4K6g8pkq/dwxo+fc2cfydh/8iCqgY+4RM
70sRmKSmPQSdXMDovR+zQ+OgLQnOikdzOrSvRBLG00bxrvK1HjMrRMrXMk6OEaFi
6xMWEnppNuhKTNdbjjR8IIMGOM4n9STKjO2psHrHb27xwGzXPNkN6rLm54q1wBAN
cQt/pOUfGGzeR2A+6gDLHfLX5og5M1AqAmbd98drORd25kuvhA02UZseeMStQ3s7
jY5MfCqpn0LH89Y2mwrQrJd/QS4xjq5SrzCZGCKb/s7TzYwIsmkriFyr5F6xfHsw
OpRfwkCYShibwCD1cb+C2uPTRFjVF4GGzsHsabwloERITh3DCMwfFGpghjMYyCdx
f3ml4r0/ZP7YVkoCNd3m94z9UCPCsCXZb+RDUQh+YFPB1nAAeGJI1q7OPTBM5xbT
DWDFOMrVFuVWe7EbFFL9ql5ZRckPhJj/Ho0a/7IkYXUC9H+WAi3i04XdbrX5FLqH
LTciaYURmKbhlWBFduC7SFcHSTq7Jit0PhtkSazPDc4IUO1+K/pD7P4PWiJWr6Xt
nJ7nxlNSBjykmkDyqhHSU9bo1PQZw8P2QVp4FCjLpq4W5034qp9IRnua6U9NBclO
lKfGRibEzURXictIGynZKPUPKo2VBcK/qUfa0Dh95ZUcgwhMiJCjXIl6XDdEyl/W
xP/4oYPKAb01qQrFCx+2pXLf/fNeiiNOsnsVMsqCBWZgH3B87sifgsWMqZagxFrz
8e9AM3lL6iWct9fcz8Tcz7vV2399Y8DQZou1rAyfUP8xBpYS8B6TDNbBnQpCkf4h
2CuFZ4yrkK/KaISlS3lsHGI6V84OQqnWRSV/M2opRKiDxbKFjD10TMe/olQNAjt3
ErDG7K8fPmHHL00ujv0XVKItyj3hvlOmERuxQNP7gi3XWD0MLGMjNybc2lbtejo7
Jea0Bp7btvvrTmJdfcRKvSFRhh6RRVEqzqFciewT3RCCTUr1Ug00H0E65jz1Z+rO
5IcHSwrrde4qY7cCmA74OWhIc5tPcdS0kiLHScT/s/x/KdQTHWuTyaNHTOlWza/f
2/Ex3XPiDtJrE4gQUvobaQGqqhY1Vuh4zOc5AlZo7bRWI/JCuMp/pfthqg3PAYcV
Upl09QKmqW8OvoY9LR+B3N3jTv0piRTOA7CuwhwUjt798Nr5bkgfKIx51xZGIrxr
oQeam1nfxwo8fj2bxSaQCXQ6nxpeWp3GL6GMfdXsZHf7pMa3Gxzd6Em9f6ffTnMK
qvukzyTwYVkIpu/NulNopGfEfxQQhfY1XWSqIFjQ0o+mkNQo+RGcrbIDI41m7CwA
Ae8TRRmRyEc3FzNFTSGMsIpibPTCdlDMtDCFMDjxA7bNU762a+mQu3oPJgemSOua
siDfYjdKdI06vASsT/63WjIbRmngrZ99Abw97iPscqnJXckjlVj0+vheQlkO1A8A
3sSKovoxBF1I0I7h/1knIT53ustUZOLuAlHt5M47ekf0ODAzFjqVPT+7+/B8D9ZP
9HMqj6sO5P23jyKOfd5IKkca2qwmoyklQDsDtdE2kGxmsko6XYD7cDLDc56Tl17p
sufB98ctVCFn4g7HCT4rx31urW8EzvzTAsatJlyaGmBFebqqValAiGJSC7HZGBxJ
VV661syusZTPhbr2B3I1k0fd3cljjVTAOSxQ3zUO6yxDi+8BGiMehuVI0yiZvsml
hrcu/1N9ZbO2Nl6yWyr7SB/efrMjhrDfKkSNESITRwNvfyE9Drxs2KtFFxEyChNi
p4fmx8iGFCceIr6Ul0AFpPDg2tf1shgHh63g89C5ovE/AAVYJvwcNxvDHlZpixRX
kCTm3XQJMIx9Je18DGvLMF+fyfOxQbicE3IpBy1vYQzxL/YyHcnhM7uPidlQWS/z
o8dHEYsfb3kOmNAF1zmZukz9kzbQv7GwHJQN9O31XvagZ/gKZVbH0RHapvw2k/Qw
O8ZZ1WDvArdliVMhpbUl9SR7WjkcYSiE4O2tpMKwmfFAekH2R51duYRfd/u+Kx9E
lQAvMPRQFpwpX510dqSCn+qpPZcqiNdr6VnPKPt3e9z9JeFw73fPg8+oEqziQlqf
XSmVCzWuSB6te0ZxdvaW7gmevdHd4UaItixXSAzeCHvPNHZ0+XUnrsTNUJMFzf+a
OVbEKFWJC9ALVFX1SV/b//gMGlxyFEo2iXdc2yZ1fSkag1HiIfjAXX9kbjMVXAAt
J7qNI9hA9wcwlJ8FIaV7x9LcKiVdDUP41o7SVcY+qIbGY8zGJCLNxORTvu8UagLd
629aScErjkgjJdgZqP+h4ekn+AixxklC5Ty9j8sAcpL5p5YJCTmENdvCLcYjnnHO
/HzlTFYwfFpB9J+zixCuMyr9xGYxmH3KIk7NvP2C/j/NgoC8gEjw5a775yIVGCnF
tko4I/l252CQ4engxEgC2LbVTtpkiPaSQG3YKTUjEe0++QowTpnzi0TxxJRR2enM
yAef/7JVCTr+0oqRHdylqvEA56/6bDj05KCMz5OwbHk7AIHg8jPNnn6sXiC0j87Q
fFn6Iv1uO2skygWh6MOHQtefQ0vZHKUaXY/HmRt07fHiSwa6tz7eVk9L/b5z1c+0
NMkpKkUjLHlIJ0DcR9HtzsCq7Kk7sVeKwffSfDZWlAKiPShcPpkdmZBi7Mn+yU/a
sPYhtcE0oLqLAI1JKZSYsk3hc7FMpVDnhbYm/mNyT7rPmUoWi/FOzdTaPG9Q/7Et
1Y2hXMNkTuk1O/VOSkXo9tYANaY5FqcLqF130QJCeM/SB2qYbM4MUh+7z+Z0tpb7
skIopPqqlEsVbDCv6rd0oyWZ9S9581wU6KOWPyG/9abiGwFjk12BvWikudtLOkgT
SW395vZQ58o6Nio8QVHjA+Ope3d6w4qf6oSnK0EUP3a2DrQx912wMvzXl5qVCnw1
SdYwHxybpNiSBXcu7GkCBnALav3SHJHgY1Buc5xksBcSaXRquU+VUUtHpMyBNU0n
b/mR9AMWsbj26qByDv22ZIlOJ5oh781e0zijmx7EiuxKWh/psLiWbZr44HOmKVKe
ge9gwkLERr8Gog0VfaAmxfdFnHV2eVMReVe0fzbVQ7Ox5ENo4MWzrhOcoT6Ij+ks
7VRxEBXqZpJtLUDpwsjzgDDYiQg2FjKODbx+O3AifVrtSJC+1E/nATFJgDk2VVSo
tGtxLF+eqwu2x5wLt4KjEypiY9iObknCZzykrTvQ6lL/m9Lq8nVYUqo0uWHsDPIX
ZpOtttPVeByN1P2tgcBPiHdJCElVPzj3Ju12kobiKXABZ7BvI7c67lPvKI0ewCe9
/nSJy5+7vJT7ox4tZyK1Ydz/UJtkulFKju4dfFmj1I9SoDCn8kJbaCdADQ28K0iG
R3zteaZpgmFs3sAAlOHXjdwxUSYEq4HMHyMzJikrYMFAHvAKoob9XKaREV+RTh63
89GXvnKArnBmJH9gMKvp/QKx05skReIiGSoLrr1oY8kmPOs/BmIA3d7lOaz0dmF+
apAa0dhZ0r9EQHOOjcsHu31CFjIJOAarejvVpQqIumaseP2NCc+vqHgA/lXo8LY9
aoTpj9BCp/LzsBHyBU19t3AUuVT6E0j3s8dWeDTufNOfs1ZiZWANgqjaV3o0Rr7V
6+EX1pfBahuXPirfizs7z1Fl+GX5L7qbGDG0YjIVZVc3UHIZbiacoap+YDrNZPf9
gjqPQ/DIpyjvnMtMAUBGQmrMfTnG3S6/JqoFKZT7jQbaPWs222jpE3/RKGnX9AH8
O2T0YGAgQpS5fR64PyFu442xph/5/+cP7ihKKxgP3hzHJMEw0IuiojwEoIXHHlWF
vhcXRcWNxiHB+Nda/3ZFXteOIdvFCpGeUlTZvJ9bascOfZVm2nE2Lo71NK5qK4ux
kbOm8rs/PETRtkeRazWvVAsZERfBhSitouJgbzd4sfPUpxSJkG9CcfhfdoF91YxE
h72Im1ULmqoWr44Qoa8gtlcxfDan7fdT7aY4dQEe2+oUUnt9xhbKrc95/C0dIU5q
q7IsTnXy36Xe/643a3Zh8pRc4ClF5hTFI/n24ioO3VbK7kE7bTRlDOrOMCtlSXJ2
DE9ZpaMtPcQpSeg5F4LQHljHpM9lQmGIYUWGRs2qxeHbknh/KW9NhvYuLHUX2jsC
ucklkrgpnPqMacLZQKpnf23yAiI5loK/37W8ywnXd/+dMW8L36nouT/DY5+wZZvM
YRYfEo9G1yhTd4+5TL0Pnd+TYRlRXELqc9SLYGMrX4Zc4if6WI8Ad+PM+8i8pEFa
WACpaoa1ve+iaTqXtFIZZgyFAjMxAFXOWLLx01vXUzSByERWkZbupkzmDliIrZSW
FwPRuLd/sOeJZQw4lw0Xl9e1eN2+bXnJ9CzG/jdxUDiwnBvpEKWTkWYliiPdbpJ6
P6xU4vq51XA6O1jxSEXl74dvQjzfqbIf17hWf11IR6GaiPV2BCplawAmsqiZAtJ5
MU3FHeGuNLL0Q1mXfVLP9wBbEkh2sd/Y9Cq97k+gxXmUfBG4RHzCAAAW5n2GMLeE
ORglwdXahSNWHTAoIHJpy0Jy1owziV8GS3Ze0+LKGlpLrKhYLAbKxUTIwnfCV2SS
Sfwr7XcL0x2qjdoeoeY9N7IawFfddLn8PHlJbY4Dw1ZgqM/yYAguIUQlRESdwKEc
d05SavyAry5oOr5zbvtdySOlVMRp+Nrg+lJ/uH1ufydhtpqzXxIlZaEF0jLg4AWR
o1A19F52UsnDAehsjRHeOhRyUOWBIu2QhJMjSRzicwJv/kSmbXGVrOQIW5DqKbPY
w+tZYtp8tIq6BhJz8epTADOfSqRT24vLXw0QqMpOM8fY8xUm4MrAvwA9EvFRUX+/
2C4/4FOtpKI1Tpyh67zRFikOEpATe//Af4Rr6J5vwTlC+L46bTm9nGfhoT34heG8
4upl7rgb2ESoYEs5Q374UO0TH1SrFBVppLSQb5pcxHNpuhv1UzNfcyRlhu5yHcgE
OZdPWf3mzOAA93Cjw/E8pWqzTzkELC7ICE/eIdHpPJx1XNsWxQ5tfSSvI6vx//N5
xYqVmr6RT4fmGVefJMKFKjjcApY0So/u598kItThrdX7Vt7JDELZpSZ2m//9qcce
qVkpEbXTfLIiDcRcQhYdsTX8Np5Wh186TkfmUgee1LxqMg1xurzzzL6zKzgNrFZ7
zRdPrnVJzldizoQEKVZV4EUGTjFjj/uQT7PH0YBJa/QEGqRK1vXFZDy/jJJIAoeP
jT2mgNa20XOmaC+wvmlYAX51FiAjBPN+lEUvcAjxZD3lcrO5zzQ0wKIuRnT29jJu
re0KA0gkTmWIDMyoQzH1Q1D2pGA01f3U7F0/YFRxtwvfiOH+8q/ouv8je0X50Y6l
Dj6rECCFosaXWqbRGOJnQWoyeShG7mHnIOXtRoVkXNM0wvqgDpKF3r9AjBroAf71
NUU5LfptIrixsWywNsixIiR+rqvtYJvN95cuwPiIhVDHV3/T0kovxB+CY9zRrdZ9
QlnMyG0O0Mst+MCQRdX8YNFLaX+9EsbWmqEYHOXHjlpbtZzJcHIbehkYTNZvdpc6
RRvtwdiIh1yKarklr/xntv8SR3d/ahq3X2+/CSRjKzBBE/BOXUfiifwKrRWVYAAl
jSKBfUmCslfnxtA4VQHnLKuelbw+YdAeG4D9EodmFjVdqJVNkNCBuX6sUX4QgpMz
p7uOzJRV7FsManORM2EzpqT8itCGdL8mF45j1/c/Y6SucN+5NPJp6X4bBoWd96Fx
KH9qlr/Kl6vue1Sn9zHSjSlfu5E0DA4zWVTtbtyI88KVSbQ8ndhdtHtSPGv0yG+8
QIHxuUaNhE1EnpkCQyUjWJ7csUUmQmFApy6PxG9D+fZUtDJkskYR+u+E2IxvO+tZ
AOo6qpiTznEYJQqx7vDVID7cVA8woG9gOyRCOkF1Ew4FVz4zRVgTDuEEZhqeKQNI
Ob6oJNpoFIFmkAmWydjYXXk26ioLtmTFBwpvw8CeU0CdjpHfvRs64b9paVU7mkVo
thAeguv/D4FBNUlTyPWVakl5HcnL1Fpv5QeKhGfAPf23eIXQxVOZvFYX+48/VtAG
3cIFtKbO8BvKv0HWU5yDsrxsmchaNNVaDMghiV3anLYes+/I+fGbA2H432aspnN0
b6856DUpOlO0CXiI5CUn3HwBsYBYOo36Li6J+z+0ymofLdU6MSuC5pS25D0YII0N
LD3iSvnUcQSMQPKTkoYXoTFppATu2tArdlxF1kSiRxx6hPiuFtn7/Lu8fEUEaspj
UVTgr7+eyswlvMDWnI+eh1kPcJbadLTo1LkP7XpZoQXE9HeJkEyJd71oJlCYZua3
c0hveO3epMQS6n/2C9+SabDaWoLoCvJFOxo6EeBxTrkuCQslHut2pfOXuT2Lx6md
5pLp2AyCXAAb0LRALONzeBhkPC6N2T7d8ZTLbM0af0PSQdIS73ntq5ngRy0DgQQq
80cF+wffEpJLX0cH3NiDRr06t2F0WnenejtyiI8zD70eqlk2/zVNhsZWsb7hmVVU
3js+d6zDb5eNT3EjR1bUEOtEVU086+OXH+TrwcbvrkTOBOK36+VaSQaMTQpR7v2D
z0CNzAEFNiqxYDYQ6w++JkGO2kqZEFUd/VeD89ai2Z+iyCCeoWodiIFjRIk4MnLw
fp9FSX+X2Ttvt+ln/eAdkJztOPC4pYUjtCGNcg8/gX0C2CwRUjqerQyhqVtvLUaC
5gvFVX9dRE/VcAUW/TyVNxMKlWVdSME587gfBYll5Gya6N2B7vqqEyYU7/Wlard5
lHRovZkAWbBdrm28aWQWb3YcKKfQfUyqxw+CCd2DsqulWNU7vwNkaDez9gupxiif
EQnHLOpgG1/sAPps4/vNzdbvQ9ffXdJXmY4v9Grk+D3g9C7nkZs61SzJLdaZy7Hm
WgGQ/vzsTA6Ae9m6E9YwDcE5zcjj42UvF1vDvRkVwz8d4SWfNcOBWCrZMGmwOaA5
HhzKiqQTV4Bmh7v+Ozg6cGNmVbfhFNI2KvEAQXu6Szl5PQc6GzoPOVl9dAz6dPFv
SXgV632qkqSYH8+DpfM2BEB63jla2TnGSrEyLPJAwSgwIl2zK/l1qXZY126X7w1w
lX4AFheiCOcM63azEnive/S2xZy1/yHNJOvSVVTwggywL49syI+hvtrbiXVdhg43
bAFhasdYcHMotCkoCqDZUovmabNxEGkj99/0AUyVwJxaTVDZF5UPoMqseVH0h3p2
tHGTdQVAha5ibdE9TxTzf9y9ZRwwnKwlwSUfH0FRemyhWFtaiphhH7qrYZGe+3oE
5v2SfM6eZLfHdDMmd8nOLYHvQemjsS4Fl3Ff4BZYNMMeTq3hi62s5H5sMkK0rhVD
xNg126yqFYy3z+fxS0NBSjELaHjNQmxWqPbbKzGIW1vyy4V8MgJVMaNaGRe5wdp2
YSHT2klGppIk6IKPdjOkWMzN76XJVuPte6DhZ6+m3g6mp7DfQW6EYWOwDjJIZWGD
AbqnCUrpmDWkYNivHKI33tNGZu7C3Pcymc+R5WWQ80SvTEvC+anjSX5sIveWDRIP
Cb8477ZritsadNEblwMjLAvt564noQJloOJJKonZN4Bgib3CJncG31X2u+45T8up
BqjN8aFbm1NHkha5Iy92hrbrBuOdLIAoIE5mlIXbqzO4prt3puLx5mi9DZs4MNsK
0BNf9+HcmCxo5D3O5QyyxY7RqmQiluVoDbcCTLfFGzrunv0d/2FVEmzrFK/h4S35
TQcA+ucVWNJwize3vJukqFaR2SXCtX90YlVEEKysfISb4Y0HuwE9CSJQ8iqmE0Bn
jSUqyf6iQNKbY1OKPK1typ9keGCLKed9NuyXqhsqjvGGUpH6IznMn/SpMBdA6hhD
ZajyeX7spu32gHyBPi4F8rWIAFlYJaFBE0l4ORs/8aHjMLRTxSwhIS9BRh5yrgiJ
3X/g/Szd1IaNZZsRZr5sAk00m9dCqMYvvAWlUmx8348VPmSLY4tWaHDYuVKFTGLP
T7Xk1EjZAUrGT+F2UzBUEAsedg7nIDqMDRftkynW5NLCJLZkoFMdp6AzGE++Z7jY
jN2UhT6GXvQvQTJyGnmE6sqkKlnAitlIDgST6L+gyWC15dbQN4uMN3oe8qapCHbS
4Rv9xogCXmPxt7VWtCGmcE7u/3KAgNRE9tu9QA/jNmEACmZiEZ8E37yrXJwlpyXl
jKPSTSCyHSIJwNfKrSHQ5hnfoisZRG9+LE1MPLPr2CIxSW+vw00oloJ2eo8LSv31
4krETszESAEbpuhfxpupEzw+B2cTT9VDxm2xtReFakS1GogK6lIOYwDUv2wUxbD6
s51Z5yR2xmk8ZGMhyhsCbqEjEejDyJZgvm74pxO6RfSdH5Kv37Pd+61xD4/QL8N6
tqiwdZ8Kywm42r9ATNcGwYrG+bHtbt7hHDTqB7goGqrH7GnlVnMwAmgXBDUJqSmn
cjy+8o1wH+MJxwyP2AwFNfH1cl9kWMgkMmB1QgQNOLqrT5etYMFsKslawTS1Qij7
lFrfllQeRiWxp5VFDfNtLmb0zP7sAe/rsyaOLgi1siI4co4Zme8keGByaax6Wryc
mGw/WLE4pAkrhYP46hHauoG8SuVOnZQ/Hlms61rKpvkYmr2JbHhxRjsR3Y4UUmP8
CWR0cXUCzfOickEqDL+ZJ/d1+5CGUam7BAvuWcg+2xAB1mEfG7Y69sUJhMDNz+NL
/vPktgmexy5Ynwer85dQ3NIAVW+1SkUjOZupe9GAhLOcS425Z70+ouK5izbl/uB+
PqqCUoVFuBiQOiUcRfm6aNL2J6imZYvAOauu+tpfxWI2TWlMqqY3viI0jJZXLP1I
hNjpw8Qa5VXAjBBU9ZU5g/bZW3bt12QGiZprjG453Do+O+cZheP6BKHBPqgmFCIY
rnkvfgKx3qEgZDdYFQWdqWKUpqeKeeyw4RlB0SMlV92Drfc34pYGqDgCDY6Bu3EZ
uZ3X0yIeeiEgiCBqwtGcPzGEGMqJAovNjmIIv2b00RSIbZOxl4NQH6a3mDzmx1OE
+u1r2k6UsMBGPdQBZrV5Xl3/udgoBXaJkQBDt+wfCL578L2cQCxEvTHmD1vdTti2
SgKaVIsOALz3/Ld/Jj7Y5dMFHCdoRDyCBXdOjdgJzAh2SpXtN859ZNSBCA0jy16Y
KFsK1dnGvP1ZIvUPXhg1WaknaJqp5l1goLJ4IwaJ5WHVVyPCAdQmObXB96i8Y2az
dUZbXs24IXSgw53JDJi7ajjDRuHJaCQtMqnL/o1Igx0duwWSEDrHv4YmPq4w6B4T
9I1Vs+qNY/RqAOheCYRag6UZJFR4HELXZUQKC5IPFSUYkP30AO2InrLN5zAsW20W
jxwMRpsiHPJ/Qt5eDtU69n5MqCIL1jzDU64gn08AZOqvX3A9yNv3FGB71bRQp6ek
hO/d+Gr7pO2FImmIjmJozCQlCp8veWoIePYEX7NUwRMJ+MaPrWM13PpnOx4AprHg
i3yXlFOukm1wWFWpAsjCb8sMnTiazvWX0g7nZIpxYU8XUfXWFuxLZ+bjZnJyyFA4
fix6O0uFkDbWZEs8bbV711OJxz9mz2Ih3UGhrBjCLN5WpC18PceJfHC5JEO0fvki
3QtqbWm27dWKdju0kPm44p5qSrXs7kbne9QkWNnZiSxIYOiggw3IQZtkGZZT2nHU
mLP4qzJGVNxXG/M9M0SFvv4hLIwh6TMyoQesTTrJ0cgxYbAWWkmTQIky5v+a0N5j
BwDfF3eOHWd2SNgF3DRTd1DG29qzuLxdWLOOiWOdEY8vZY/nsgyvyMJ+KA5AODnJ
eYYjWWpehMGqP0nBbNsdLWY9sBtCWNSgm+haQNzunqa8ezxqykNGFEMRYBkK/QuG
UyF/NPB3jt9YaaxknyGRq0aPZVC/3wRnXQZNdLhbw7PxEx+M77ggYoz4COkZwzWl
0rWxdERlpDbQDd79fYenr7hMJeMo+xpPfnaV4YpHBoGKRXCOET9u4iTvw29sXQqe
gw7WNYWTqEzPEFR+1GTlEe3wR/AbO0sFGhKb7ZbFT1C5yBs4V/ys/a4SF2+VSxRx
+zWFsTiyZaxLPkf3TkvIRNQwjXDFyuPwOeFz7A7MxGJPwnOAwUgvvfBfr3v5XgT6
wMpiAG4fLMzID/xA5F2sJfK6lpU8gH4J1NdsxH5/KoQIN+FbTHUvDEn80YordPzW
MIsAPe+OeYPbq3Y6RtJPtp9SuAZBT0hoSj42g1erPYBKAtsAyfq1j2EBz9QuEdWE
K6pcUjGeFMXKr2D9lj+i0vwgPTD9E/fkGba1KqqDxOr/Bbc7xiChdwV8OnWFVtLc
dvnC4/SyFpZefMF56R0TxAK1MvnZC23f9ThEK1YIyjWSt5jMHmbeSu0neaotIFS9
8oN85JjyyPfvGEThQT88FsReaaJlY421wk1O5eXzupgauApwNYmASdjCSR9kUliE
iXnO1ynqac5RjTQ6DoS4m5ylheNmO9YnMCeXdQX5LbdGmWzy5Y5Q7FxK36St/4b9
jX2YxXlBMlwbN3bBE1P2Ho4V97P9Wcl3M7iU2sEfKyyppaVnO4jVDOH5WuCH8imn
a4ibluNjGrdQ1sVncyKxuUDFAvFExuQtbHxyfgkBl0G3McZztSgtvVsvmQTyilmt
QLYnSilRol0Sz6Qa9fcCv7WRASpcJCReE7ZR29sswIlcYC4YGbw/fJ+FstR5xCtA
p6j1egDOi2tIL8VWnDcHnSJopUdqI9uFFCauZ3m55nHrupzYIZ+nY3lwxYDMxI50
jXXbYfMGFcGQZx2W4n2JuEk73m5u58CrUncW6UxtJ/0005k/fR9mtVqRmFq8aBi4
tXHbCj1N6PfPhG9CnhIloLvUpyLrw6N+/0UBFkDeBsCnJh8kgbXVQ5APWQXlOsmr
XGOatxEue9JdGDO3iLyW4Iot04nHE5dsyCrYwItTN/XU/gCye+qOfbmYUoc0De9V
bchf+xkt8JZQghtPRo17y8BB5JjMR6uBSfcM/a4JX1vGlizAnLJBichspoR2OxvT
9s3L/nkIq/q76qoVA6tOWlB7auh76/JzDMw7Uk8ckDgFK/Wg4viQ7F0zwnFyWydA
/IK8C+7lix1f0CBmTZVzfO3tLvOF/ocvim3GpnZhfTQyrJMGMBK7NK905FhG1WF0
VzbZFOSLc1v/1t7mUfP98w8+PGSircon06pzM0IDeGc/waN8lTsO8+45QXbK+Jf3
pJLL9Ur8UwgIbnACFDUPe3FdJCPVKbtN+obD+3tLID0SF04Jk4Z8gHFizwlLRN/Y
CuZ3YK7LP4TOIP2FZJyQBHVoqgarPviMrteVqpBhz79Axag3Te7cyFNmpbpSRuIr
Xs/haovUh5C4VXF9sJ7iueinfvlDc+/KBOhLB43sSM7Qqz4v/eMRWzNR4tU+Gb1M
sDFEM8JEvWXOByG4DhF9JYmAembxGB+LUSb0X7eq4w9rfdvxL6s9aBzgJ/4mX9XD
OXQHaJsYDMh8Hj1Q3i90I6B3NXTC1nIgqiraMdXRYHEsOwvmxlskExadOPMtzZyl
ssVLPUUhNFco8upDMx4/WVV5ScrJWdaGs3APgpMEYrU9LW6X46pC6ALwTi7LAq5E
TpmlfFyocPEr1qT+F37DvGW892aoN7+PczJIoDLr1vrpWPBHv6NwU22OSdbSOb7O
qYEBuQ3t2PSBO7XfL4BmJzvdRm9uWW5NmiaW4JJSiy45klK/XSCvcX5l+vIIm066
mO2BaWPFbMvF/8MrBdg89mXrIk4AfJg6NW/GZUGgpaba4Wuxbc2ozvUAWoFkksXJ
SyflTyADZAg+stWFFTAcbrVgYO1jzVr9hawwe10NHFJcUh3RhAAXc7VDzT3N+/Cx
pd1jtMInkEudf0R+d52z2Kuv74kvdQpj/R7/HAcsTyZk9TVJYp513nRmFMWLLHlU
GmYqA8Lb5LsuJU4XudPlQKptL8K9AjEk8LZpYEH5JFe28KI3G79hX8BRe124EVof
ie4J6f7SfXRtV6bkT0icKd6gPaw8uJwW0oC7+ofJkQLJRjIoLaqohpayqjjftMv/
jQ3yBlxZKyd4zvwyLYfkj9yQvK4Ri1rTWl05WjN4kjrYGvNBC3hZAkKCQAsQ3GiK
GPMCP7g9t5MAOv+Q349jJqzAlRTVrYuVNyCrbU1lVEZVJsmVDGMr8Ah/cVTB8cJZ
OeJABMrTp6iU8yUY83oMKFtdJa7KbmXhrJ14nYVznHPbVmq8BjvJbqDZPgtjTVZG
OkGxipTjkRQIGRfXQlyz9UN08UFMfNDL9bIX+WIIeAYaDK7O2FEzM0MEvQMnlp36
tki6I4ciE8zeNvC0ecenIs6a/rIu3jTw+6va481IequkJVH5/nTYJEWa6/PTW6U8
2EvMB3q87R8txDomjGWFr/kD67RA0YaGMhkweRkssm84u/l3W9RlS93cTfHVvnOa
Si8mQ321hU4SP26A4CnfgdUGHRo5PTul32FxjTt8p/seK99Hocn6SMQ25mLKGrl1
2Pu3qlBhsg5n/WE80EXZ4VeRLgl6FbDs9PeAy7SprwuqGE0S5MafCQGEqF8wXWeC
tbVnYZSE8oWJtuJW+/0/cDxI8LczCqFRYMLRCrS7+CpttmIZCZMe1jV20qVKXlJh
ufKV+sCwX6X/mY/GvQByEZsfomCfTM0kW99I/JOZIM2NCIRwgP/n3OC2PWt72hxF
h8AblhJ0YoQhloh+iHw8pASR/2s3ePoHtmKKepYTonvMGK4+OsTozoS6f/j8iXXG
UpEEo0uukxoxDT3x4XT7B9EchNKU9JJ7iR0NifxS3hJQW8rSJ435HnQIHA8Sl/Om
4hODU62BlfJtZnd8b3V8JYXWsRphfcwwjplSOxz6nn7YXsChWYfpkFjj+ZF2DCel
+32glu6XyIKjPCQP+pu6C4epqNvjhxgxddgxSN54Q87aCwrlTJatg9WvropDHDt8
4T4fihvRXYglq8ZiPKVlQ29q7rrXy3mpmVow1ursLDmJ4fbtLiJ2s0jiWBCG23XR
AqFvUyxhWAbJaZEXXAc/9xXhW4IsG/djrHMyQH5+iwy6r+zs0yBR038mglq5utvY
n8MgqEwafCukauRxn+71KF0hpAj0s0PsxnA2+xkFwz8ks/dTeg/TIdtFKJg2ZQfv
cnjJ15k4AL/Dc8TzPG6Q+Yj4g2gzPT0FmuzkGEQc+lTFNcvQli37/s4ki/20G4wV
YwMqf3+ofMUY1hZSU+e4x49oBZsMuPPcndg+8o+A7+PoX47iCzWyZGGpclBS+fyd
Kcd10DJ5HlW2MdEKt5HSl3SE27vEOBKZ05N36HlqwPNUOiPwdvYA2i5tJp9xQVBT
pOQiK0fXdMRTgqD0HnB5JqXa0BaVzO/FUziDImGB6/OCPlOyT4ZEkNlxko97XZmP
PGKjp5JeEzj5OjseOJU1jr7CmoVkpKL81DZTPOO0utPFu/Hhew9aENmZdk+eDiGJ
zkkOAZ+VMlmtCZWaZZNfZNZCLRqPh0NKUSZQrZoOSgzSMS1M++Vz4p5ruif1nvI5
OUN2h/BVdAH7MyylyKUy6Jc5LxIwjPbrfPsfLISAt1qmRJ8XKdurEZ5H+OEi54Rd
Xv1rPBPQJhMnSbTt9ifJsy/QLkp0Ro0lNN9VvofzLFua8ab2nEADIbs2EPb1oRvF
fBpMVFqBwe+p0oGUFd0NyqeYNlnM7w5RfR3WonttP0R5TnT6kZDciiswEVenYA3B
R+3xXXXkodQGUwC2U6JaLcj6odhu62Wazlu8EZ/zrCJ5pQ7gmmy6N7pa+sPB8zMc
n32yN2h9vr1u+0+v8Mx0TNfyAX4TM0VpuWx6Y/SK9fRz7z7LaskXdAO/bTedZ2bg
uIuJvRYKjiz3BmGqO187C/HD2v2YDMCZYLmFdsyrs0fioHwCIZ/E5cbV2sfgbhHn
U84iKeR5JsteDjU/vGubZWUQd9SE4s+1vhA2yjgY5tkvlqFtVSuHDUMfIwKuK9uV
wSWXEjshJ01ZAzI3bYn6z05P9g9Sxt0AymmhRC5z124phe98SrFamxESTsG9kYxO
sko0wLcJeGsu/ngONTtskxQ4x/kY0L/jvTXzG7QH7tgjNUCRXJyexcgvJeZyiOEh
UmJaX5XnoKKBUXhA8gl4ywGwRv+/jzmuKvJXjj+W0pwyEy6pK5rnq4Y9J2/uQYdL
GHJGUxWqzDPunWGOMxaHMFuSJQ2XapBOwGDB6qQqbbfw6jKPQ3g1I+N+YHRwrKsG
+ksSOPAa0YGabYEjZV1/r+bYnHcmqr2sF/BTEESa0+2vdrM/fNfGQBDf5nXG1kxC
J/4TjTdD1/PTii2p28sFl4s+hqYFCH2ZYrJVvHYjtN9xxwDz8Fv/ZrkMYVWEcATH
athC8Kx2KN0G8itHE2N6UEiDcEQDejUnbSGvMmuMDyJThNS6dsNGbkFdAQAP4G87
BWLrv3Nbei1r0y7HEbMX4nNPyFr79KM61/m8nI5M4ReyyR2AoV1SRqBGmYOUPZal
449OpIBLyvRB+pC09DUJ9xS9EREv8pKCfbEU2hrC1mySPF/cdTQ54giByZWvJi85
8MmyeAJ6FLCyT4kJk0Ib5fR61yKbRxUIwNAwx8i5ujx+mC0fEaYoNRH8i2OFuKjY
+1lP438pJGJd5xRNhQaS5Wkgxm1YLUvBYkdBHHTo+IHUnrfIEDWIe1UflVknkomp
+HYgQ5jR1bDW9aRzOj9nRbRnUb2lbDubROUfvVAKiNcIIZTbXA6nFdAv1BrWSBsK
P3nVKyaKEJKMuTjKFZFZ0xM54W8eN66e8aWVil5DfTcNPKfRiPuFg3cax2MkoLum
RK33qQgrcZoCxR3QbwMNks+yRRYhzA6traF/r5ONZmT4cJJKl0t5hefYRHMDU2/B
ZnkBa+pKU0ieFCEQXQ+03+QiSczM/CytEpE7Z+2WcnMtXuid5tMPFJP3CqC8G1S2
U5ZVynNYqnmBnxRSoxSCKAIxI8Mx+xceu0ayj9fxHoW8ZevkSgEM7Kjsc43HYJwy
kcCmhOU18wnLX3+i5gSVkM6zLFJnou13ltziZ22RR6CaDFiKyw+gq6W6F8yUKBXw
c7QxrrLeUwvpg4Gpq4lAWuSWN+QCByI4M5zmHwelYK/7Ra+pKe88dIFiAjvL7pEr
OR6vnBexzAgSwcnCBhdVQK3C7wp0WTz1n/u21F4IXmruitABNK1YBADfXMUTYJ9n
DFbWvAY2kbEq52pVhYyOxhs72YFpTxqzwr9buYpPsc2aGb+PUlXj2xKIzqfC8To+
anid3mmUWLhIHMzgiSsfCBXtw0ES989v7ZRwkPJvaaW+iPYQK35Cfeu1Hs44qY7r
3lydHRrNg2hLdViRQDklag7qwZMqyWiUliQXPuB348TanbBNykoXml352n+R//2s
Y3tX97ULW/Mu64EIluBtBqPGSsCYa33+2SuhAZ9XyuGRGvAjlz9QqpV5Dx5lYAlc
SV5XmwJmoi9KHAcE6XlbaYr3cjcgTQUgUm/uZ1vcUofbdqa9rmVb/x6h9H6ECBzS
oI+NDLsXwO+dMnOmJHxUNZw8vXGFEtIwBSrmXxmFIIIl5NM9yBWXBxNOmYRvXqs1
N5Ez9QIFVIjL1U8beWiHv3c/b/e7vMNhpCJzqlPE28XSggpTV4qpd37hDQESt6s6
/ba9wFGZwD0jz4oMpmWjLDJEh+OIftDkFWTQ74D5yob89SqkTPGnm1w5ocKEHKY1
3Dt/yos3eFGUJFFxNZdrR670ixZfrtvEf0UmIpnZm6qWbHu+wIkMMcsCuD4Kvf3l
XBnKbiqdzxOXm31zjMsWX/ZxWjlaz/fo7+I+myueNk4vAy5gvmXQHaRpGjSrtHtT
S81Wf/6fED6yd4zO+uoWqtNe6hNe92JUMl1Mb/kOWN+ukxMZt9gka6fBibSFn0I4
n1jjFm7HFEqN8i9Y3AUVJi3kndy9z4DiicUmumsW23tv8DdwNKqIsiQsne4huz2T
et1HdPCapXnvZ4a9lYPqgB3CQpdABhLidN8s23rPrnDf1daua2wCZMfORVh+Gs6M
JaUeTPXmBTvazPtW+U8l1PSLOqrr7sQ1025QcXbgeVakGx8BNbcUIbW4uTv7yR9g
80DsGMi5J7jjPuxO86bAjtKvQigrYIK5M7vVsAciMs1lL4C5PUksCl9Ltl00JiKA
cn86Sbse5nTCq/xtDAKbA76rTCDDfOxIz+Xs23XisyczzfasbtvLJu9eByziOKcI
d/x0EpJ3WrIPgtrb1oorJqODTgWRkyLNFzqQD9acYAQSOox5XcngCmXwBhy2A9+8
/ENdBPYrwHkoEFgHO07hSsJvD0A/iS8tz+SVOESUi4HL5WZ8yqRwrRmTIcEs56Vc
UDKdqXUeTKNSwqXc+4j2vIberd90sHJfPLkNDdPT/TXv/mnURb5RZQXUBSP0BZby
815x/8iX6EOlfiaPDl17rQz5PN2O70SSLaEZ2UW4z9xHeobaKQeDmC4oCzM2taak
E6OGaNOenU0h01Glqz9Rbr3qzxWA0r5XJyRFKvl7RBNew41tqis/QItjdOobN/Aj
p34FT+1TYOEnMwTO1gVFcUJv+5OS/R3C6oJDng1X/riKiFCjsybvkv7Rp9ONdMVm
ptoDOWYoPy61IU5OXPRO2f6pit2IT+6CfmqAe+RnvbM+HbcYkZ7yphcq9wvN8AFu
17P1OmnRZ6dLwPqMFCXC3u1lqOjDzq3AaPIogowu+6K68zmtKi3bW4H6Z/Pxkm0I
uFrYXh0bzFDCf/6dedZLblPQ0yultGtKWa6jNCLKC9/P3aA0g44nQbMdrcZ9eSd3
mSziULsHJ819LJNgc/VHuJAMMWl0r6n0MXAzShLh71Lx1llxUB+jZDRpo/l3bieN
gLnrXkCjxaeMKyf1rd/3WrpHbufegOeShh8tH6b8x0t8bMyEmspfiuHIxs52oLn1
m7JVCvRo8mh3gHzHNJgSImZPzQeR47vCUIRMxyLmFO9+dP5VO1pb+UWtbf0m4f8S
nR64C6jJXoLBdS1g4TjTicch8VxsHMWfjOZt6F2x+66M0UWpsLDQfuhddPr/A+Ny
g2IsgRWRD83F5N08szdwjN8ElV5RbDJ1ICNEBNuwsbpIWe2v1QThPbho0sDMRVwn
seTTuRXh4q/sJETVfqwIwX5lm/Kf3Fh43XzwDlwRyMTc7SdQiTa+LNbyoW++P+Uc
O2SiAYYsFMaXAMuBlQUApC5F3V1ZOw/hwPB4Akh2zDXKCIFUjAXxrqCewQP8QjYL
zjRXKt8s8rTW02NajOEe/VJUvgodUE1FF3WPBW+zpfi2LJv6tiK0Np6hdxn9cWP/
aV8Pw8FC8WccFys1CnFg3uGJgZLlce9baiaSTlYqJAscY2mDTapRNwpGGwIKll6r
Bu9v4GbKtubaTfoBFFDs+zO/Ir3qDEijbVBlScLKlFZa0jOUYQpOLyVWHkaL20zD
J/fZhM1VqhqKOTDEspV7ueUnhrcxt9kGRNDIWDjNuSloS/HHyw6dfLR7igVEaXeL
/G88MGz7QktQ6l9EvSRXYSeHU3hnsmaRjMSc81Way8zsMhKR5Arj2ZGWG+iugd59
9PCul8kJb5n3LPu64wgOntrI14YNHFXA94RzPE+jvhtARh7Kpd5WRocspY0kqWYq
LpRubUTdlbbz611/FlrsJzxx8rd6NBlKPWpfbrqiwKKKfznn1goal6xfFIHH7vFl
jc1ZWnc8Lp+riERckPjrcoL6wwKUJiX+Aavye1FL2COr3cB0o1Af4uqCXhQWne0T
QQrgIhEAZSwWjT5baNcp0fycaCbEh0AAONZgZhDR1wjDg/2MmdqPv8BbwN8XpBVZ
T0lFu2BtOZAcJ7HMJMYDi421IOKbQzR/I98Mo9LHTOUlu8x5ruSwg9BBeMYRLBGw
JU6ciN3nFUdknLAneiaF8rJ9u/NIRIIuSJ2/2TavIoA8ZJs80w7R3TbNZNUR5kZ6
oRNeFYF7xtuk3NSDM2CFMgU1/YMUqLht9J1HUxap9qkncSsrME/G/agDr9uSfb1D
Fpwy3N8QTlFJvJ36AUPuqCZt2Jp8Zm0tMAqIbHnA7BCI5MTG3Q6Kt80VuKE+GGc0
x/DM1o4Rh6+pbFZ8XG2ExxwPJxll/URsNWMRTpIOfqHKD1rbafjk4188TnOuVcgS
I/oroWSH0LTUcWVI3xtPP0HlqQmjwvBMgaT9p2IFxH8RKmLH9aw2cisnyNOKFXTd
nfBGrzSFtA/FdnL8v99F67Y7aZIfUcTwnGMsJFaU3Pz5BrBflO9CYoMCBg0N3SMS
gODjZo1PPTSu86k6S7AI7sbymTP8V/J4gBrcr7XIDGD6ZSoi/N/502CefHmu5m+N
cDXW/I+7nGETKvPOTeMEPVaimuZDTDeju0M3EgQhZEuoV4uJDCpy6jkorUAj7Ihp
0Z99p9OuRnzlSx2YWAhvB7t15srhhXTrph9KNXT+1B5FSUsi2AQ1GOaSB/L/Ftyo
14fDEh+PVG6Y9mj7kR2WsoOTc0+Tx+Wipp0zLpFJReHpTqb1t+IqDdk64hTFvEwn
xeSroGbGTctEmXkSGqnSweCOgwrenum14XsvbtLU2rKL7bT5BvwkoOK9pxELOjI9
SaHkR41D94ep9ior6fV4faS3QsQZKh0iBb4D6M2IxDCfo8OrR7sAvZ0e2+vK9YtI
/JQQhxHA/vBWJ4+6NSAglk4fY1Vo++Kh/AZvrlGpK69wzidPIh3BW1t195e76C4c
OOiS64u9VY5gtzbC/glz24/TltsbM7855sgkndtJdSmreLO3NJxnSWpCp1ILG4Ty
MaKxJsAZk6fpj5IKTxYSyMQ3/5HBSvU6ednochQSjef9KqtX4OdvSgAHC2soHT6k
ZK/ndgoMPPGJZ0Y/b1ft7iFgtSv8rTPclyndi6wIpGa3XgEo89vHbubSXYe7s0E2
ONe4wkFZy/iUcYx8gc9HN6glWTy5OGfForR286MBOZ7k8BQRZru9LaF/q2R7jx2l
2Ju5RAx7vuaXHv07ybsdMF0fW357RCuDjXh2Gzv+PUqpjVaaXF/slkjc5koBCF1L
bpD1m7DwY91woj1fUbToSG3tOkA0ivL4S2Qn9hnC8oUDYzQVtCC9cfz6exbicbmJ
QW8u2BLEP/SlCfOtu1vC5Bi8e5iEDRH8WnoF1lQUEV2eUHphMOZ35OPtayES0K1K
WB5TCaDElCe1JacCDRD/wZGcX0gKusAQjsOAm+lVtKW0jbKsCiKVUDRXJvxfufT0
UhApmRmqVhnu+K03JA7SE2AqVDYyaUC/5qJy9RYLvOuCeGCGBsoOFjarAvPJdDFg
cIu97CqejE+2ER+k8BXekhgjfuRHtK3h9m5JCLwCvFz6sDjM8nxJieiTlvZZBiY2
X8x1Elt/2zM3Az9Gix9n0sHNUbWHr55ZaR3dyv4kjfMdhZbkqAoTv0INGXAKzUP4
xU7KN/tkfuHpGCYdKMys88X6h/ZurxPKl6GiZoNgniUGxKw/68VnJZNTjU1GY4/U
AfIGH/Z7s329k0f/HCwyp6L4PboG+R1zOrzeurhX5OTMooA8JcaULTr3mt408lB0
hoL05mBr2slnlBavycppLDSSjPBRVFV/jl5ebqTq0ukeOuW/19Qi1oRrQO5Hzgnd
8npecFvItFSEXEtxndqdRKX/gvzJpc/YH3bFObuTfHjlnR+6Z+KcFEoT4EkYvViy
sZjT6nGgSJ7YPyxuntUE/112MRa4e8q5ZoTu1xaWqqFoviispU0Yzts+p9WmMqU+
bdpQnnI3iiDtrbUq1En7FJgqpQt7KDgo+2hQ3jB4OXF3RmXYETGRYhn9tDdcRTt9
PAHAqGEQOGJakSPgy+Jci8QX6/YmBqE6RWR413q/i2VDHNERDBUx3kS1GmgXircu
A1CVROGY/ltGZnieHMAhKxXVOJSw6klBNQT3oNK5ZXwBdIqTUPkZ5EJG6YgsxYEP
0/L4wsZlVYx3aHtHLphfwVJb3d5kaBjHMvge19xSJnjH28eVtiTy1JDGNhrMW0BA
2WAh1uYiTeRENY5G12UaxIWzGIIJmkVRYg5LmKsVOSj55YVlCkqnZGFpMjOGHAbF
kS7VXikdPXQZ3KMNGsmtd0LEEkKJplAPRCuDwbq8F02wjcYyxki3WUsEQv/QliJj
3gLZ/6srOUqYBrKtud6Nry/B8aHPAiEzol71o5kPEYvULDCG2huuPh7bC7ZKJkjM
tBJWKLdKk8NhBphM8UA5PEIV4oITp3i5dHt5Mtnvgo5JbNgRHN+hkbaaL2bw/4QN
dr1x370agXVWE6xar8Senx+kN8HIz8mIArU63hD6Bg8nJINfNd2eLkzp1rkxf+/q
O7PVUJ084TGz49M1pWRfKMrv6h0b9nwNodrby/TlPCMa6ESfHFkZ6EaI94NGOZ82
gKDS6+9EnKZJuncpvzF6H2q2dTjB4dkkL1aPxP+YSxRxOm7sH2HDdcmtmS8n2rz2
kWr1h0ndMKx4X6XR/mC/YQy3dvJ//MlcWOAW6wUDZaDdcjOpKS6RG+ym1/F+Y9er
sr9pG7agRa8+AcnGyl+54QibjSZlZS4A0Zucn2WAo7DSp8KxOiKZ0fR6WoYRAPbW
YIXcOFDAI4bR4fKCkx5LyU7acpwGMh9GZX0vkaz/3CmPyrviamtGXOkchZ0QhZFv
m1GNjJDCXVOF2dIPUwOhU7mr39c391RrrkSPKac5uypiqMgD9Oyaue2Fvv0VQ3pT
iBoKvXD86flnVee3VUVlEQrbGnvYm7PkUaAsTVLnZ9neqG9rLjtfi2Iz5V9rrHvR
2Wg/QlgyVk0SKKsux0bCN4MrAYa+QJd/ecCjoAaB9bReYeCSx7ZOrNSX9I1BDR2g
0HKEpCfjS5uPhivb2mWog/md8CXvTCv6FTIvp9fdYFEHpdy6Y3kPT4IGjkBI1tcK
Q29ZMndib+K9aCLmQ+4P50Q/2ndW+vQltHrP0bf54H7qZjZmnoQMrxT3xr3bBSof
Wy9D8gC7KAQjJK9xZX49Cz5Ip3D/Nr1B1uQebEnm4QsJGc7N36mqYCy8eYbsenyy
W8si3+UAdXfBog4FMnJxwf9w2oxjf5mJVfho+3HidHdSLeGIKoDHYo5I79S5nmG1
5M3qcw7LhxyF/taxkuIdsrByjPqT33EpK2BkM/2j7EMptwJmaMjcc9HrpfC2FyPj
OLEvBTJU5l1deVVhyD9xPm9vs8d3Zs7m7x2Y5CxgUOKbLdkJypbpitjHRmdiby4T
ANpWRoFxuXoCoOvIAVXBU3sqa+o97R3QY3V1BuztC6SYm3ZqGlvnpg1cGISYxsRJ
2fxmgdRYoePNFXXVR5dj7igWNvvHdhpJQoZfJo+T1TeGG435sh8fXZmEazmcFw2S
sjkq4P/ixnjUfj4jyQe02rU1i+fu8DOZUVEztPKxgnR+4BLMxoJSa0kLvUrb5Ta+
0wej5XkJQl4Wo2DqxtjRxdLUIhvGS7/2Y13yTQlspw7q2FJUPZTf7xrJHxONydxv
OpQtZq1aQyiXrfZccwSyglfomJVhhB7nzdRbJMyAbfb45qSjuyGdmj7FNBahNRJd
Ijy/gSwjx1H0oTBk1ANkMu4vi/HqNqUTqUtFGaMVgB0VVGpTcuKMdX70eK+uYEry
Qp9AOw+ES6aBtgQEdmdjWSoEzaQIHHNN2/4jXcxQbCz2TmKEfDkn0hMxrOn3e/5f
BKckPpjkDMIyQVm9n0QbTK5Uv8DsUVVBf6M6n/J9XwaZ6GlGLO3YUf9k3KQxf8Dt
AketrB9oWfl8Une1ovTmuG0oheNoTguws/p2ZryH3w7eGmkjz3NkhQb12kEZi70A
1eMuuBgHM5tM94PZVF/fSAnLfKjGVGvsT6SgfV8iiAM4VKDtJxhqs1Z+5LDW8iJO
8M2qm+Q/fsHjhFQ2x5Ij6100nNILYN7i1JGQmvvm5i/irULOrUKI3YOvyiEyZKUv
fnYwjXXbGNjNzs/J3OP2IzrgwVmbWD4eMGzc8xHDdeJEtUDHHGTZmym+ji1tfBrF
pYUQaIu1xZS9JrCzPzRMz7b0pHplJkcM0aWcsY/NnsB3WttbpQmwLx+lw62UuYm1
REz+I8rdSP3imkiShjvwKXtNvtpyV+GVqOb+ByI9cPXKY2qC4Ksm6ZKmvW+xv8Y/
x/5roXPfuHSSCJ8/M9mQ6F1tT+8dFLSTnMnjxcwTz/wjUfT9IJ0foQ42SQ2r+3zG
j65z9TP9uVxTkjn2FnWgpTQxNsKi+2Ru8yuZe2dGCzel5lyY+Et8+Ao990L/yew8
hov1qFbnFHo97/zaw4QoLtjicBdb2bizW3sHR0kT0rWK0Wv8RX+Kv1pwLG2NBMf5
RLY8QMZTZMVRH3Ad5kgixLAn16DK/IOCyK53cV94Zf7M8ADoIBsKcAXTxr95j2Ap
iQa3TM2G7614euEQm+RKeGqJfVftLLcmATqp0ppBotwDDJa81L2A4O5lR/CfRCnz
Ew/K/BlFwRWFlWwlduR6hhcZeyiLdWhB2VLu2mE28ryrCWWImqxGhbu5Jk5LRdA/
x8rexK6hCssl7PKRRjWqU6riJz4NUNAauLLrQ1W2Jn7+3OKw/Kv93ZRFhbMh0S87
OzljBIcfbex9aC92smYcr+Omgk5T2N4HTTHIoE58ECKGIEPHPQEipa+40f0WfdmH
6+8SKbezZGhQAjTJulM9ZDOzwBWFHdmY0gEEBJKtA4EFAuz3EbcjUWhx2JVS44f5
+LC5t2AKeyta2IKTsgO8aYw8+/gi3x8V+KsLDf6XfyTIOopn6xssM3SHyVXLYPSQ
5coUfIhwMUtsXN3ihkiRMVcmP0W1D4pOC+jDdXkfn8sxXSk+YrDIL450JlUY0FwY
ZZARO65C4WDhQTFIVC4ny16CUlK7NWrArms/2DgOt8lhYAK4cFJ2ppFLnjcFzd1G
Jo/8j7IdPPfcrD57pcLYWiCGZYZiqzp5U1lmbhmmM6TG/u1NWzShlPBXq+hz+W+C
RgRP/XP9JZqdQ3VWG9NJr+DxlQlMHKICUzM4rlAHdsJMwcLL/7JHeaHJl3Bn2z7r
A8dRK7TNJIxPpOBfrtLOtHzbdzMBiAR1lpXS5ot0oSDnm7oyfnwh9rLEZkXU5yfX
Gk4stY7CL0h1qyke6c+pdSgwXMxnCYcVj49K8ZzrWNIyIEKXzlMbsmx5uwKA5wNK
va/V2tg+jPaux+qAJIfGjDLVyT5Te0sx5r170D2iLxozLnkFhLXqbVbBq96kuacX
j6vGgfseFBB4otn0zkz3u3tKaBLZ4NdrPaI6oVoNusVnhkw8YXzJpM7hF4tijAOg
/VBkiZuw5O47ifIcVEkxZ0FjjYkBBeg+vZmXteicUPYDNbLPH/8RiqcyjOsReGIc
x0meXWu1NyXCq/+b7FmMUsxozVWO7vad5zjjVHN3MOitg6a6X8J4/D0nYVHHJ2nG
oNCZuE4QPPRzHw5p0OvjRwIc4n2Ioq4EeT0So4SVvm/W0OE9uNlHc6Xl72dvhQSs
Kau4fMbvunD6119uFIZQ9LLehVSNzeP5caMDdqHSP4W7wXnaYUTAmlrzTAWqOPe4
I/0riSQTWKVRLG4FEtLTIuKOnuBeR5C23O6wQpAmrEFyQO8KbHpkG/UhCZkyl2rD
+cyH84z8sTBGMvbGyjvmJl0O1zuAwmFzEThZmJREJ7icbm3DaTzV2xiwo82mzCCc
jfT03Vpw0qFEGc/tSS1GbBhb9WG/yRrsQ4tY2HAFT0a/Gkki8wh8A/5q8HKyxohw
FfhnQPR5zadJ7UIvs6NjZAJVTrj2q/tCFDHEG1TO/hDTzct2rvCmqNXMKmmUgnOX
vGCitZHjidEqGkz4KygpUaCmpX6RBWjuV9G8Un1VKIYPLuXnzcahObdlcsz87LM/
w0V181j9IOQh9BNHU6HaPrs8oR1MENu79+PSPDeIsRfIMyYVqBxZiJgv416tCcQG
x1abejRyt7M6S6hN5FRrs/aZ+RYQu/4MW3qBFOSwtwmnZqy/D+bp0fMQwmNKOl/c
iaQYGS2JYPaY7B19Jl+ZeKemlCYvdkck5IIXwT8/R4S11Qh4y4ELUz9F568D6qDW
rp+llHLWMPzlpTL+n60dMFyA8nEoLdA1Kzu0MkJkGXReNFKNN6G3A7mPUke4/+WX
hqDcLFEBGvWqwx+9pDNOl7tKVpGSZ3swhTLpddLOOFjF+Q4oguSa7xvdJCztC0TP
xpBpRGYZS2FBPNTULqt8XH36FPDnQPTm9K06IaVI0eetwEKHS5rIiNi/LnYza97Z
12yoY72DnnteiDKRml0oT84XY8TCDvs49PXPyzlnqtCSnnBJgUFXQkoRSywJeMJO
fN9mCYqc13LMzSSki3R6TtRSAJawbaGojeG+3QIFk6/0uTmJTTUVPatG+Ot36UyL
CzrEjez9rj8hArRcREA8rLCoP3VaxLab38GHf0sUpSq1FThjf+/ZOGd4hxwBAx7G
3+pEUvzQRCuzDjpv+4/45Z8sqjo/5CCgsj/8YnyLCIm3rz4lQr4YFvvUhdKt7C3F
I9w9WGlWhqZTm+dOzE9k3Is61QS7S4k47azjbc6aUmoGKrFBpjNjMvPxF0ksnDKL
TdKSgGd7ya2gs7Sg11pTy4KAoYgPWuy4BH77DQuRL9Fs4Tchfw6eAljucYdh5+z1
9GyxzVRbYOvaHbHBmrfL6EJN/vKRp1qcKKH5mCk8sFIbkyqfCOOHHQ5WB1tFlbMl
io+OIsxX2Y/YHYkDtHHSLNsE5Nio62uNW1OaghXhBZBlVhEyYNaIULvApXYoXCLV
T9aGxsMQSdoW4T/CEVNZ/BO/HcbTE9XSTYUO+c7HVzklClEbbqqVS1iEnB6Os3oo
7geR7ITgSCBiA5aclm7d7xdfIj2OHDz2/mkBJ4O7lOQai1E3E9z5lLj2xY3FABOc
4UmGRDC1qcE8D3bo7bAAoW0YSWGcB/+NA9H1dmmR96pArA1dszlS1u7wYovj4R41
+tvcD86CDyllbTPtODVtKBQ5UrCF0wzSqi6l0T8/L6eziBXu+6LBJ91LbJzS/b8t
v8wQQ5vdgsS9tJ+dTmppA4UfoSNgHo23ZhWtr3ZKrB9AR+Hn6s3mcunbYPW/8LO3
G4+L88M2RT2AsxBU19cGMXAi0d5g61M0TY6FO+t5cjYPDybgHZAUOB5YDujp4VHu
BAYn1pnl2Icm6USMM3pvoSURV0iFMzxYYw/iQj40rYn3RHwoaa1W98gcsOfQ0DuD
3CST2JvJ11csdjyBLWvSnxWPMJYOcjv/p8jXIK/uHy7XgZ6mPyNcraKEcmO8HyKJ
ZeWtASzcHHkSPoiTfyTeSpnEMt1gXG1Qc0IOp+MS38Tsoa//aOYT3UtHLAQx5w/R
DDokPNjsKDUC5bp/iNbJsS7byjEdG5SrFNvXVdwTmL8mQv26QPwABMC2jLhAHbkc
prXS3kfEZLQsjpbJgcVCigYYQqOffFob+i7m9Z4L0ZuN5yfDW3rFOrxkUdsyNza1
ykFRbPfY6zSZpWTJ/msuEWkiWPMi9WZX8RoDQfe7cRIXdwmWpnEpE5tALasGLIs3
cV7QL4jJAap+cj26HCxfRg9c+LZkYpFdy6UiZZa3hhYLv0m9iqUqKOht6G4keXG5
QQakS0sp7d6+qB7gsDbpweMxp+u1cAsUIPLqRVbGm5T4ys2t3TkSXYX5VXLVH5ek
8qDriT0agyB1nMcjyu2wGsvdj6LdyYWnL6Z5aEVbaWrMtAFb8x1thlibna63bKCM
SqZNrGlPvOTYH0VeH+kHNIMaP/icfePTbz2FK8OFk7Vv8AcizBsLLeyFKf+7Q3vP
L7vySIyd49ZXG7ZL95lFHB1PwPWNhHG3ekwb2OohgdQQdEXdj5l+9k6a2MjhRqio
jio9T/xucFnUuf52C2hYmIzWFzuTDkTgWfNyDDg1CJzfZe1ERnB6M6FmMGXPltGO
PzDucXy76UaXnLxKniyq65rKbv++mBSmyW15NVOXhGnlAGH8qHNGL+HJNm9W3Df8
10DPWPIYi1/aonXKYAPY1pzt7zR+Vtift1hXn07mLMjgGQwIn4jNnJT/UNvC5EiF
oUkMUTgCFVojjHvB8IQEpydeogl00BMvFY/ft7bDKy2DrJ38WXHbkqXpW1RvwcSC
4/zv2yhTB2e0yuVQljnJyfEFUWYpkGvA9/jJIcNpNdHWfDUSFtwg+rRBpJ9zh2WK
5eW2enX198rCpESfcNrVQkdpzqapZMnbh9/ewZup/jyEMu9Nh1jPLN3aPFZCJWe/
IHljx5Mnvc/uO3DPzcVk+ag2qoESf0Cj4fZPXToqBI4ijWioYeIpECon1djXr+p6
JFQjlKpfodWzz3q/G5bd08V+TzKbbsvexmtVq2Yz/JOslP74RS3c27kvTYcryX6q
SRRWCdKMHaqKU1GO3aZ68NYqUQvyfiUrhUYDRNXdIR2zY+LJ2n9mkyfAkCh9/ynb
e6M/j77dnuQ+3bSkiJMOHOO/hVTW1LJ8NDyKicUvhIxHiSujv0lVnbH5ZJJQE9LJ
1KLW4rmECo86eQvRAyQrfvu85ov01Po70W+t3kJw/HumpVSDPt5GD0o9K3+O4pRT
tYH79NNqVcrh2xoJaq94bWS0hbdvofJHp1UrolAC+Wfox7DBI3ptYYx4TNu9sFY6
f1AlitDPuNtxbJVcSvQ3YiVNiVb8zWxkiPz4Ui+RJTaO+1L0/4NeCdVbWY33ebrL
v94erTVR6j3RL4R7fmLFxS+jESp5SJ5UjdL8CLYx6czc8nmyjcJxnpgxmhb7H48i
KRS/Uv/deASXXbghwEnwraXyTD1nG7KZWfsUW8czD9ga5tXrPXVdc1n2pea3/qS3
B2NCfmPS8i6dqGUIji/61Up/uCkC1tpWG/nh/fx64vjSQXDHtJr4z0FRL9FxlmA5
XB4V1mFvs4QwIuSikAzbChLLo4GeGxaTlqcFs57+xFimU9NWY/CRy2MQROx0PyD6
skB1M61aAOa1EsHLXTKBQQY71QRqPiy8hCDB/USsWP1HEOwSeQxmnNZ38wtiXLJ2
PGGAL/o7xcVK+oA/lHhjW+/romVwJa8LxYhdnidnMKx30D40CBRgEYTl4ybzMe0q
uu5mU9oEO5zKIJhbARqcjIFz6WrN6cowiW6zJ4cGZIJ4+2RY6aJuRwawjYxtRqlq
6DVVUjZl4giLE5Qi5T8HfXkOqry8eihcGz/HCSnMEaL0sp4J8BffWJNZKG6FZ/JD
yCMiVMKAM0hfm79e448ivhjcetmPwog42eQv+ZW6i0wJ6xM43kNdFFu1+o3BIDHH
rQSsV8XS6lCtsZKQHAb7t3G9wfsv5Npf2cArCE7KXihC/JjB2DzXjmizjGNxUGVc
WTZRBLfKJ2X0Md7gxeM97hmdmvAU1iSHJS0FXrdS2GtnsNL2c2HtVPHz83PfR5sK
JKV+85TD/10vLpebR1ZrpZr6rydmnuxX1MDLxO5auQiUicO+n6a5VDlD5leE2DBs
NObhvLyVYbMlzgWK0tiKbxgdT2kRdaqU9gXXpUzwHU7qV/cZwvlk//TGI21wiFwt
4M2uLfJDWBhBAFGdLvLCicKSurq9R/ZF9qsM08Qt7cvm2qvmWC+oPDTqFOLssgQR
2Hk//gpAxa8IlfXXTbLHFMYL7rl841QwN6dxajzUpulmZbue1hELc+42yBjUer6Z
2hvfUaBM5+donrCT3HJ+DFrb1wBs6G8Z7IDPs/3HuwTl4fG/NwQwCKQF/ZgGpPPb
20di+sDB7Oupd+hkl8b4i4OKDBntOEQS5j4qVTAMrL1v3skzN+QGOZtiMNUcqk1X
2mm7BKVWpqgOxFy1BLqUrpAjnVdV8AvHbHBj2vEmKz5IRGoWjZs06OkJZn3Si4jm
rjGHlKuaqkZRatkuiuY8oYc9phiJRGOTHjW6GRfqpzc4RN8On8MqZK3xNIHfPQDl
S7jxeWbnpKM0caad/Vxmdl+FsGY82Q3lVOY7OOd2ZKG4K2CTqMK7yryrDsbuCsL3
9vCF0NOXFp1B+hr4oGOl1xCjb01Lo6nsVtTTlc7TNhYMaEz88d59qIbkLlAd7vCx
AfCQSZaZpUKQ2XdPvyPLen8yPVZL01jaqCeK6sm8Y+s58LDcqAGCGCE0hWpnxndj
w7HnOLgHQHtCMHDDyP7H+Y1SwpFUoHmB1YgdQ5xXTaTRLz6qHKfhHtHZfHT+3+t7
Q4CfUunmWSTL7XxRl8+yv6+BAvFaNX0JURdxcNPp34BMiAIq9HhVoQWKS0vClFiK
LFDHJfM4sJifkjtSYVcZT4Reyc5JqTi34ccIBzUKniRFxqheZ9gi/xnRB1ypt7s4
lXiB+QTw32HKa/REP7BbYleq30eSgP1F1+oFN3GSWx4W7UDFKtRqtF5KztQoksOb
ZAXMDB7a+vVpepfPz8o609/zkzV30nN6lmeoXxQwI8wNNsR1EE/u618rZm28NXCv
q+vMxbvdHNwYU5b6cycAy4Rs1shaorKTbLDW+ZS5bqFNptwUQ0rgP1OYJlAlGK/q
IaEAbwZiQNomcArmI3/hLSMF/I5FWyZWp7cHqYWT4yUbvM9L6U0I3qXiPOvqbljc
Lc0hf6g4mEMCi0+f5sBavoloI8c2d04MgxNqzH+OpXdhUHVld2zwQRqFIJkMUymA
gUF4ayulOmVKQGuFw8Wf1a24NJakeGEsRnQR0dKnwk6KPggRd/vN3Uzm4S4TPIxP
96fCTxRoKaYTlrrRihOcmc0+S2hsGo8rEU2Qloe+BEjWiTVQwVOtaVH1xd+/G0HA
vP5w9IHC6SiN6hSOUH6IX+MLOwnl+beyo0gyPjcqclkGZLHg48H1oh0FhqRfSEDv
TUQojxvcQqS4vxhreCC7VV5elHe3mOZkiM5yYxmv+xuIKSXkGuXayXlbv36G5ex3
FrPXGTe7wnQwZzg2C/vVpKShhyjOFCvp5/dTayPjcyC1IVXok2+Zq+zO0+TvqPxL
h2EzwjqX8gQbd7jAAaiyV9vFmBh8Ycgo7Cc7vVHPBzKJbB7AcIjlR3hO/w57i0Qj
hi6tHK/rhf2pw+9pvqDM4bZpf0gyen7YiNb5ZPvgCAgpmZ7KzQA6UEKlpngF1fRZ
TIHb5JOUbXVHqsJ3B3z7hhKaSJtnF12yNzSJRjWzrn/7U2eAvkoQK5Zhg/hXEdCm
md8Amrjm97T+73L7ogKv4xXiI8Md6Mbb0Xbn8oBFJ0tMo7/hsV7iCEHf8B6R3cXY
7t3FNXNnpF5k/Chxc3bLd8HGxLL73O7PdNsSRA6EAGLvah3Aekm1F3NJtaXlySd5
9txwhGKfBezZj0D1C0q7zMfMGn2k5tjO4fVeYn4G/FZ9bSw7O+R7z6IIGYLXyfle
NpXacMKF7+Hl7l8oB+zmPB5vkb4N1GKOO5bttpHsLhEF4V8Zepb2FwzS8ag1iKMF
ONBgkzlVQSjYy0wsIuxwPoh7xbvTs41IfuSDRaBrtfCBAUM427Sx6dtB0Lhnj1JZ
g9yE05VqqP4ecT7gy7Z3jmfxMPr2ZhnMSgML3AF+0ZwRWIo5kIUC336/o1c5iS3e
vKw5/IuUPqAxJxx2EwwIlxDUFfWHdcbKb5Y+e8PFo9oOKCQDtFm62Vnf0MQRmsob
uAj7f7/kklQrkSGGC3yAcdXJ6Ln2aeG9quIsWWEnru9AaqSCoYL22ie3EG3t4IDx
7KiOJyfT5FujuHWN6nXCo6MR+G5vJ+4pzxT5PNzCkGeQJF/yAfm2hRap/Trlk1Im
BXxuUJcbHnbHpJ/aDdeARY60RVvI5CRXbyGWOiPdf6igdrY7O0K82ScfrinZslVb
ydtuISQeyzj77dPP9tMdEse0VP5ntniyrqMioArMZkySUgjIRqK1p7Vwh12hlhuL
f/IbWzmh1FS1Ko8jAwC8i8wIGwMUw4B/uU6L6Ff3S8wnnHtH5b3Ok21Zu7/Vh+xj
TMDmIlJBNGzaGViX14/bzPUAeBM2S8lG9E4l4FFbx3cOHqeJa51ZPuJLzZRMWyGD
hA4pbkX5m9cDCX0Ig/twLB0Ms0hUfpAl8nfxSq93fW7SrAxZ3dWP+b0oUPthzv3j
ECRSqXgmZsyNpykAzDuC3pblzMwS6Q8sy0D7fG4VYQ80INNnVO5yH2Izjag53zem
7hxjlfbmY87K3dygvKbATdVFk7UAfiDnG2V+u3S4vAloGJnMr9veZrIxcbSTwOwk
8HrWYxX2MZZ3PFaHgSiSV5CevpEoiPSGrZkm4ZTnllGbva0Y1ohKy+LcTPpMg/RJ
rtZKWpf6x3QK0t+7/0Yc3h8VeeHcth8sNVCZye0Kqu5v1g05yb38R5uEJZQLCBlj
neBZrLOTYc8UjdFh1UunN7S0KWvB/ND5lDAoPjmzhDEImJRtFPUEO7lDbVNbE/PN
pv7dzrSGkKUs+0bqUqHpZmRhTSRkhDNVI7yc6BYNMyZnnw2ziUA/vuUR7KJQWF71
urEJfxO+A8azw8Y3coyhfa8R8Uh5B3yw84X+8aqjJI4bo+wLN+RnVZYHsruduQYv
VIz+aKjtdg4+MuAitm6qd4ParZrRLViSgqpJmVsrGPuoWMFBytami4SLvkOk9GPb
nBxT2xfW6u0AjxUHfiHW5LCbQyoAC/HgOl1cS/1kAZgRkg04/ORpOhvYdDTI9aRH
nq3dltdWXMbNB4q3GKx5OA7OkIE1rZlLdY6SdWLTa4CdlKmxy4grndOB/4SsAU94
EkrEynM3MQgk6SZbsdbaqiaq8PsE7e42+0yVx/j+d0NOHvnc8nA321POhWZ2q0A2
ze++1Vn99309fHWhyKURQbcWYRo9ernjcf9N+YpoiUsqfo2BHGGDNrNO+HC6DwiO
njDm4OEsmyBKoHAq6d5pARzMfAQmamIayhvLw3myo9NJZE1TSUDxsmYmWycKAqGh
trD5YQmxFkTz+XJZoUlirmyqvZZFevEEGIYMZCKgNC2xy9fpav88e7UiTOlYicdx
+/ukbeqBT/Ysma8wkhbOFcZT0BW+QlF+wi8RJBlj50Lb64O2jG1YadQmplPdpL5b
vBNxl6SjxehfdAxx4tOEfoA30Ok18Vh9fPGQWOyPyq8H8CPFeqRsOBdaxchgyZfl
OD9CeBt5TGVfbQDxgH/vHk6QukBNvlYlpp+ed+bFJ7g9MCmwFFliwv4aOQ4XJ125
w7hBbq1JZ53nFz1CmIMsWg5FquW8I2KisA77cgv/Mv3A4T6SkHfgF8+d2LafX7XZ
ry/sHgd9+1K3roPyPHn/ge9jgdYUReh719kINvqKMA1ncKdCE3BN7fcCdLvypjzn
Pfb0Uv+MC1JgRh/ZRwKjqaVskdnLYdIKSNgnkZwL0JHHAfLrTHed+lFhlvDV7+wD
/15a6vqhyoRtAjEzPJV8RtUsZTNsm1BQmWVdMZg0vrcGltuVM7cnvCEXUncsPw8a
sDURKrGJlb8fp6Hz2QONvzgVUKLxMrJckwdEh45fU4VxRmtnnYoh1lqE89N3I6rT
Z+jnprGbf7R51dZ4DHGDj+z6QV60wGh43PEktql/IDFN3TMsSpeXY1eeoEMA6MYj
aAz8ebLTnwXh0JcrUI/jb8vgBxAzmQmEu7vrKYQ+n6aGDin9te9Jap66gf0WPMpr
FIUvqI1p6BwWs0vkgqm5mUK6H7xVJbIgiDLtZH66QPYLVYQgIOHAdXAqGuAcm28q
IgNAhUTvJF9UcW2SWc2VZv+67S3P9kWyWpq/iuxSgcR0mRp7g538wg+8Bf0FeuOC
o6UTZAmk02ZVCGSsE0iWbCdT4kK3azGQj3Whilc0+C3RKiPy8YsRiihlF6yV6cvR
BgrvRADM3PHx18Okl3lDYIudwPJJ+nZQCogxEfyywptsttDZLTirfZEZoqFZ9uyB
bfTbxcHkO2/eQC/oY1rDDR+/1LP7I0fS+bleDYLkUgkdMQliPjbpEjamireCS8rU
5ybuAByuG7tYkvKEdEVFgDocbamsKy9/06jz8Rhg3eOsJI9pi0ZBYzGnQvrhih8E
QUtQGBTZE3nNG11bNR5MWCkwDCXiNWdh9BykCF982L8urlYKYnL8NY+8hJSv8hkr
QqfrFHwMK8rFxNfoxykjPSylpz3bqCKbIqFxc7FfMB2C0Snatpw81TpfZEZYAer8
bxf6XECAS27201AbK+g/VGDS8UhytRJbItjQp6CKbbKs1EH5hs47liLcFEHfPcSR
KLC+JxDZvDz+13RzHxq04AhjxEE9f9WcrVEV5tNS+jwJ/Kvb3Q7gLKYHErQw8/+3
HYEgI9DKGC3shVoc57adndz1+N9mhniF4PFKWongEO1+qztN/PoAIeI5hMxus+37
oM+840A45DdTXKgRsgXvtvFfvd1dOWbcat92NL9+NAbC2/0tpSCypb2WcyzOmD7d
bI6oxAdGNF5YKGkOciIL9uIlYYAXiXpaddKOOjWdv+8TjsPpwsKMIwoKWcP9FDkR
MlHeO0XJyaW8jnftFQadcvL8wSH+TYTgLkQgkKM56KT3K/xOT1fOe0LULzooeMBb
lqlLNhjQGozIWolGJ5r7lrm2abmN23QEKDJOc3geWOoqh7QjPt7GHlGUrWmwxsJg
RQcicLrd6ghLpwNqkQ9LZ4LLUOOieuW6nS7QXIbNR4uVZoen7pUqzYN374owZAjE
Z+mJ0IQ9UwzcXpKhrJq3l6UksalzhQrR0Zf9fjpMXl5I47DT2uSxels/mRPLsEqE
4CbYT93xAoBzOoXV83tejugjSFykwjksV0zJ3DCULBWxss/J7wBfd62+clVYb50H
Ej0x+LaRNt5SHyWqmc3gdxvQMo0qR3IJcSqHLMOabYo5+uapZ2qft7HACjvTLKZp
v2A51+WQdLGtUFV2F7YCNrbaJlbcqSViYhgCDHiHaUxC7ckYZQ8f4ow7B4VQsxoN
IdK7PVjMT8r92BGKw5Pc3zAXLIrDmqzb+E6NNnIcJsGANON148EhEPmXKMYCbSgw
updpTz43Bio+ngU9OxSQSnsmGGBoIZdsztkp7bJPd1uBk/1PU59uI9FT+s3SvWiF
r8mGgNU3ZJDUcvaq8zQvFlEGx8cihhJHeVbjNxmCbyVSxjD3horWxbYDjgNguTas
vlbhHXtUCzvwZ0PxGYGDiirsb2XMeCqaskBRAMIXdnJITAzZZFhMi/HAWfWTW5Qs
wsbNKG9jq+gNn36DQ/dffLlEaAYMx5GLoowy57w5ajfuibkm7NspO1+ty1LwqtGo
/sUpj1W2/D3tZ3G8A6S0FGXh0QVfVfn0YTJD2ha15UULCf3Tt5PRy3+EzdIIHXs6
UywPlg1PQShpXAbRqckeyHQsXixHzxMy72kMIyQBFH5uvDvXNnC4FLTz/2jcc5cy
80ysVjLkVOs2pw6dCNia+PPcjhztk+nrLAJmPUa4VUntZy3K1gxTtzzKs75tZeqI
VsYJJ/lzArGY9hcf+RvSvkEaTvfI3+z4q5Xoqc1s3lvQf4uRmehIj6PsisEHdJbk
H5XLOtoxTlHKNlTy7ClLknJkxrsn/YfZYmo0UgHDOj+4JxDhJS1EkWA4fP7x2NTZ
n36emyNtfX4HmrwrCJ/1I4jJaDo11kePAd7AmWhH6oATEkyrMvO3SC5672t15iJb
DRPYe8N6oH5Pv7HTLnRtyTB3GkVjWLcSGEoEaGn60D9I9J1QdGVgUnDPrnoKv9IV
E1QW0xX6fLEsGeHofvseU4y5Rftcu4E/e/+Ls2A2HfEjVVFgyakbHCl11mcbGTHP
4w1VYomGJTEe+QIEG8YFOGZs1yr8EHj50CNi4H3VPCJt7yfwkz7QIiE3r3rpI2NG
NZHgTJSekl+Uu5A2C0lNTSQdNN/g6EBNOaoGKN6lVqPsFKQfRPFoP13yFliqCzgj
DVLq68uGzWcRor+8OPnDcXUenhQCv3HUDHQ+gn45490wa1z8TKBhqsD0JP4Kt/G/
T45AIsZ0aFTi8n4SVlcrDSo/gDhkAxUq+K/n2zNr16BX1rncTWwstS1RxWqkWjPI
OKff89j9TcmQvxEQ3X4SUTJLvWSOW50sNB/4/3lA+rgJ3+cPkLVdtx0lGi8XZctR
bYZqmYVv6uAGcPd+iXVeBryJlBmDWhIkuvs5BalSjX2RekBVc6mRxLwa8bNOLQYy
8m4anrDvRkmQsgRDLSBRhhQXJKYjLr82LkL89OtA+ixKhi2vbORnvsDNMTV7jw+m
mUCzECs2iHDgzFCheSShv5XwA1MDmlcVjRLkcVQ9HZIKtlMZgO4Dpup3SBlzG/SU
Z3dip9QIJ1oor/ry4MpDiBgIGSw43elFJeQDxRmT10QgVTG+acdISdS9+y3IDq3n
Tj8covNwJn0nYtk5zYX4vMoFQsaetBBVSOKIZN+pMlWRFzvfnnVCEPJyYVY6D03J
7zHBYUKWmkKh26m8QgmVOLyQIruf/1VARNEt6txbEDAGqAsMXut1tiL+J2GhiOB1
5HjbTMDmXEa7Ld8W86CCvhBJ7UZVOF6O1+Bzu5A7ZKw4gPn05qXr3O8ZOsj+1+/2
7BTPfwit/9au3Pbfxq1i+Pf/pAgLJy2+eCy3FXgj0XAqz03uwLj380AZJNThPWbi
pNtkBfVwo3ij5DhS0ST+gpwbDHjVCGH/fh6vrcS04mlQI7EJ0HfEgDzU7JQtSk39
v8WTRQ5mAV9iE1xF2Yufs1DMCjtMWOoLh2RUMjjlsfEG0iRO2s1DXMBO1pygUglj
cPkSK5wajcJzMGSBJTgMdi0ucy+XJldHY4Nk00Z77d2MBDD6nX6iJ0jtZcnbLnMd
sGXYUhOk3UOD2BKxB2FRJLS1m0y7ZBmSRDxG9unDbFgF7iDBthqqMNhNEFIm/pUY
8WPNxfVSIksh5Y3IK53DI2IqvEbdnK31KWd4lgbiWYxWllGEZ4VHnQd06Cf3bdg7
7QVxpHZauUW69ehxvYe4t+YMIho2EcQYOUdybJO8WUxX9ebfdryUIZXvgt8HcRas
Dbk5U9duchh+e+76yvQQ6J53rnS6Oqvb93kd1YWBxfRCtxhcew2w+zzDTSDJZRvx
bvKShEuFTBIWO4gKYfUChh3hpWZYxNH7GLAkqN2U6/rE9C1Ht/l4RuHlMtLq1YsZ
NgBrTgOW+Tj5X7lxN4T4pyRiuXaKhw5Jwq9oJ+ErjamJS269cKePxAbwmPY7FSg0
IFm+fXuhuZVOHlctQczF/yG4NN9urxf2+sEIdJaK1j33UiQ8r8ivDVCHE3T5jr1a
QNhs28PHU2j7Gs0GkfuPzrmzt/uQMXOrJ8DnTGpFEAorePK3MCfQtCiA4Xl/rfFN
gVZkFvjRLs0qxIK4L0e1APpq4tUZldPEGtggfKRo+cq7Rk/nee3OOspNFikGlsTp
FipjCXU4y2HJT84UTiKMZE29ZNy1y2eH0+NMydNL1e8XNC5KbKIlil0SG8wsy6C2
S42qyar2zajdZof7SZX3IdO0kzCX8rQiD9F4rWuD/4ZYH1qvxA49KFYW8Zx/J0CG
2Gn8aN/Az/ZSsURgZuXLEzPkoE/esX0LXcV8cyZlJR5MB257bX9RWf8tNtcdSjpv
RXxA3owE+r4nQwzXqkeYjJ4agaJd7fKeO3EU3VbH3v6QmZz9nx+xofooEBm6YzGT
JF+5HYxGwPdlqLjKi2y8iDd9G/BHqTKeg0upbDjRCxfS+ADvR2JpOYdK6svfLpsT
2FNh1WrbH33SnBh2YLUJtq83DH5vLQO51zK7FFPlvH9Gwra55GjoP+l4pamVvtlM
RJIkpd8VZmYq5jcbuITexv4YNTp94HikD5lD21yUa6cVuCWhuGpwIPtq+Fv7vIRS
XaTBGfvIfQUDExR6+aN9RcsFIxZxHF/AU2kJXbQbJvG1cDVxn3Bsl8TOr/TJV3cD
hDD6iXktFXzv3z0I6ZowU63LOCPycSAH84jWl+APRt4S/p2u0OW0GVWc+tMIIhjV
jTskYRv4mB+T5Pa1cjTKNDMECiWo6zFB/am6PLvNPmPRYAqkZcbtU4qqBxNylRdv
YJgOs6j8xHcxjV3aUAjlIO6cvdjSz1UEtZtVS6K90QxxiFo93aidgspf26NhjRby
G1bXpQkt9pQXqm0W3SiB/t5Yvj4YVG5nUpw44xRxnexTScMXDFCwxb61pS8nVMzo
UIR+11/UrE0RBiV8lZBIR9AUXcvsBvmxo+tN2q2Juoh+wDoxf9S2XXDiio5HuWQA
dVRcaPs+0IIKzBDypBb0nVVv17Pf5VMJKB2owyJ9xRdbfeTJggWRUD0Xws1ArPDs
K+Lk1ZcNfZTD3yo1vP3cntxaGyyxQ3Ecd59Oz6puA4zapS+j5NAvcut0dVSBJTnr
S7q+OdeyXOCMiGQmlZjYdA9AASDmmKdo456jDKKA1ATU55/P09lwyw6QX6uTrSQw
SRlmzeZAJHHKa0UjLbX5dsRb361Rw0a7AxN83EpWToZ+q7qFYIkpkd/76iVOZNqG
xavQp4UADKe0nQ1Yqeo4O6b+YgEFMZ+BIBblN5Txz2qCrgbAo7ywIHvfRGD1qQIY
pxFUKvEUdR02Q5JWyIHYw6pyMlgH33xmvCe6dyHe3TPBlMoAdNGvGHzgL4F5WDtP
UMLlaY3A7vgCdBszrB605AAeErPv/dhoYwcXmXXJBhLfkzdcFJX1F2ZdhsT68qGt
F6eDwK1MU23J+7HJBKmEo1225ciwUqQNJTab6ZZWmZ453VzqOeVk3uUKkS3sISd3
EbXsa/p0YnVNBRnruTN+q24l2P3fCksrJQYZf3ntju/rU2mdaWqXACLSmql64v7l
alLqxy8cCbk/4FKo/TITK34MiwhJ7wV5TJoH1YgC3pZowV67MQoEYbPsRytdZeKq
xn0/CESGIF9xiy44jIimt/WfI/FXeNj/d1hQ/Gu5cvxxYllT66F+m77vdyxlYNi1
V2KjE2UlWxgHa+QzMu+LBymvfzoFnS/IS5g8DU65QLe5pKwCue171fPdXhgYGOT4
2LkbxKNl1Va6vp2gxsRan+QJU0kh6uC3JU9pyq6MaJM9xHz9r9/EJjFWwHoMixMf
nHOS60I4Qx4r2umSGQL93XKX0yDBrffIDJdVGcHEgh4hPmreySeYVNRAsDHfwe9m
NNxvUR+QI9a0G7a+JD4TX3T8HcXcHL1WxtBmOJQH49Ko6rl61vIh9Fvx1/yS4q56
m0oErjho9Rz+V7N6OHDHwWAe9ignN+JRxXxkbOFeMy+Josz/fSIQrK165vjs6Y19
6Bf5fJFvLRXx6ZZ2SOpmAlwZ1IUBstmoR8jmt8QFSSbA9ZY8fzbw1elcDoY9fUVd
KAWYMnWM3UxkiC0E0HVOMpOqAyeml7fTZrVsKUrpotdSHAStDO5nqiTW4f+c5S6z
Zejsmkfeu8WxrBvG88xWRyqi+U/nAbyQjxyreExjTuDUGxeyz23BTazBeXx5OTX/
+J2bDLstrdQusRxStJR3AjQM1QDCom2+TB1ePRhL3LoHgrxMwC2giivczG2N6VXJ
N4U8AVZC7C2Ofu/PFuBHnhu0NxWfO7mL0JWniwnekPu7tUVGotXjjswRqN1Dvyff
dP4bZchUsdGBKwb4wY4tcKn6QnHRA6V4gO/bm/TJBAISFmMz62RWCaz3CoMGBHGd
l9eaqDaRrBxtCNsjhXl0pJ0rQTYsR06vRgwfNtj0/7SqdZBpyGPFVFCZ+e+TyZoS
gU6Hsm1QJVstsl7xsXlPcwTxcHu8JHlxhJ6nXAA+azvwu102Ne8owj3m0Agx2IgL
MY+4jC2+0jj59r+HR7+ukq1DtxnbFo4z/7JT+0BKPo7k8OHn/OSn12i6xdkvDn/m
1AhHneESvE1wrCGVgx30ocuoLos7HuJkwvhGY1STQSGTOCK8AVR7HCAxmJ2e+XH0
Ges8u8nWmqGCxjeIaNnNzg6pDlO8fK49yoQr8HXORxS3dFl8ZwtM0SHSn2PbSo3n
m+uyOHdEEL/PCZDqUtC++320aUgbV/2jPdkG9EZ3kEQT5Dke+AG34Ae6zt9vis8n
A35pdHpECHoHJ0eykDz4Wt8F6nOoyu+QPlqBcRp2viXr938HWwUNMiKkIo+8miCO
brAax1XlFCFoOjVYHXpJcSbfraSCCnxwQS/zQOvy6QjBa43jmJtySMhchp6qKUN1
LwyDtC9siyBCz2FXQbcPb7aTe91/Lp91Nw3yAJsndmYr4QaO8gBq3oj9Zru8DbtL
IOOiF5e1X7bM0O+fvkzfV5p/2Tsu6+rGpECd/dO6WBSDQTwnZTthWaH8S0zri5Oe
e+kTnuvZJJ8dJOJgTQAjHO1jPWiyiIBPkmdwK/Aqy670P5wWWPSt3XURdBT2ACVX
K3cf75AWxhSxfxGGpWoHyH4w0A+PIbZE1HITDqHPSSPW2bimbWsZ1imzGSULaobR
hL22LABYlyKK050QzOo7y1bfA7p/Fs92rw18bUqjvSY+8xy6Q/zJx2f0UzS63WY7
k1sFbZ79w/hhza2/3D5SzCgU17mUEJ3HdSBX9H4/4rSGMrzscBh/+XJtsysKMrXb
fcKylpYzECrm54uz5ZHwo9Wdsgei0ja/ilYMj7mUXKZbbISQT76qd6q2MbkHK0Us
UQQYCAH6SQPc1cwkteuu2jN510O4DVyK/oduioghgZsukpC8h5qeyxyjD2VhF1Fn
+irlxtAcVkyoouEznwWts+O91nrpVu3c6mM8GXB2dxJZzustXHLcThVeivMj0AIB
TsZJ7uj2jsFHv1l14d+gPJ3pz/IhT7du7OgSBeiRzPYitWxYchwt18ZSsxa4Sefe
xgQZj/32MPKoL1SGc6Bf7P3Lc0SjRstJ90OapHTUxxTs8rNwkDbBdyd40oCPKlgT
Yoz29Ac1wtFLhYgmH4wZVj4q2d8EmMMBK/x31QGIinARzitRAm2k1vWA3NLVzjjd
eqSE+Y+jgm+dhHghEwPigvBgLBNHP5xrc6gd7huem8DCz7cZXtB2xf/R7pYqQGbV
JSr5vpcnzrhRkXPVbI+P0y/qM5xFDNDHySWZiOYy5y9LX4ie5mpNfj2J5AwuBFmO
y6FtSC2r5Id8QrZHsmR2nhX5lYprghlsZe//5DAiOYMAhLhBB+ErgtG0vKDie5W0
bYiRmUMB6dsUjSLgGXDiO+pQmCOXhFLv2848ksa5NQflakhHyGUyqMUWx4LMCSvr
jCBKY4wA6ruoVE4RCcIPo8CBGsI8qcPnaQlf4OHFUtEycZqSMl0qdO5kqyPzyTJV
L4kVLSAESO12NEKY3VbTfGibRfqRRne1ShAQMQ6UbWkHGH1+Gn75BkdPH64mfe5T
f/AzKEwEIvR7KutCqdDicvuYwljNJSZg7QIByucRk5IH9YHI6VBqWp9mVW/SXXxp
v2lAIVCOLP1whxmQjq3CmY1xBdKL6F9Prc1anS6/KlVgwVH3ezOqWYkNRyfA/c49
xYqJhjuPEvUuK1PnqcOQGh+WNyuI0jCFffzSResyRBHHtXjefW5CMYOWz48xMHJD
jenQrIxr3R3nuk2i7Eazq4vVG2V8W/IBhhjFAADyJPwF+qsW0J9JysxO8H/6LmOL
UcvBpStHj/NL1lsmuT6s+MnE3yB7yhLGpE8309kdfZwYEjR9WmVhBoyYcsiTYa5r
Xgg6PyOcMTTVg09AhmO+5eGXAh7uYeEikK+gNg+jlQVKy2xZzvQd7FdvNoXnRh15
O+gM6ZNJwihetSKNeuKukIEQi2lvv7pLCAOxyvC6yj8nRLUe0d+Rh0jvzOYLLxmt
DGsmAF49GcyrVXoLdhn+TBuziAgG+0IBzrOZmXG3daENa9SNLmt270AFUrsusYFS
Lk5/qgTua4BXlSgSn46brRdL4fYG3Tqt5Zg/PWfXgjqbnrn32IdR55GKaldY9RG8
3nsp3vuhhOxl1vZQbMtV9TMGfjwtYQ5Kuzk3oCtnNNQB2fNpWVZb5+RvuLaCOdDQ
W1DXo0m6h3e2sWGbnzMTcx+Nup3h3YmU2p2J6e4sHmz8J+VGR5DT5tHo5q2he+SF
t+OASoz1hZzH0pLlTKcslw/qLFm3te+A9O8hyTxTV85WjXKDJVDHkByLTt3vbxSc
bcwwwF5TmQe0WDSg0PX2d+GsDgq+sOe/SwGnz8b9AcWcs/Wpn7lNF194xgKUytoE
GRZebnTt+Ugu6hpotXmpAR0En14tVHRqzx17gxBBNq6XqiHqXh8yBnaWDjt8D2oU
EwVuVRo6OyZB/+DF6AyAuI6njHkHGudacdlZ+FrF1nxJIDTgTSKxMf11ZKnISdKq
h8ZKNQtZduRKuI1U5kp94Ek77rSCdfC4ClA26MccPgITPv9n3rL9ZWeDUpzgY5Qr
7j5fYtVo53jN6h8iMa1btNeYSxzS78rPHAsWn2MzQrfMO1uBCHVuci7XSdWeS7Fw
J79fybbLVtWib7RW/D39U68eIqQzw+YMvDNti1VkPRHSW8uOcEeXwAGHeze4PmLY
XXjmexXFQOubTgunliIBap7E5703BY6rnFHrgb+K6stVh57UAme8f5CEV9xSpTin
QjFi1UK+sOLC7KxSN81h5ieeW1WiszfWzuzalt+vgl2BFVeA9+eSyJsqBkfc32t3
8Rvxqirk7hNEzAQvq3uoAJMWOTirpMjXIhFs0w8yHZ9agLOObQumHWPi8yOd2j31
UNKyeGhyGzdrF4xv3s/lo+1CE9rqLkBMmOlS80biN+2C30knkFChlI0hgHYCempf
+4e5cbYZ5gZMH2XiJGzrOPx+f21UVrmbF0WICjtksYJA9WujJ/Ao45ciJYTQc46t
aMg4mQNltoyzyWl7cpWj+MNpiSK5Mj0MgTcvSPFAm4g3Pu/91JhXu684uXGfNv2j
z42qhFsoBUduwCmE/hJxikZe4D8Y0APDKXvsH1t+11dSHzySLNgtHPq3ARJhXe9i
ZOn9RAdaZFjbFoPYod5sXhcBDhl+CcO6qwOK3ttzAP++f62uUmvySTrXK/bIO1ZL
gl9qq6V5WA69pT2h66ReuxBpWvG5Upq6ytsBIjxq2JQFkznnyBtWoM2ui08PbVAT
rJPi5jhyD86RacAhqSeBtjkXgDa3UtYUoC4HlY/8tb40IxBjkz8JEgOtcskAS2DS
6Zd7dVuDhJzUgsFLCBcpqGd8CZC7CRT3lp/mnpXmD38ulfP9KdafGHIXRVk7TcqK
CvF10ycteolpbkWGcGAUe+pnD+nCZ7avUQGvsQer0OPuZf01QLzq8znVZKoIAqkX
Dh0CURmSVF2a4uAeE4XR5euB6gEyRcxOwuhARh1DHImLBV8i63aZ78pgI0wuWNbh
+sjbz3zqokfxetEDiYsXBBUBh8kKohtZwudryJfkSV93c9BJDzbfZwvJA06izmzu
L4ZcojWGzgpMPyurpuV3MJtSPdX+jSXCFoNFzL1laxuDQ63oFwfnhNfqfNglV6l+
Utj2iT5/0HSxNp5ktrVQmipcHyTSrxdHYaV+8RDlyQa9iAXcHlEFeIMoQgxfkb41
qPDYoYnUIR+Of+S6vOVtRHG26Sv3Bb56KWJby/aTeb9kbHgNkJcKtit5EaVeSxCk
KR0k7cK7o4BG/1oorff/CBJwp69PwcrIWfGzFa/Y6iPVWBE8mESkrF2/ijLtintx
VQw+/GwarsPSYMFW4jiPikj71iZnyFnMjPqVanvhubNQp0U5+TGf8oJi9z+40Uex
V05Qn9GyuZ6kX9snM2EJ38HwPdYqAVsE79ZIbKyH7td0b3mF+qPQM+NZ1Zb0+ImX
bS1vsat18YfcIrTIEb/+qLnjbK28fN4XY10f1qUdAwmNtZfBQn/QVi7qGKkU2+QX
AFaZhHdkLck21AUxT+99Wu1cLwuvi1IjakRHJS/XAr8lysSERym4VujKJUPb80bP
3nhKyOUSTAyuCpRISnk3jPGIxnWBOu2JLeFdkk5M6vQta2nR4VP+0xS9izOF3BVn
ahzHtCOGTt6mnyTw1zxSUr6V255n5G4G7RYy3NSkpsYIwiU7EJZY6Hqm9wXXmiws
MM8rcomSwWl/T7tBsaOhT4BqTegtpm4TmtP2jHST5ZJy7RMtCi/Fh2vn26gtf4Vz
znjbrXgbHdceLZ5SpGx3DCanSK8maRmMnPf9towDsyELO/lkAjhhAYj+3OgiCNUb
tFS4IY3z+V2MN+HJWe+wTD937CQgQUq/SwqSanWDXzfwwPGS/1OzNtRpD+1xtgqC
lGwIHEH+MIgNHjPoLDKSA+668wB53rOOp9j1TWjyDSfXjoj6ZbDmUHxG/79hE/wE
X8bnYK4TrUE6Ria1mj5fmtj8TuKGqrDXA68da8fsbSqS7tHW+7Za2vZbQDw5962A
eEmDwJMHFnDxT2uy/MrTEq/wxWTT+/L/p6LXHKY2x0grX4+CzNZt0/NTw/QeeR1V
MLn1Lq3nJDB3MNCK1Hc1b7xVrCmYsOcgPqnwdRkvXRpJPHT4kPw5hDCH+WL/+tAH
S9xCCBRYgetWlH9Ss/50wfUI+lGDQ0ysyLFvil2a6F97DlBL7Pci71HTnk1MKwA2
ohWbKhiZZcUtP37N0tPbqKVppw4D3uVVVVOSbaXjb8Wp57JNeSNpOlHLv2Qu3rTT
u4/7BMM6HsXOJWIlhSk4eBTrGwkaMJPfBovDrk0oIvh2pCpys5vFixHGyb1HCAI8
dtP5ahT69uU8A81NyBfse+AX+GoDo7+6An+wG6SaJtWmz08Nj/dDQrjOINLcysDl
oEpzEpS5EHDozulPRylAq/zjbF89PgfSOUM3fDKCOblcCCqWOfn8n1WatYtZxIL8
zX75DjhF5tGS3ZJ0ZbG8CPYmyEbY9TdnWC9zKglUsCaFnVbvX+9LGJWLXrLa2sy6
shLL3hImTW9Z37hLLhGDPrMkOzhSCss8jLxnI+hBwqzorlWk71yCG1hQzCKgZnSH
w/WZ7/TI6cDLZhayh2BWlajPWUlYiH41YEwRIEZSABgcUx/BmYgfRGQYF9tlj7Rw
Vo5rxYzugULJVmpwFhdx18gZla2CMDv98a6sfi6sQYSo4XwAf05Y/JFQHd+W8V+9
cyHX1Um34OYkkjTeEkGRWkQzwKzj0gDwF6BRNhNYGrJksy57igr/jN25Nqbs6Owb
Va46ZvYjeWAVEFy/+qokim8YfyBu+pGdEXBayLzu1SIN5wWI2q2EqDpx8ezxpt8C
dRXbpmSrMETFFUmnztjzHgD0yLicHIbJVK6aXC9vdy55jYArYD2s9nyKh7Ub/M4p
ITAFt8wqXyp4US1qike57soXfITs2V7S9MwPXTi+1KSnZSRJj+cvczxMqUe4cWGA
Q+dqxZ79e0gktIjG3N2EiWbb9tPKc6Lhcw2SDt33oLa84BfofQJPBCO4NddkY57M
e1oW4URMNe0ZZG7DJafdmISe6F++8KAQWqkYwaBxVEATH71wziMdEo5GWjOho/16
yz+N3j5+gOsb3hkdCjeU2IkjX0gFBqjWlpHCdI6f+0JSWuXqRUdYFmwYMkGUAq09
ldLsDm322tgF1+X2NNzTyrozg9SZzFRoLe724UJ2vMokc6NdTKoFDpgjHHjrHF5p
W0l32SJPeo0mhJK1Xles41JFUAo+4N2nNUbOqG5vNQ/5WOCe7JZ6oomyi8AxNHVZ
51xan6jbbEgSxP0cVvAAHcjEvVFHMKos3XjNfg8EJhIiibs9+U/FX+7y2PyIEE/t
oZ0tuF0rN2IqucoA7lQKmG50z37Od9mRkYZj34bURDUdNsKw0sBxIcQEN7juY5zy
KoDymTPSQqGhXt2KUhChq4Dy7un5Dn71HJRLNKBzswQJqR+NtQwfJ0Vq59klFAUs
l7r3t916hx/V57vG/oX01uJDPLx52axRzZf8ObtIosh1/2L7tPSqgZSTGDGkkCzG
tmssNvA3IF8WEuVgYaP48sntCqlUnJl/V4O7jAJpiT6gFtXZ6cKGHDoPLsK20jcG
nZAvF6H0NEY0y6GXPcMW+HSlKOUfz8xrdsbfAeur+HtxSbhIOI+LB2IVLto4qo7O
bk8vbpDddN7JJN5EPv0gbsTr++KloLIKU3AZKrSnZ6H/e7eihRoks77xPPJL7aHs
5YiVAII676W6rEj7bAFE82nWg65dbg4BzifOraurE+19IYBffWUoxY6kYZsNiES8
alzxC1gPtYUp/rCloA24YfuaJlv4/W8jwFlu5EPIy/C+lenkln1gc7g/55jpo7Go
fsoJjw/L2ZDbTXvRaAGaxyOKglsY0/gFWoRVt25yTkVXV/aF6HDVOYWPPebz7EcG
yMAxKqlcnJSB2FTSlxPrjAknofbEvCJ/xqw2u7vjx+agAFvlf2FbYSb5/c3JwBMy
emMpuhsjL2j+PQwEQ7qa52GFKeqfcz6+IL77hDyf6/q3xmYK+hdigNgrbDa2KXuJ
20F3yypa8o5MtF27kjgXYBLk/506ZzNBaOFe8qXfUlnH2UurvC5fo67X5MyDUKIA
ABQk1xFKCxPz64FQUePWAAc36/YQwO0SNhkJ8aGX1V9hfFCXZhkhADLrVfrMu/ny
RVK+wJxKoF1+Opy+sYxX8K8XqXRWCAl+q2Ae0B4n2hBfbqYO3gveC5JrvEIOTkIl
jWP8suQ9m4BBMcPJ+HsdOhdwujJiuqunbT7ERRbyp1l7kYkKTC6OrnoqF4Xr0HH6
/09WzCrz5Go/skHquPT4KaMKV8v9Nops4gzMVVx+2Se1+HDQ+QwmkNCt5XT3GdS0
zdkXGJHRT5QmZimf2MoD6EKBiUJg1UXAJqBVqV+CeLSkf8SptWz38OUTPF4wf9sD
tcRSl7CGd1TuO0jJtNQjd2hcnK+IxhLgr6m1Kt4YLSO90JBCLk3YHDz0BYYTbwCG
Z++IVqcFU8b8RylPYWVeuzUG3XjY/SGhH1fGMjumgywn3bz9OYoh/D+pe3ycZM8u
FqIDJamaZ5IMBFw4LnjeCmUX9lCJeB/ipTml1f68njPrfe7vVSDpjHc1dIVxOGlR
M72BYfZAdqmZkqPGsA6r/XoPyixIxgGsm3v2MIOjVhDGUsu+H99zHL7RipE7Cg2/
unNK5DPMbxFhSV4U4nerknTXQEQcNPIeadtCPhu7wga0Q2s2fiHSAzi40ffs3H68
y536GvljYdkZhIZEvNxQouE0YWk3lrzWOJzRHSYkSVmL6do3dcGbc/wLqdlzjtaL
LBHUiS2tW7NC0BWv8m88q0/OshAbj0Eu9M5EJTV1hOuh/yiKUqzMRJyXLRx0298P
aulzCTHRiN20CH+r43FpIXbpQ136NSOZmvkgnU58k5ZfW5tEPy9N6XmHeGPD4Oll
I4ccOpkwXWA5f20PF1rZoJnJNPisnv/6YaH5gQmUqaZq7Ik/p5XM6Lvs43D9Ga5i
Cl/Ai4vZwTX+2lSDqenY94PMGz9YmdwkQ/5gQgwWy75YkYQv5lHqndfCx/eqmpe2
S35hV5VU5tsOUYVIvQM+0E7Kggb92ElRW0iI/ZqkIyyPVn+IqL350314sOlFPvUw
A3IaTcl91+Vb8f0sTKLmGOwKJxKpEDfZzB1PhquqrJ8y4iOdMw7kJJCYSHvYoew3
qedVnOQvZO4kevYKWkAHqxB7ry/CH8SK3HJnD9zj2zrWj6YDRmg3vqMXhwcGzRGR
xzpXheBjevoesaGgzmFJ/O2LGgdi2jaRWo9Oib/oROrJHKttv0fno4u2oh8zSQlq
mVriKeX3CiDUyF3jVL3EQAqFpJDl5VIeLPu7rzJOemSBMLK+xRmkV7Ogg5cuuF5P
vFGD2WCEVv39MEIzkvygWCAPxsC5Wg87P9ihBFM0CHXc4d5EpjsAdVMr25v+liuL
gpsTlM8qm8zqCjM+McCE8t3DE4UR4caPBWhze8nPiuyE5vsKoenX48Iu+tkCRwCD
3h/hxK2PdFP/Bq4y78Cl2vVkRTDwNMuccFYk23/tcbhUuxP/o1j1A04/iBSOe+1A
RXQetjWZeGiTtqIGd780Wk8O90T5hG3mf2K/wI2AOeLm6XTJ+aFArawu4rKSdn8E
pac188EtslHsOfEuu7yE7GK0NSXoj+MmJjQZVP/SVwC7UalIE7L92wsI44cEUejG
mAhfnu66DzO7MwsKQ3uLZmM99kLuhv2HAWYZ5a3l8cvfD5+gEcr+4GTDggVZlgp1
DkcUnbVaBeRTcCdcXfNBA/iHUZwLEk120sNTp1lgkCc5R8QTdXH7axyYafmcwNzx
XLzUgx6G4DTK+nWFIPSC39nIb82mLVpvz4d8aeQqaV1iO68IYRAX00pn39Luy8t4
FjDFpdTFuwY/4O5T4IcKeoDYm560gQa52GhCQHaw8CwX/wMZlyarsV744Qfr1H5g
liUy0ApILXiE0Hi2lGZ/lXricKbyzKl57k+CclR7O4zBSFY1a7eZbbxpftgFlmo9
KTwzKdOdmcc8W29Lt2TSOoPcCBPtIFLfoz9Gt8VJDyRK+8d1twjuZmlbnuckQA7y
b9ltBzJUOqnYR7bihd6pF8QiqER/SHoG5ww2up+dA/pkIkUJEVxEMz3knokJeq7h
XmNPGNixfRuD1F2yLZNVRAnXmDFIHGwWB4Y/j7OMPLj5YQCyNb/H5IgF83HZqBJP
0LDBEBL088a2ByFpKRmCS6lRDW9awyaDmdT/K1XV/91gteyrOeSgiios5PEGVSjj
RoWxKA+ryfn7cseShtHXX0HjntxExLt1WTEz/6xL/xHpVUu5ViVOs9YJQIOBSGZz
/6eKqdVSiMFHrsCHy3d7VegUIULYMBg4W0gLQVMflhVlBXPk4biei5bUY7y4vECq
DsvaHMbH98vbnryX7+10XBIBVm5HoYaGMO6XsWf0x3YMKSywXkgL6rP6Vz3EcnyD
ZemC1fkK2774ZOAlf0MwaENl4S9DM6X+gODf06n4uQS4SHHlNrkjEyqXDTsmgAD9
z0nYZsL7bXizJnvmQqymUQnmbBppyD7MVvRI5k54gKFC9IDwfKqkcljc+PJCIFhO
FcGENksqS2GshI2pK7I04jIGytF0IjLC/Tuib5Wp5flTV9qvD0rE7R+Zb5hzlOW2
Iqdp4m+t0qJBWkXGlOL9BxjXV1CVRbAe96MeF3o961wDv4VacRUYHQcgdrDSTMIJ
d3uhcOl8gCvgcp1Vyq3hTKdQXHBdAsoYb4f0llngWOip9p99zPlYndSH8Y666hnw
Apdxl9BL6g+cj1J4izKR/dMp11AXZzA+fgZN8UTiBUzeYXcOfw96+8O8CgDspt3d
SwAq/F+LeUIyVU9XOaUgGu+uREccPb9bnUPBbTR30FcHfqiT8uxRPciOFXx6v8nf
L9FVq7JvczjIfFG0vX+NZ5w2Ofk2aABbsR14ZTHIi6H1VhKArb2rMeABsK94QmCg
dW8i9AdBl2SPe2tj3Pfd9ov6kfNtV3V9xH8iEQ0qUWYnBRTGf+pjGIwfqUVTRpUZ
flhuv915ug0yQvF2v92QEQkBIBPHcLtUnVRyAexEcDCLw+HdQcejN0X8alxk0gxl
NfWLTzDYMQL/nrZsis5+qL1YzaH/O+/LPtpEJRclc6EgwjevpiOHbwcYb+bpEGuW
ejTwRM4QMUKhdnsw0ozhSl264537KRK0NyVphPl35g0NGhAn+AjGE6WjsPYM5HeF
rdeRHR9rMdy+urkcYdd3otj9yr5KSHOyOb02CPLn80M3gB+qxrLHhlKTiDVhDdyx
bUIr7aMVrXed84jR3Kh2Ia4CmVssqWVVmJtk2uUhyOT17EE/Xd8DLThTZKerIOFC
2GF9mA/kvzcnXoJ+jg0M4keAYYCZm1oHj9QhqeDGKVj9d7hEOutwN6ivKMkeMdPc
PJsOqzVUSY7ST/ZOdTHmDrAwNCtl/Nhiq6ni6hdjDJA2jUT4lLpivfL/Qhb1T1Bd
+XtbPZpB00ilOuf7Xgw19E53IriJtUcFQAIxP7t25hk5jS+Q6KQmSZk3zTZFKxws
GevtjnoYqBuPO0kVlBGxiFNWBo3l9//4dBr1/YPoWClmPEsjqwY+V5sHGsciMmPm
LxG6KBxVdfoyIsy6YMHIJzd0RDCk+16nXZ1V+Pz2DufYjHn461dprTmrYJkdMS1c
t9Xbk+KpaabhQTla+CrQliLUBpfjsluOiRBrv5WHtIcZufLwbJcMmDwIxJLsaAr+
ExnqM4GnNWAsT59IEbLCIBzSpF8sMmx2iNVu1FrxoO/OKzmyRWD3D1jSpYAOhOA2
jyqj2a2LNNr/ZQpELwZfU/I6ndMu8Pt0BiERxMcX3U76pX0elxzWgwjQLDxE3mW3
ZWG9AlgHs+o4y/Dp8lSldcZ3LQbGLyFple3s/zO3GUSohFoWPpvqUR87D9z3FevF
2ShQjBmEotmEtSToSLLn+nbB2iB9wRz36FY49a9ER5iRInhwTNWdJiMU3IdhB/uU
G+9LSb7go2OyXzSgFsNB1EGLrxaEP140UEx05wihTWwXDTK25JzmxL8UzfNCtIEZ
6r+NCTDNcq6TQBCpX5cbPywt4kMUDCl+WZtmA+q+v48Nrk0VrxToPRp5syIzxoLU
Iz5K7dk6m6I0W4dl+qpscdE4d5/c9vk1DQV9JXPfLWEAc0gj2EmnCZSKCD03HPyN
DAQ3bCLXcn2HBqsiYtOrPT20U6tdsZrWmpFZvZozPsJHH/lk9Lg2PfFzLLOAE2W/
oShmeVnQALUZCO/zfUDLzz/DK9VK6ZnpPQj5xRuKJRpJ9CYf/SXbYafbJo08p3Me
ys6KvtK6We22dqMxa60dG84Kicswr1x47xyFfh7fyk3oBhIYpiUkqIfUGrB4o6da
gHRNlVgjlZpkOA9m+5Sam6YFSWK6DYI72a/ilNWogFg3Fi1gW+odhThuIOiG1aYO
sOYGNA13dIwd0iaIpnf8xzc8TLNQiRteZw72w+cy+QJ9T4budXX1ZvUfQnfW8+Ac
LR5rKEMpT+f6x3UeMaLJVISYJLmWCXi2mc6QDpfsBB0yVqbioUMbQr1FZDSl/Vsc
81ixvPq2j8yFLBhNoXPtNbrEClGdeUYFsSvu154kWMD5hBevG7Q9TK0jZTh2MfEi
zcabNx47UnPiW5GGHz9bjpGolwrw2YQxpEaIZjTfcivU/rqcZRqjwnWCfT/ZdVz/
qxZlnbQT0LdkTJi6sYiiJYNZxaHaCyRkZc+PxOULopr4Oq1Rsg6e2KMrjU883u+6
9U4WZEO1Uw0Vz6DfAczg3S6kXgoE7nAirWggv0/SaE7/kFPmIVqSq3WwF1fCIJfM
FUHjPYWdi0xByg0ElO3wrBmJILeROznBjVoliNoQ0df1VIZXKf3JQMOD/Mb2Lo0X
h/KR6kWXCb8tL6cgTCiBPC6JRbjZpc6ZIDo10Fj/sJEl11n4dR/8jCASGarpWnKk
rStuxNAaT5tDH5x4cLR4dsTVsJ4h9KKgsXy9CDbDonZZqM3iMjAEZMItgGN9CJ1L
6iS3jmd+ygmNJ/dBSvuUdNwQI/MGCS89rIm77bSUr3u+qHTaYvM2zgSdBoUNuZAn
+NRBn2ED49/YRWbbWmZOIybFhuGBRypXAxr6N81X/rAFR/UVBmywBYGFbX884LP6
sKyuD2sXQqPOYoNHylmixa1SyoFJ9DVcvWsbXK4pbFrWU2GYqVHSn8XGLXY26cJ+
jIHI2P0l8vwPSI0IajnTyHSQlMeI3RSNvNIrepDEsEyc/30bGMrVIEgyamfeLmKL
G+J9mj7GTfqffaldlQnjVQbBwkQ0HKKSZGsavuJX/tot+5x5ayTO8dYZvsASptF1
jf0Zo8PW62KuGhklVcECmqd6lALnTpcBWHFc/fF6GxqUAcqtYCRkhKfBw7gmY5TQ
zR8mECECBL3EO/QMrmZd65AIHM1iaEihfhi/BF52gmeaRQ8N5I0zrPh0Ha6s48NV
pwsVH3uPDEa0bcYhfiJCZJnfmrZs02oJAHIeKBqZRXk6of5eh3FJ3Zz12axdVJ+a
k+6Jo5a/SXTpBPe1/BEtaV+tYMPJLt6s+6F4xWb/8X++4/GFjUJ1dh7tLrsUyhiZ
z9OfsDuLS5VveZHSgjlMF9QRJArl5xtYT3laOh8H4U3pEI/FBD7RncRbaRKjXgJE
WFOZJq6+UbWX4G04S+/Fyf7UWOVHzhFzwNAAWi3cNk62fppplu1lq4Q+VLjUjTMn
SmYG+zcPdbDZd7IUIQkUg3bEZ1oFt+HaluujYFnjF7b44wa1dY/2dBJnHTk4g4zv
ojySZfzfLuugoTiqt9YJvpjiuq6/JNVFDufTn/pNyI6XL3unUmX0bSHEyj0e/m+6
Toj75OYzFIvGsVdjW9wKyJYIRlHaaXmAhAdrZ/gkeQXCnbgwRpoVqyIvwRHA5FNE
Sel7usMw0h0qS0ZQ1ggSeAMBNLFEi7061u4qE9cy3/T4CBSpBsX+YVw+fTcBKcci
e6QXJbC5CjmkbY1L7M0/7u1vkoBrZ51LOhS8iik2jV1Djksi4yUk0aWjrx7CgMX3
1hueGiV/in440RjNT8KCrR6MUxEs4XQVaWBEBV6cm6t03Kb7/d2k/AYCJmsuAm5z
ey2A2ra+VmqDFawuCfwCS8iDI2RAWviiOT3pz0G1ubVH8fQPjJ3maoFXZiLeA7lx
zJWBmI5T0AkhldoIp+n1Ost329pmWvgOpswGJaVaYw3r7S03joJzqp4klmQALusW
azVWpPiubFH5bzCFBevscRAxyRH/yAo0YZKyep+qeTCEW0IqNbK2msS7+PtDCOlf
nznO31VeoCrudu5HTUvR98DEwBr2gRGl68+Du1XQUHk2r/I4gCpHt3y2XkV98PHq
fB0C8uWfvaZEm50zlEATsYi6PeJDqZCkEFz4dutPXCb6t5l4v3cvJU3/uguRMl/i
6TeZpKAYn5XlPIcZjg3B2JjpZfwPC7nAGSOuidncHFKN9ZE3PQ+/CYceLFWFB3Q8
mxGXA8r6plGQeu3Qm37TdfhU1ZnGAJuN0DQRByPr3Lyom2ux2WgKyg5mk485bHnP
CAh1phh/A7S7xYQcqlWiofvl9I7iCxcsoM2qdTa5UIDDNObdkz1sQTqGsRuIpD4u
FT1ahAwyDDnF1Tuh2ldZWOJ8JC7fV4gYA0rbj4x0bRkoM5Vm+SbzEwwgFF6qfaL5
ajeXWoqYAKG6m0TvGYMJY3GKUwkIau2oJ6lT39p+Ux+zU6pWXhRc9/78mbNe6K06
Bs+OEBkE7iHPWhENoD6KBVJCjDpYIGBb11PL/qvs+lH2Yfi/5xPmJR/JbAURAs99
42EoIUH6Ebu0pLNJ0piJY1R3DGkeMS/Z/W5kDo2n0P4F4fSn9kS+H3aY3FLKdF3r
3V51PNE0tA7T9DURCfSUY5UZJAjPIvsjBELaFu4Z0HPYOR9ykWFoEYPMkmJeILg7
QF2AoYtqDFOjC0OHcCVv8wD4CXQgPBdgsnKwblBU6P9Ro7C4ypOoqXaS8EnmBkg4
38RL5RSm8BqGYPUALGwh2dfPMQTGRXTxB5DZNk6U3imd9d8Ry1CxjuIleseJMNMV
PBTkkSIpKi+owGzBWgX7ifCmsXjGM2hC1Ga09ZvD5VyIJpHMb4t4QFZisB4xB4rK
VwR30B9hFnPEt1SssGjayQZHaSf0HpQw7SgYWkeylr8P4Vy2oNOKESgfMpHmgCiL
2px0rQKarB2hZ3AZ/4zAp+sBON5QtfTMjztr4dhBQXb95O/Mx0Cv5BOB2TIvyRYS
qWcoAo4iySYzvsfNvGn4g97v/UV2SHkuU1l/ocBfqbuI3X3eUGB7DiXQLvYKZTbM
5edaQKxchF41SGguhXuTQHL7rPzQ2LcJdvnOKqJ/8gBlcPvw5leiBMZG3o5QqBWq
JEO8XHweyM3rTkTGPcEkpDiyyve0S09jKr3US1ecHj/D164IvRNr6iv0b5reejYr
SUzz104uGL2OMK+3gunKwatVvovVZ6QVlpacdaXcn82i60F5hFqV5KDxcXt9eDDb
+IGGILcy08k4lXkmwPpIKjHuD2Tj6UNXIMwqN3AZ/29C9IuD2NheBsicOYlnONyK
q168ovlzf4abCVbF4CS3TeMtKks+WDNRjafymIaavxM5cCXERslvO8Yo8zvLwFi7
XIJwVbfxbEACy8SpptgYTykh+iDhi+ytpX6OADLq+MDD33BK4pX3eoBoBs0ESUqf
6CZbcIduUIALM8OmrfCx/tEEAU+KKwAFvv0+zSnq0KjeMmzz1Jd03TgKbwIF6ers
o8SKFAX7Np8SY51T28HjNG16QVxmh4gAR7ZZfAHkN9VyFzrQcLMRSv0ySawrm6rA
NHNcRFdLnunQ6iNU3muAHCYdYzcWnPZG6d0lNy9n0vqcHWzPVZrtI/fmymP9z55K
7BV/gQWBDbsFOD5S9/4LJeWXiD1Q/rVUZPGTRyql8zCsTx1gcybcMKTjoNbr6HQl
SkkBnMHeS5PNdsq+BBHg2C01CJA1tmpw6o6bjkeyCwnvVzJbQLlm8qtvRd6XPfuW
feRyiyOCfkdmV2m9R6DSq6p25KZo5jELNmhJDfMl0PlfbaFg3w/dBGNON1E893Nt
JHwIhy2QOemm0C6LT6y1kKZEgcGldbZTtabvP4y7TdJq8ivTv7hzp1TLMXEqXI79
Z8e2i9XE6a1mFy7WEVtkgl0SAwA9CQqAHDtjEqm8MmajS8tFNPmhY2AEW20Y6L68
yahOujbwruZJ+RZwF6+eDB04ALhYXLu3nDFcRwk/kA2OlcCij6rdODEzVcu8ADsy
6ByXaokUhBC2gTxLO2hq8gkqmi8S/4GYFIUgRxgEK/txUnqhoBBvJc89xYtH2cOj
GCk2QmT7rHDkNDq/hmoXKjhejSTteWHVO4tHKmKxaCKy4Z5LV/Z3UHRLj4oP2ePo
oaXk05hzsfxPEqZsrEzIXsAuklJWUBoxz+OB7Sc3+3KGRhbhDXWjydF8+D00F68X
KQk2APvWVqXkPAlQmkh4OfIrsxt4b7jUWM6fxTJaPSsh9P8qmBTYkCpnX+i/m72H
HL5c2heryihBIXUn0Vytwac3RxI6YY917nav+ok1kDms0MVzrUqZDcMyxZcRtW3o
0Wi6NUVQT958OW+1u33ZW2wv/WTgIpqYrnweMGafeljXZruy4y17SLgNFJP2XUyT
gGwrLH4ZBPsSxJeD+CvjIyVK3XiZGwhbaHLbDxdrSvkCKTjWYnypkS+kh41NOM9i
xW8DwO355fWTpjBROM6LRUCZP+rIbGKAmQdeRkMcJC5Vst6/LD5TopmBqgWUmcee
gDQErAuEi+/ga65885oMenV5oqVaVoRzyFc2jB1vAc7diYqikBra3bqv3jzO1tAW
AHOruYp656547PP02KMJORLXhFmhpFiDkS0v60RkPKgjNURYII/bVz9+oMbseAln
C8C6XWeucF8/eVs2CsbI0sSL07oFoq4206AOiQaOnDLNAKXrvpx99gFfLrbHip/A
l0vsyhAIdzVVlODqd51VIkjAiGL1DL7CPzT5n1m/aQeLZ7lxOaL+NnKm9mCUvvbC
2v8ioGuLFD/4gIPCxx1NWT7tzabr1uMVW417Bj6J36lm6R2PAhGAgxPhSffluKIa
+Zre+lt6ZnUxrzHJEZP7Zzx6FPN3eVSx+o/Pon1dceN1rn9IEeFhyZCZDpaZN85T
qqKbQT+hj4qoijacynM6NRBiNs08p2ujiRAJTRYBbv4duob/De/aSzcUaP2yQ8NN
4MmrIRXSDxTDQc9vwAtyFJXM9yddTdWHPJ6KueJCYItj5qHhz73tXQZ4rDkdoeDm
ooyGnExjKW8ctSQ40DgkdII9v3fLyadmtkGeR0NIxf1UJoTHxQitaluQMbutNutL
T02mQqsCeJoybby8t1V/K80apc8uBqZL/knoCipu+VaNl96OLYU/hizCodcROVSy
t9FSiUB9V8qM34D32b1BJkiax/Ti8QNI30zZ/DlJGc/zRhJwCdBcrR0Bx+7QIgxR
Srd7LOwtKmGIjtnUK0aEzxjeODCupyr962smxLPj9z1VHI+ppoeDNAGQTxung52j
yOETbwnBecws8YNH2AFlUJwiSMXMz8Ku5MMaJfr5pWtJ7gG6Rj2BykznJPCyqXZ5
VWsxOzJZcb4I5icZyT3Mu+rVgmrIQ8/jK+aThqfCjw78qgrRUCq8ujhDuaAt9MAz
z7MywNI+gS8w+xqbfNkhRoOGjy5fMs1eVqYM2HQ+QhGURqRuVERo1Je82LlHdZ4h
RdDqOpSC//udEnWbyKoOngr6pbYwcU7hkS9iDNAO+KeOdR1H5nvOXi1vfa9ZqzOB
xZVyfv2mm8O3Ftqwaaqyv0mUAXxGISK92dY4X4yHJOuc4Syi64vDFEtbkzM/KTu9
X/iiHJvXGiybQIkougQ/BUhDob1gs6wHgme3fCSesBuAtRKOQZsnqxwN0v+f1QT7
FYna+6KZBfmf67Qds3rX6elPsOqgpNn+zjyHY8TrSoeZCsZLm2J7FY487dRS2tCD
tFv1ORq9j/CmQH0osMfLn3s7Xkjhe6klfzFqip9ifa/7idbGsMQ05tHVDEN+48K4
4u6iFm+x5To/3QZ/WreO9Cw4paBjSwsl3//5+tnwu4HC06XuQnZKGaFf9AsphcsS
QEH6AraQWqys8RYopEivP67G0EHNDmpbZQBc/Kf58o/lUW6+ijIT4ZNfFltIoeML
KHuZQ56GZraht9kfYq5CHrr/thg8VM/vbNuECYtXTn6dEzYjR7y5flvVl0+RDnNW
0jJMzbUbAad5KzhMjiJBNPYxQ+pM+qdEqiG1oFMm+fUlfYyKzzZIZVVHZxhMbHD4
p4E7o+OgnAXZwWMObi6mciaBm8S4TQoNaR9ipNwD2EPVLyJmHMLiNi9ZfrSAGhA6
nJoUcR5+rYc7BjVCDcQM2UQt7sI62dbRw2zErg0lIxjqBW1C6wAzu09ngoVwWLN7
Lf8XCrNLCxBBiPw6vN7BFjCLkX1jRRX8MzcJjSTFtts+3j6Q6YSH2ReoeJ5a55jA
z7x7IrG0XKd9QGlDR9VTjBxO0nf2nakXgA+f8d1Z5C9+qAC0leolhkiKkNQorl/3
iV6tSwKtUiMejDhB9MdchyYfw7/5K8uY0Pj8HF+hm/oPlAAveHXFOvpcQXN/e/cx
QTAaoKoD2w4TW9IqYKLUOlpzf134B5S3CKN+Wpw3FXBRgNTvuHRbTEMYrYb0yftS
HN+5CsFW+IZ3Yxa9gZgBydQblQ4pgEQxFeBvFDBc97CJlMVqBBdlK2R6TsHq1Aah
OyjRAO3EQcVi4pTEFDziFDkd39rIj4MJF0Q6JZI0jofKVTYWECB3DgjieeLI1jEZ
pHS4qgDy+/6Hlnzyan02FdJKjyghltwCxTXCXC0w4S24ZuHWLjrX4txJsdNTSE2z
rkYz5iikHMHPECwg89lwRmXQ2ZFGCuMIF/IYL2Pu9SUb3LcvUuT+qyUh2aba4V8P
8c15PpUO/ROY3mW+m7Rn2KnKZbVIHX55Bfv0dx26/hAmEyt4kaQtdBXhwS1jHtNs
D8tpt1H2GGtD+3AJ0oFxwkxiUEYefwl7wYAL+0cWsBVm51Deu7THvQlC0Z9aOWFy
kV/yhAEwamyw1M5AseXFLHBYjEjLrXZq6i49iUF6HtOkTeQtPo5UAJ0fywzcwsPW
rukPcNTASaG0LbdiUMhuisiHfZ8S3pSYfNlTSlK4tyMyB05IVsTOnltkpbx5Z0ms
a59sH7yp/oly8GIOktcJMBDO97u+m6yxN72dOuC8U0Sm5FOG/uEPI3/2yguUUZ8c
5241v9V61fLvIbiptr3XqDjjtSU8c9sdXaXJ+U5a1ZZ+Ct1XyX0YEtkvUh1XLkFK
PenBocSNi2fFluxaeWBrf2E5RiJpiwDhXV0bjIRxC/CAR7KM1nGlOUfh09F0wHuk
4tmwgU1NMHqmZweydj/hD/81aXk3WXv5oxTj1eQFb0NjpGJfzfk7Z5Wa+MBfWdbB
nb0U56DRK/ZsMPoHmriHuIewNonxAdUXfC1v/SiYplDVY0gyv7Qc5mayB/V7/sq7
XB2EwexnLqJmwvrTePGCjrBImrdNcM+sSToIL5mwN9QCucYLle+pAgW0q/hUSA86
9/zhsYjAvcLU/Ny2eg+YpjDh6dXK8+H6D9roYYnsLbIoiKeswOA+N0ARSN2TxQzS
8/tOdxdAFqpYj2foV1upim7XUXOZIktSlRyktPw7uzM863a5CuNRF+6C0rsr/Zcy
CmBNULEdJzdbB1prukpfNjZCZpbvir4DA9j1SYKUKlBXP9uHSCp0+lOI9UncPzFi
JUkABR04zquEp86JYIEN9yTqdpkF3xHF+ySUoqGzJq/JXLjrMqHN3XkPEbC0Yl+c
3Dgbegy7oQoyP5Okqd9imKuOkNKWMfoo9wqMwtIf9g3tdznE1JHHallbzDikLARQ
VzRVMnSOZfdzvMdwc2Gmao7sPB2fCfeAQBNtJlkKcc3DNv8HSy1hVexroSxIn8Ow
TFfk868f4L6KOxT+2KsH9P2XNZceObYw3EQ0yWvV8FebAUVkx8oQ/xqQJ7Mz0+TW
o/RLaiSY4Z6yyPTqsCil+QD5lL5T41aBs9/AFQOiecdhkp7SU/3sVIU/SPY7SLZC
/WPY7ugT1xx0O2VdNEQ5ZzWkEV13B+N0UlYx/wwa+vhiiTBE5gGL6PfTiRCoRFP/
8DvmUDvf0c8GVbb+/xcedJa3bkMd1N5RGcxJtduZaV6wZ5EgaMhdWMTPb5Xcp0/T
5grD0M3pAm8Z5W8CvGCzrO6BmLyfzxb7wjqYXL+XOBY5wDImTGO6G8rgmF/xcRrk
wgRSRxfnw2PV+BYIIW9CIJgPwDerIrcxd3Wrg6kF+DGcBxHFdS3TykAOlqXvxYpT
sJQnRUeBbW4UPFa8dC9Z21m388SgdzaEE47BGoOZ+kWXWYodg0zeEWMGMcfv2Rvd
qk8gGDzJ3mJpjuZUTlff36kPKrj/uwQh8Gm6vhfo0ALhnVPKI/VysZuGk67u1mm3
TurVvQFBeln93EFsfasLZIV8v6/3RTu7zfGidTmmOQlemITTw7gS3wKUM+WdU9eC
oHYoFnFYJm2ltm8L+0NLuG3b6anLyhKO8LJTBt5c1df8CYQMjXLWXMQSJsPJ5DW+
ZDiYOXJdx4kSRV8ejGEPBidv2CcG/AHHTQPggcvd40lY1RutfJAO+kWBhF3nS3Ax
14ZFnpbtvgrlrPWotxplODhCHim/sJ56c+sQj5/OfDmJ3iVnwsv6gj4745aPXtop
IZilvy5zgqmoNiW3S4DHDJcZHttCtGs9LGIAGOvFfoo5TMiIFdf5aKSKw0TQxQX+
LpxfixF70dN/eTkCYE9XbEWWt82cFeQi2RNvmDHdMINsuNM0ZnJ1yVIHQkvonDTj
02Fl4TY5omAtTH9lFdisU+3BIVCcY9/98Ijj8d0Ol2bdYgsGPV7b8MzFCTSBCJn1
f5c9F9H56Byguc1JYcaCgeNglzzyODNXkZaqExVwJHn+MIk890wVMZr1CMJzuqIJ
q73+mR+Ei4Y9Q8Cm65oXXXdP4HdD4e8k4I+POeo/ZzD0DryHL1IiDx9TKUjT54Mv
CAOIXYdj2P9F9+P5ZiynpvDmp10wktgjQzGLhlTbApHlEFlKIx+7PMQHXmyzJVuz
54Cnjv+EUWTL18wfifcesNw8aNyBynrUhGNA3UhFgMCsUgzFsbBeKriVDZ2qzESV
Y9NLwnn29VwUBGYuMkF29s2HnCSfmb54jDZH8/oYiDT1yVZ62BuGyu0vPZl/YM2C
Z1Z9WeAofXc51TGDJvToiX0TOqxKzUDpBoTANEXvZXs77eu3r1HtHERmFj47yrtc
taHeLDinEA7uZ+Jd6Ut4MCiak/Ick4mpSrPsyPCDwLWWHRVU6GRKzgjbeo38OxGr
dD55Z6mkczRUruytiagwEz8AyMbuuv1f4AQNb6h6oZmTrUdCG2SP7XJIZEmpygKT
PkwEf1kQGh2os/p5FzneWS3w2IiNHYEm6I7qdIV2RH2YXgm93kCKNutSRBo5xf7W
mE0ihbA8u5QBaG+dtQjnpZLKjbFtsl7ln3RAwFRzizD068ilnmJc6OXr4puWQRR5
CcvUuXYZC6KVzPs8kv3099HM15Jm/afuyl6sx2Bo8fkZykSLfysP4CzuVWbGOrzh
jW6M8XnjuAqj9cmO2EfVvMql3oCh/6urBklxsJi2lYvYZAJDM+KMOm9SAue9s3gn
mCi4csAAdI0po+W4l2gpP54j+XZpKGg7uw4Z+OWDXnrYMaozcOGE1X3Y2GjwRh3m
tfdgD8oOBUDmO51xIxB3UVQKRGkEp9oYK9PUcJCXnplIKLZPBFVRbCxnQd53HF9+
pRgpXrwm38PWaUrT8QQcdzTA7kEQfeF8nyQt7/rwtr8G4T+/CeKnU037h+xKtD3D
FswFHue7vMyrdaAaqWn9PzbGQVikeWrpZaNbkMaxr1ee3XgEN7UkWJp65uXljhOg
aKo5rw3jhNSqBfKDWtSF5diM5Fs1QQb9enQ/bAF+qmk0VOd/Lg7TCfOT/wmUtFyl
qmrOzy3/4K7Fxe6MiyRuNdqXTrFR1FPLOzcTx88HOejyceWUOyNMKOnT4rWPtO7d
UeCWx64ju1W0EoVNqm+m53ira9naHGQwmO5Ejv9wUqSPi0IpJTfmpdUuQijp6b4H
o7RCn2iW1IDGy7K9R13UdqusUw5KpiW2x7w88f+jn/VA0STsZl23XR9gAr8qnnii
eLJtGnCAdunAUfGkK/Dc68Um6rUbOpjOLHK5046Q6x5GyhQ9ipJw39QJKEL3fX7R
+Y4Iz/V+wpCtppCX3BGQiS9YiYd4aEYoxa1tA2IcNsIu5J99VH2QJxcGOvy3gmtW
oQIS5g51kDDQupgBjLYO2EdOnq65i2NGuNmjrean0rBNjPgMYuV0UY+hLUYNUGy9
Xeg6165ej1svZvMiPETAb0+VFfBZY0hPzp4wsBuoKTXlV4QTcbCZEHxrxzE8JD9m
Ll9DHQ7VUyQJySmpH5IgAiKh2PfW5OXL17Tqz9AgNMowmBmZXK2ilHDH6IzXXvWr
uE30PTr3kGtU2kuBNZyqQeeZE86vF4s2qX5xUXmMegxaO36KtAnGxXqzhXWi7X0m
NI1eIPVHXinFwQnyZkJpTjG95NkIUeI0d/FsMLC/JdDS12WuQcOflWGPc0RVMJ6F
FmU8O4xVAmMVaQGpJzDsc/j0IoU+5ErNc9pja/QEH1mYHXkmZx3fP8oWMo5JSZL0
k+tr6bRuclA0q/cmR8oGQJBJ5vvaEJJZsB72xue8OT18YkI4YE2uCrOKZ5Rb3uCV
+gA37EzFJzBLf5iqaNhZF37+suPMZRW59YZJ6KGngSNMu5HoPqWWC255IhKOlFvL
kOXwNoJLvIFMgmfA2Flv5g8PBV16o5jbXUuSzvJM3cTlev5yzUbuxydY36613ZyY
bv0PXODk623q+nAJdnMCTUTk4GtxnHzIX76X6UFEgMmuGnVZYX69MN17oeb+oX00
jqFlaXYZVe4EmqAeYUoM8r0RjtMFOU00mgolGMXrgQs3QURgjRYBgBbuqSVjfBsQ
2m5jcySc7b8JBN+mC2Aj1t0UQTX7upro8dwmuHqgQGa5zrZytfxErQb3co9ll2va
3z7tTRJuRzTIp7/LUCfBDFHrsOT1f5lzpMjWTmisChkwhHhWQLOAPI+0ueQUwzPm
byvER9Ql/K1pVn5TVpWo7/X1J4CL90pG3BT+X0vFd17svOeCCphmTagEd272F8Ou
rNIgIKaS83TPxtP5LylQ+xntiPuKy1BxEDyLUdku/pzuyYTNL1tV3mJUE0VlTz2s
UztTrh1rebVUMosOBeJyjLkfUmcgg28C87h8wxAztZX/HWW6kkWojjQnpxbJLLYn
KYkNgL2ZdbeujODGX2tclgZBxOTxXi9n95qt+i+KdJAqANMDI42KaMB5Pz13altB
XT7TH4cZPrs3R2Rr51Z0ZJao+Wca7BzoM8vXdXRKZ7Wf9HBo7J+zYt6mofUYey4c
5cI7q22OtHM2ajozwLH7LYLnKjPYavk7KpTXj7V1zrj211rQsJOW5L863yv+Evu3
HYM/slW9egPDxi4R35vRqvg2Ik/mqp8+tqAYFjz9DtMHVMLyuCI59VIlX4Izx1SQ
we/1AKuu4SLPBpIbXSYjIECHrhLOhBx7WvqXU7tpWkhK3mq9uWaEX+BAISv0iOCn
uMbdGOFzYBwdI3+wUDUHeFq9yVG6163RAmNTzhSWZjIeqsfNshfrWokd5ODBF7ZU
TMCJ9o7TUjwEWX+Har8vqZQzHzgiimVNXvYD/kHSBPj/USk2CmVoH7EjNhnUddDd
S2aSBIlwuoQ6KN6I31tIToRPcC+aHQyPPWXkUV01/YzOeDIsIQTJIJOHcv7TPkUq
2O8feMdopWjtny5+iIEZOz/5pgePX3g7gTt6/9RiBVW4dzLf5sVaxlYJgSoyif+d
2p0ULKz0fzvhvSLfhnwtBVzDLvm9sHT1LTGLxaTz/46tqgdD4SHHXlFk40Nm4uhw
OjFZE0Ro/iM1Qs7GXLI2yUguYxpdve8dtyCN6x50VWP7jKyt1HWzIftoRb+/Fl8n
8gbinGWh9W8bduPa1EBnbBbdq2YkVo9B+UFiT/uiUhdIEXFFagz3VHi1JTUuanW7
ypCyCVH5FXes2nuUauUdbtVM3VXft4ERtwEscXqjgzL2KSinrILZW4/ycwLlPRPe
XBZ77uM9CIqSj4rXvDA3r9kozHqxoFUNG1DdGvazffFLMx1nT0Bv+66znKa0lyVk
3rFN+dYyxk1u8+kl2k7MJm4X/1jFCHszsNu+Tkyo2qF28xmKU8GEU034fMfw1azz
W7n/5+xMkxBmrsjk69CeG6qKAw1ZkcFOqBxe3tIqkxys4UybJrbNGrY2hfvdeyRQ
3c/jKeELw5aM59nzZPzvLu1fOsQ5MiwLCXfcuSHueW1PDjI9Vx1pbERer4iYsI7p
lEV2eN0fmtHs+6avjSstnH/NmTL40kuYsKuM9sgJNKKZ+2JWszn80UqiCtcGo7UP
3G2Xd4U5kuIslPzwW3O660FcxDxYwUgdMVWyVH3KtF4P4a17rDFs3Jxe+cCmeHKI
XVyp8q7uFk77ZXvPOpnWZFN6Jjiit+Kkzyc5OMAtD1HOwprjmelDno7dloYCBp2K
71Rj8tnWqUKJd/Rd7NruOvMBB0kJTZydazc/cWq3h/bxpquhPHyQnUY9ZDSoDcDz
REvCz3gFkSHiggCnxfhvJAi8o0KzKDA0YKIj/JfUWfBN/4bJUDFnebvBFXcjmTpD
DAtG6et/s5eUQ5A2riRJN0RarsC+Q92mBdm4eWrVzU5YhMUJk1GmjT5XrX1nntM9
Tfyq2UBTVgK0Obc5ELawrJ7jQP2/N+jAwIb3BoCmKgHN7HcW9LyPpNaE0Ui7Hh11
+Xvb3TjdO9RBVjPdQ/caXGdLHU8m+mGnYOXqvx7bTZ0rJOJ5/JTyQW5mw6BWQ6Er
SeoPMhcfAZGUza+lQzg25Q7f8aWVS0w+71xmkP8PXpDTVtiO5l8UI+kmhF1zYHC5
OUnk5844Ak96J8GygU87RdIh4eVmBOyYwBHssPDKk0fRAzVOlbwg/sOgSIybApQ8
wWLr5bG/uhbU8ZPhvmVMyEMd9GSMvfxBYY64X0hxJor+t/KqcOlFW9iDWEtFUoa6
5PgdOUmZpf+wMb8hNq16oQoGnoyjlDs5H2l6rypr0AgKQdMo+NpLEmYMhS9eqfYo
+SnHz9/ntV6GSNsYa1U1so31Ke5AED08BSV8hFoqNzKs6Q+omxeGgg67tKmPHckP
8fAv2i0vxvGKh6G5S/c1062r2qT6cZoycu8Ux55N0IC0Hy44td6N0x2AZ03r6/q9
8pe+wAsI3ElL2PvLu6h0xFwr62gNHoeGbe4Fqp27etNyUjhZTVWExVKQvZz7TxW9
uxp/mOGI8BQDnkvG60oP5CM3DHKIRxbpEQPqVAKw1oX/DorUiHnHt5RVJePvM1/K
8U7r72q6pxQmxdbQatvjkc9+rC39Ql0yzDFK3jguU/pB8eKvwsSvhJpDRdI4uILz
E3okcFSaZeT7eghhGQrpB8NoW10BbwJZKmgS1Cv1wBsE7i9zug656BMSn6EHRtzO
SZgP7GEQxXEI8jZq8Oh+hW+k7WxcSTEDc4SeVdTm7eq5Ujl2OlYuCMn09tyMXQd4
sdKjIsmtJU4XjPowtmLczwQRILWyr/AqedkEID9VA64aE52pWzxUoYZM6eupb2lH
lUtzG9xgZgEWkbYxI4Q2ihSAuclAHDoY4uH+J9inFSReVYOPKAAaw3G9duFDDp+v
7IoJQdtL1EkSxwTJio9rhmNaVdU8Y9sMoeoxIvtnO4qxtwAxvxwnrtxp7EDkXrtY
UgMY9myEqa1+tUD0hI90XJzpo8ZbT7GEBT+QNOb2KlCv7hkflMzzPGGb2K105/tA
259T+2pJZR+bQ6HgK7pLhHF5Musf9ElfNKplS9EbGhjziK2dtJkLYv1EyzhJVJ+g
jjr4x7C9dBqErmtrJ88dJbd0zh0ut0aCTwFWEpcuNyiVlZKTp0xAOq7pLs46GJbQ
/g01XNvqimwlO/C4ahSoYdfDPtvLhsnmP1+KXDNdJrbSaRn+h7Q2YuoG/GhV9TVW
mLl2A9CK+IgJDzNLEyrMn6NWO8t1KyEVHY1zPq+J1xVhsEBnSSO9S4h6SpN++Pem
WaKLJk3zPo7xBsp465GQLEfda+nmX7ofwxxRAmTFako7AYZNNecmcEofwxoULeMq
2MoejfFTNYDcnRHxNIvrs8/ca4DYhF8pV9oIuPMwW0mfaSykj8i+3DfV2kmS2rOO
Vd5MVXP1K7tX9LQUY/lDt9d3oY+07a3gdjzpy9WQDi31I0pYC36DHIA2yk5GkDGt
3csTBwCKfeY8eOb8otQiqexh55sogPQKNjXqlrc40c/kY0Fj6OPMkAug2uL8bDVM
+9QCH9WpYb2LeW/VF1Bnr62/zmx+914upAjos46TsxOV6d1hga5UQ93WUQu7EaIK
B3huIUIGDtqDrN3sA3W4D+SAqgzWsj3WiVTibdmTMKI3bVbTj90Nu9hZJMmqnOZo
//ZFI8wufUDbgHvt/XNW0ZghFposm8m3XdiVSfYFOoVXa2ID0elWw2lcSEKT2Ftn
6NGcWOY1Kg9MZvCCa0H3S6dzyvLvZE5nSpksDEqxgssWQN/wNEW9xgmZYTo3mDU8
fiZQZNeUi5VqVJHH/gwwhqbERBZXrM/RfYVycR52//zDfv08z4YrwB5FNS6cxKff
Lp1tQoFRbYOG88tznIj4FlKCThCrw3OJzJ/gosJ7Zqqb0kJXcQRN51eAxU2d4I3Q
xc1AwAmUjW1gVBGibBFcEsVVKL3z9MthdLCXW+hzK/EBNDoJwUckYRYZmr9HrHX0
wPN7LpVIZcPAvLIN44G+8pXSUwUliSkwFxknggJDG1eCGUgPGBxCC1oVW8mzxuHH
Yy6DVW6A0ZMYL4ULGkYRlVwgkrUgtlENavs4iGFznIXeEKyI+bIGfQ3QPyCyuGHW
NKo1qtryZdaWmN1fLrmdYwrdl+vPnCnrSotBTZrllVHGLPLceIXwWaVqAKyyc/mz
aUGSNL33Vd6OUWo+0wiYBoQ88sGJcgcT47U/k9wBzvOHLOLFgCbV9e+ix+RWi0xd
oexy6JDcKMLDvhHuvrfZf05UGC23mnFPCOUavX5m3gcduuzNa11X44KQmGbNZ1Bb
V2nDkM+Q3C0ZObvUEBgOUDmoAK8C0Vt1z7hd4SlvtxXUSFEdYFNKDuBsl+Hy8WqL
t4BnVEzUL24JLnCtBhgSlnEANE8G+AHg00uGTf3hv+W8cAK5KjgQSJiMPExwEf8V
Wie9UI9x+3XACQiGwUG28tiZ6kgy4KGR5/94pdmnqRpVRxX9rS1WlKtAT+Km6fEw
FTkODnvUBJhwcTGAoG3VN8UOACLFcP7bV+sKK6jnQPWmS1mH8HXdMMv3JuZ7C26Q
WjmLStcUGQZEO67vi1nUdUutEbS6MNyGezUgF6xK/ZLYP7JS26Slkl5CB3FFLhXj
W9//CMhag++EyVZgbCrQdRtBykkAM446SOzhg6WojOSlxlYT8FE1yqqxjQcrHz6C
GpND3behveH85pJjnhhk+EfDdbDX2LNwK3tfahHEDLq9xZyJFQDbF/wYTLW8bpIk
SUFKyb073ssj6TlgoUSDlqjwRFQ6fMy08FXJEhYUDcYzdhYyI2Rdkqk3Hfk90KGn
k6tAzgSvLbaaGLOfpgKS0c/FOeyRMlhiNELbLRZfnNFkGHQSrZeACpTD5rYp6Coc
g0+sXaxtyJALyl31qgxQ86imn1gmEz/z092SpxMqR5Bw85rwiENTMcKbajsuoPsT
XqCSzLp2MDJaly3tzwFLe/El7YTRZMY+t2RNghvsexywWl9l3Niucs2GjkdzaAax
+TYFhgBUSL9wl9QfOt3MYlmQZM38sGCnLcAeANg5U1/Qu9R5wVPHGUbu77RKhnu9
1LOv1V+P0GFyVN2Za+QDUDwzC9kq3CJB2YJ2rv0eG6VIEgMbVssq8MAPkIATCgrb
K9kX2Wnul1W7u1EI95dbNTBGHUTF6XhlStI2E5GVPccj3YzGCI37LxQRKmaRJPIW
lxVHSX9GQ3uauN90oHRxnxnSMuCAGJKpnCDCB4KmzSg8GTPdXGqMcVIOEC4B+kme
72hjwKpd+tNta6lG8mN32HdIgoI2T+vu9HGUJu/lpKoozVFT1meJtpaEfBmmIChm
i7sWzrqZxUCZtlaUAUzAcGkYpcuMhboYZ8Y89T/ZQQ/BCf97NW0MPtVb7RCw4xM/
upUqARRG9O53sKLjtErKK6hGOCVPpV1An32i+DVLufn6oJEzEgUFnYOeHWcMHkWb
1e2tgTKn1hl3YjywAoaa3MVKlw+InhjfONKRIR6UJuqFHqimVQ6xyPnFrxkLzFwn
o4KYvG4eVGs7IvJn3nF9r7bTi2ppm0WZm+a1KuJLyXaAbTctT+YZdshMQvkAHFMg
ORYH7tpFqI7H6Yn4UbmygeUxqKHWQxXJXAKh9cOtvJDkytGbab1uihn02yMQSglA
tWv3Tza4wWoti8tqUSu0ed5j35YYRalNZnrZsIYOQ1xRkHBGcAudOR8O1TVCAY4C
pvdoJ6pktzddw0SNZF9fjpTjy8VKtHm18PW31BpzZNGgxwxedWnidbe4/aTIdFjs
GwzxrWq+DweXOrytOotChfnaU5dD6d/EC9jawboMDexYDtZkljFuXUZkyY75vp87
g0uuSWRxBA0co1avWozHWks9M2KS54FI0j+WHQuECkLh8vZZSnCQ2m61Ki2AYddr
XcxfFxGUpZPui6g1S7soimWCxbUKDBV9wY0or0at9vxn08/I69hTd+jMFN10YdsP
be6htClFHXTGpJvnwxUjhwe/iR357Wg08G61BMENIAvczyQj2z0h/sFIdEwcDVoc
VD9GiE206A/mfKpnk3NXzkRe+fq0iLZQKDR6ctsjOKfIslYQ2pfg3I4HltaJ4Sjf
rDJOzr1iXJ0TwWNV2Z+1aDYo3DjU5sDKQPR/MuViRuWUHXyma9VacbANHshVStA/
KGRi4qQlueUb94XykRTHorQcgsGNkhu0XYgFwNMp03Hm+5rccFbe3P/2t+XXTMzh
wGQlHwUVkmGazUILSgRYLBvEvBii6fizycsH9IutR3LvS1tszRM5jA7GDtkUprs3
hYbNPXU97mKM06fxGaFkW2WV8HLaKr/vWvm28nObx7BTKtHoe9YBbA/3BePyaEaA
GPjyhGq8nasqFtwJtAbMzEBLBoi9TpJO2itsMPDftBUlJaqe4VbsNpHfvF31D/Ln
h1ectfiWUsp8i8DtbrmXje/4LLJaZoTDHiwsqLrR03Pxp3PvmfRaPHdhKzw4Io5Z
hpDuNXDfEDRj6832MNrNGwv20t9Is1ld+oV/Gr3KM/TBqEN3uyQhHHRKWFGvCtbB
6YKT3+hbvk6nwlEwsHzR/jbKsKZdfkOesXoDFoVUEnJZdY8H86KypnweBwWQ7xZb
upQHBcxckq1Xiqx9IIuBiAzH3sT/KV8NvYJVh3e2uKPJy0nY6IbEwoyRNj+urQTH
u7wwsLwhcIIiGfQrhueCdbNKPRrQCozZTQYe4El5f0SzNq/jznaGTBULrjP0OH1m
MSd2UB6mORwTRV1rdInv4wICoVY+Q5G+ufeGSkyzokNf2kPCXW/BFy1QUnttLL+j
GIieBbId4Pv4+8jy5UVxVrVfukaCylX5XvScKGGwImTIGSJlabDmwUVtE8Bl3zDi
mCq5UqX4sTwsOLVKVl4X8MuMNwwcdTpENkF0Q/olQSdTUqiLuvxl4lBF+yp3Nzp2
NmRPF/v8BMO8bShNzZvSx4CMUFkkb1MMXXpLSZdR/SU/+oCrIX9NkWG8Ou3nLXuA
gIlvVGwtCEggXE/2IiDum0SoQLRo9XFpQrSD7V7OH4Or7zMOR/MVdMo2Nu/1y80m
zsb7d4NddUcDdkKERYJi7Li8MTPCsTtOGDTWKRvOyMOWtdN+6TybyQ3eW6Tbma6M
0g2Ac+EHp9wmnfVQBBWH2ZjvCAtXpoeB6GYsCA/VdOrNTAhVSUzhIccstFs+omr8
z/Rq1dr2xQJPKXhTvsgwf2PrZ7D/9mrwhmjhzKRAG5M9ZEfcuYyk8atp71qI5uHD
ZjMr8d+kMAttp9SPRx4EW66IriJ2xSq2kLLP8SGZzYV5is0ioyOMVcSQAdyT6hZ4
BNXGPYTx09CL/3OAIC9Mi4PBZ/NCw/qjs5rsSEIIjjs5t3MpfzTnEnfDoDoqKPI3
KN5JBfGH1pNZ1SAeRE+dfNabTghudseJZchFFar8RuHz3HyloJU2QXPRPyVGz6yC
EclFatIe+8a+Vkgwe4fy4pZy1/kEI8H+iEfeqHs3SIL3Mfm4CO/Nn7iER426x0PM
NhfCcwLDGajys9fK7p56TO5UYHg0F8ST4iq6wzXAIcE5AFGlZCNT3iXHXI7ytNb1
jEPl8phhhyBLJxZHldiNhd8KIoabbJqqfZ83mpSVJBvUdXgV69T6qTh/uzgh190/
Z+SuW5wXhnc+5LSldc/5mCs4cwUX2BMQp56mtv2YUi7zSyrrHJa14zyo8EdjAQek
UojLS+Hlbl7DSlqQjRxSDwBDpQyQZoAgemOQ/364Ed3mleYzZxa7UEs1iXbv+xk/
kyxr1v8rlZ0R03D8w7I0n9QTQLvPS0y9eqnHAvuxPq5IXd3KUExUscgvqy5Am23i
ZZ98pnPatrLAaOz8jrujoOrfHz9wgPU24Q2E2Dy5Xfv1TbFdiZjnhSCvTllCTHo/
7PLfByKTr4JcVdobw53dO9losf3DO2MFQ4ZOCPK/yafwWV7Quqeg9s9ce5BEIok7
AF9mKRX5DZe1yH12xmXZQkkyHGwfiY6DGFPfIGyprluY7GZiC5ToVakX3Gaa88MA
9fiAGiJ+TMDnOuv31Mp7fWvjlFvkXovG+B/UGPzrNigVjk0RgB7+xvEqqnNJK89c
tZZzfCL3o3rI5RdarfsB++/TDM0QWkn1n0ZXuQDMownOCdmqfAxpgb2h7gHKmUK4
iSKnQTmVJiyMVcA6uephuGHFG7VVta0tzLgs74Mz07aHIXjWNkTzXI6ZOMziy70c
bSgwL/eOzb+3uD4PoQ128iew1tjO/F3UFodr5rDZIjEH0fnQSg/bzmlkPjCUrFSn
e8nl9vt/W1StJJJkHX0iskl95hxtvkHm/fY1R/NVYV/tjcHXx4JsCWfzmzmpEgLH
AEibM2EnMqfE/ZAcm/KExJYflxjpuPRLcmt3i9cltSDz5PP1tXGP++68fmal1puZ
aa2T1p/AqHxIu75pkMMcP8mDddYs4SJH3o26F1pjRFPX24a6CzS+3Hy787D+K6RM
CU+kKlPLSs2+xfJVMiX1vDlpGep6+cymrdZ7h83v6Tq3dEjCdeCMubGuFTjH/KTK
d0o926BMzTUxn3prHtQe8cWcfWfXFZiAUrtMA1sDtH0q6aU53gqOU4R1lR/PkSeW
WjT0vBGc2E4y83A21aabSFakA6xMJUyFoWz6Pvz68/ZWT67YBeJdvMi3cE7UE2Pe
aX9ZUyOQb1Rn7dBon4h7LCz4WmSA4itfwWhqfnIpy1urYAjszkyNqaSvgHirtqqX
9jGGufbnQjbqQyFdcjaR3nh3rnl5h7kr8pAmq2z9NhHYBvyS3imp6SgsDY9V4a+z
9Tcd9L0asSaW8YdENdDsJ4UeW9FD2mV6DLiTzwyf9LjlTLzO1HX9aF0PzDqRCfLc
nOD9odzNN4fh9CqR2ligfqiZgg/507hd1qvFyq3swOic0vYpR9iexJGRBaBFupig
bFMRSVitWMU2dNGNrT4QNqhr3qJO++a9JyuB6UUijhBODxPzKgFyQNzT0mHWsa75
axLPrnMq5hqZ6PBFgnQx7FYbbnisidE2rAzPCDRvxMDlm+lXXQkSy9u0Wu32MUsw
hZ/ZN8mUssqMVEuLxFJY88ZkOv0+yJfscl8Z+DolAn86YEpgZ+7uxn4k0cadq0Xb
OXeZZRqntjfXSac2cQYLQOrKHyFbjhBcMfFGMZTidpFWEJBdyMVWJySbdHDlZc7f
+pWYrOyLsHWXg5iwuvfuKom2lpfWtnrT1VQpgMKdwuV+Px1q1ebqtHk3qnjes0MZ
C2/UhWV3VoBa3Fgt1RqYVSszQ68UowWbxEc6CGP4p/nFDsLtiL5xQXeo5RzKVL5x
yUmd0dhkhMpZYoIQrlMLTsgWQAAwDuCNzZNacwRLXBXhPtUJIFxYXP9973bIF2gv
2SagrqH59ttxf2amSYlTnUnNhFJtdW1LzA/vADqoMkR2s7UJhHPCV8RP9sJ3xMMd
fWJxCfr0vCt+oJDts1S/6OXlz0+Nw3rnpKm3BqAWEJ/i1VjjsqotkPLq6SFsM6Zj
m4b3C100eoFziEHQOdMFlbth9qvLUvfr5SyDZ4nBvQ3XCqVHDwzfmQ323D7EizZT
FgSWLvJW4Of/LJQO40yV21x/oEc3Aq6+WCOb8ClPX4pBE++4Cu0MIKbgNi1bOlRC
pdtY9KSqFoqzCykjKNK+VgvIZGB4CZkDl/r65yXtN8Cw0d2KXKInjYAKeB/r0uv+
TkI6+8XMQ/O8L6Q3UDmq7JbWSbZWZeCQjsKXutTfRp3X9F39ox9V53Wmpo84FqzV
Bh04p+DsyIp4h9wpVRaAb81VEVP+DlQ3fyeSKEvTSf2fbe0DfnLBMYTwrWhGzYuQ
plmfSlWY1yt2GNDuqyK94LeqTzLCiC9HERGscAIW6JLaUPUwHWWzUaiI3FjuKZ1A
4MLw8Hmm/N2nD/5PbzuG08yCTNQGlegx8eG6MW9PYqREZk9DPJ84CYRKbDhrYXco
zslL3o7sIW3P1SE5NSKmpm29JzPwd51cwc6HRoC4XCs8Tr1+aD6i2GtYs7isbHQ3
qG+Ttq7JbBNVJQndbofnks0iRdCHle9haLfi9JwP4/CAugAVOkB7y/nfXzTPPHg/
VOpXboUNXeWvnaP+KLtWmUDu/hLfDuh1YlYCpBgR0JamHTmTq1acLhmzT59Xc9rE
qImohRyG2UBKStzBUcN/flQhorLDfxilOYxElQg2bqMzSQRprh1nuVdFLDU7tPsg
Ih/TJMSnF8JZ3QlWA33YbngdriLQ1uV+dtWo5KdLozDeYECslo2XRD9Jc12XOdFh
+CVx+d8IzA8PAphtWAd7mrGxKvvGHMELFjXwgEGp3fLdcBxoUxHnkR/CRaEJXWYN
/jjsokUxN+zeVW1jNSu116brWGyuRblQvrDMEk8tOAJfVf5QJrCHzjJq9DaeI1th
Y+UyWPdfzgPvTm89wihCQHqtg+VTE0nqlSscMzynH6CJ52OhdeSctImvq3vdlmws
y3La6xxjt2epHXNTPbhHQCBCv73T8dg8hZkT/0ibOTPgZWYYiEijDAw3in/RdSAi
9FlzaygFCjGS3FhorU3l7SB+E/kHe4v2Mxr5t1ik8mBFsHCM2gc4NMf4aIc7NOBZ
zB5oLnuYtpUUC5L1qjUOCbMTwPKzt1cAq718u+upqEQA3/i8B3v/BSZyFKwkGN9o
2lcCtU2gp0vMOIbpsTFwPA2EqQgwwYVafEzobLLC5RuvbGJiSGMEzNyTIlNzjnV9
i9b6N3BOYAnpc/6ObIkCOniMYib9+h38XCVeG0/3olHs9z2JK+sfD0J9BLInms03
dnhQFiJ1Wr4cXP5rnn94A4JYgjYZfYPVNHuudEbkcwbbvJxa/P2iyqa4h0juRfnN
6PdkqcOK0FtXLLNLSFKg5qgzq5/DTwe50tI/tMDXRu8MiJxHVBiCQrmH0tyBdzJV
R64Mg2MVfBWQNW3PV7tnSYxQYkKpqQtj+8Pp8TkvRiutjQA5GO7L8FC+TH3AdP7h
Jja5J6BtrtHHtBA1gcT09A2uD16VLjz7j6El/+rdVWaXcx+gykU2lppa1dGF4NPH
Loj+tCpAGME0XMzOqT/0hGtvVhfWhuLCA419/AEeLwEU1xP5QzZHZpaBh9Q0uPT3
VNbRca6PBdYMrNxUpweqKG7O7HVtjQU71C5cbkcBfUVwdFFyDZMWMZDVJ3+zKnzB
vL8ijNgXqgqIcyl23zCRQQ92LXxDP75+jQj7aLcJXVsX9z8RFFhVLt8+MuR7Iuju
+7b2TqthA8tggAI8T/NxV2Wfhhqdla7+wTs+bDi3p1YpljmJ1S62jc9ON4mypRbf
DK9HGg6ajsu8BujbQpyAseEKZZasoFStTuZzJ34cfGEq595VHmSiJseTuf16G97D
85xl/t9yNHXJithWuSX4W0z0Ahhhfs3JAXa2ZokvjmZ8Fl3yyrryLOtgEVulZ6mK
87G1O4iHNdtPQexZ9pq6iIphgRp5Q03ton+gLBVOj4sEqU0fdrVtkkwpE7dkE0QJ
ucuBFobsMcQ9FgO4LAUQentFVwxgvpiSZpTsj4lii1WmrWQIR+7IG2fukh64Cnuu
VPFZ1M871sZN+uGdIZP6sQBQzyQeau9wpJ3VNddegA18Je7uU+aAmLgkx2i86yNx
X7P9gbJJckFExO7RTsTXBSsrxm1Qc9zXRdpW9R9vYcCf1fqnmeWU8az3tUOLYV4P
VT1ABRQNuYZGZCeEQ+oZ2zCcSmlSihE0GgFJ5ha37bDB4ft+SmMJJqI2HJF6Fwvo
n9edTco48xhBwp4rNw5L1Fdrhry0FIM3V/AFMWwtnJOwe4dF6FVUNT5lRQ9YSJ/4
qWRI4J0WKJilQN+NPv2hAKI/n4Y2ELRtz8teYYOKUM2h/wmZIWY33V2A91W01bS7
HRZgv23QS+gtIcC8ZDRzdjSHkLNzMG1x1lH/tsScNGl1X9slhQv+f1AwuUh9W1cy
QIwXc/KLQklw/RLW1M8zCefk8qkjs9bkPXv6VeWyJYuPXodagxpSSj1IQ5Sah+LF
XPzcmBTMxQN8JsST3NkHybaW2SomiYnC8yIpK5ovPEzLbXC2WpFFigo1vfCHU1nP
ZsEbFszn4tDezK2IQugHgdV+VY/EC5lOnUw/4iiiyq8KypzRiCot6J5ijGbX/qgV
kqq+cW2JLAUTLat6H7DPzVshGY+3+ggU2Zn6qwy7E8x/q2GsXkQAZFx+71NTTnXT
WpdfqISXHEfihd8FYgE1jTTRLClSnS0L6lt9ttr5l3a/1mX/aIUwUVNaW9pv22qh
dWD6Oh9qWmjaIejjNTweKVreCzB9BASppzBjHvpuqymkOjR9JImJMbvPzmu0dRK1
5pudrOw1mfdQeX2dhUyjjsDrR8D4k/YWw7AovKAgIVimZOAxKl1qQ7KzU8UfFpW9
gUKnnWCh1FlNA6OW4qUFPiAk4MuY+siGAWYoP86IFJ4VCcGWAT+AIkkOKgBLlFRy
kXWpKtnqjijxt2yWZ8ULyMtrX1HHqA9mkYXPne8JaBwWcO5KxVIbw3L/emaFzK2X
tNZPUeV8Nv/eB16Dl/gjlJjPQePzJvEp8mOu+5dAbqS5JXqYHoX65NmuZWgYDe5r
12mgGIVNOqpube3dkxHkbTnh3U/gs6XMWh0hQp0BlhrV/ZBNZVdLR3Ft2E6/Jg2j
q8e8nxxZHQs+BhEx+s3/ZKMvxgUTvQLNOo7xxD3YX/IHN1N6+FnnhQA1fRQhrbpF
sbpdV9qP7Wr5T8tQP2xGXuZS/Kl4xQhgbE+Yf02EWYQZeoZeBeVFqQg4cfHpFyOy
QdaTJUXvxbOKezV1eLlPmE9isrczdnIdQbrvAMJ6hSD2+VOtGhimHKjQmAo7IGNZ
ZlEabYpxJ92VKadQDa/ORqv+e+2aShkfii9eec4Vs/zS/vJa3FFdCWbCyWmr+via
sV+MCxLbGFunk2ZO3oz4l+0fYefkEoGww1c9a4XwfrL0+Z3VQaHeBHbKgeSqb9Gd
bmJ0ubzXFd1YVs5CQt2LpquJIw6D+YMmoq8fXmkB9MeV8NWfojGrpPC5w+8EZyYF
G8dGMGpuUCdlQlK0exoilvdJsupu6aNf6KRk4BAGfBgUvAYLzISTXsKPMWfGAMUY
hDTu5C7aZlFeY9u6FTGLjE0Fzpm2kbuxfNvLWOh530N4N8+x4wz7Nhf/NH/45WXf
V5JgH61BtWIdKfAZufG5fQjL4zbQ+A7naKKcYCxpxOBjtrgkd50ealv8+mcivZGK
gtBs09HZyu7a06+BfxqyNf8ADt5g+gsGXHWDMyEcMN/Q1bsM+NkHWXt/t6lOPGuC
AQzH5rvaT1a2mqzXfDooO3UZajTwVzTAm7JhwjCzM9MSC2DgWFkWeNHqLcFdskrG
nnE/jOd4tQVPJaLJ+0Rn05LsZTViZ+1hlpPtjn3Nu5FP0kDGngwqz5B6Jk2mwcJa
Xh1oVQCbHy19KJ7RnmbcSTy8VXtw7uI1Gatxyax/4fU641sDkAbj6Lvba6oSSLzD
7+p6aW6E7U7v5cKGdAu5ssnZ2mVN15RPJNcAiZDdzAKEQbKF97j8VZvOayJfCyUa
/eY17sIUBKAau09MT14CcpYpaU2+OJrbkK7VyeMIxKmcIxpElpXOIKvjGuAgh7YI
URNtAH0gEQsCleyXtPQPC8ApOhJM4MkvV5bCArnRVST3nsXRM0sF62vzIQqXQxo6
1DRNaH3WeDC/fnGWDbTf5OCg0NWkSVUpdVmTmZbNqflSwFa6jSw9XPPs0KnA5Syk
zrVaDE8WazFKalp1ThnHJAnHqNfSlS2pd5vdboQCult6P0mpfzAh2eDjoGaKHP31
XnMsyS1p9KaWt+w5VvUIrWU8wSxPhh4yGskbvfqPSJTmRlUkA5THnljqi+hWXgFr
+jcubr1sy5/23h/bUxhP5Hz1JldLa0beI8n+WZOF7lz0ViUn17dnHborHlPdpIFy
ee7SK4ymzyZsbWmWvX/H6ALg6d1OYopDg3+Yyw1PsrAAyreAnSQ7mPmH0QGHw0PU
nbTCYgjExkELVTAU0z4wUTVyksv/ypS0fFrQy0mHHe88naMctIPVvhmZA2pnoRhj
1015S1SKq12kc6939sw5Waf7HYcpKljOCwYOUESRZaUvEKx5Y9T1ttq/br51yfWU
EqIOuCi2Ubw+U0mH3rPw2YtFnFMkObUDocskqFa78JN7kTswQTzRNh/6US7Bfacd
1++6T3xJi2QYj5hGHPpo9gh49+jxpcl7w7E5z1IfCIeUMav0DbeYz+tA077UJR5p
bHO+rYVMmdYdvSLGOEpMTIYC4xrB7zIhfkeW77IZr3SbYim9xo3JVN03o8hIdGr1
BoMPjjpB3wSSSdluZTI5a+CNmuwcZ4AgivDErkF0AuOCpbvZYHUkJp/bVU2wzZJ0
GGmV5Ue+b0EYUknYWkMMaaLyF6Wjx3B8PJuLll895jJs4tLsue+A+lBLV2UHRZOi
7A93JNExD+LtvQLCoPnbE+If3wyDUtf/MKOA9M2BM1WvcZA/ToDm/Qx29qqW2+BZ
996PYPvRRPvXcLbtWdT7CroVdYO3EF8Jc1fjzxD5jXmJVgA3qJk0nYnlYm1doU6+
ToKgYfAuMUzKwcAJMVfpqDbr8R3GFmh4n+CQUVQ3IR2VnWhCaYCFOrLTn4BQ2Bf0
Z7F7J69r1Y3dL8M48LmXq5/qYnUxOAtL5dkFu1BYGsyEbY3JlEzL7L0jAN13pLBl
cl2HXcjj/hYEYfVoJyiUf0EWmwIMGL60nhpTPxP+uLF/BEDJZAuxoyy67vrJ6o3U
62Nf69WsKm0h1qH5U8FOozfzqDbI0CVUaXdv4sHFUgIf3iW73w4H42pSc9BxxEo6
iCxXbC510S8vXGnziRJ2haOeKcXT6Jn/6lHH9pXUZ4z3O0vQ5/5RjnbTKPSFZ0rs
a/BzJMV4Tee7hRiXlHvOmyzjiJQeIeFP7s93vG3dsLFeFvxdBNdlkDzy1Ho2FZoa
ObH8DT975aW6HDwbGl7Yt85h/ZP5bYO8X35Ra1exEMGrQUqpEay81Kx6mAvVqL4z
7YyqqloQuX0xcHDFDnDujAJpgExZALlyvlH3homROHkv6LzVoAFeQAtshNmmqI73
U6WzHIgGcUEBdAaI7/NIG0uUJ4ThIwAbaqUmh/DYL0048YszhS+uiFqBwYyOc2ql
c8tOTjUoeDDkDEsxkKHBeEwAuSAGhvT2GEYc/+ObhXy7KtOzSg9Xv1FpsnjbgRNB
AdbR1/CdO4wOXlurkH+tWrBPfXUqrdqcMoXrvysYaAN7sI7HfQONLasaIav07tv7
nmOaDWm7e0jN2qcbIduXUozely2bUKAZaRdPU/TEUbuiE9YpkfmNWSCEcd8Wparn
6eYG3KbfYzsYFmwB95kK3kd0bxv04MtjwJxpBEcp+cvKVt6bVVIjUqRuY/h0rmoH
uPAB7XYKVWj34qJDq9zQbGxMgtrR7/JbmNtEyHNK99J/brCPMCfaY2NGvje9Oi9Q
KNtp5qhoyG+gI+rOBaxYn9aAR7HSvh51Wi/Yd/08+Zv9RwGqKpsadQDlsiTSFlL4
YRwgjvJURCHeaYHkKfg23gbfTGEFVHMKqCjX+kweFzkiIgGy2I/K6zFo3/FE6tmS
Yqpe0+vNDsJAWug60ZCMJ9ok7YsPnhZVzix1B7N6mXsU1v63Vb/fI6NMI1YToyBq
wKPsuQWj5guKGCb0SEtbfP9jC72BUr3FI3d6/WC6DHTkneE8HVxBijrVwbFhYCHE
o3D8TvmHT4FJFW0IBzNU2GVeuAFKMhhz6GeZnXnRXwOSTXn4Ki71JqS7BQCrGqqx
JL0a2uBrYfBT+71SvIdPHaYqUj/gucWZF9BK0l9v6dGPXTvA+fI3Y6xdgUApaooG
23RjRp4FJYcc8xLneR6qmYqVOZ4iPIVyj2NAX7NdpHFsx5govqkbjkWM8PHHibYl
HY+WO5hDPwgQqV1xkGLc4EPkr68MghMhwu05w66jfRQZILK/KX5bUb7ECMsrmcyy
PXa/tYzwfWRqg/rXfX4Tift1ZqpX6/Hva/ZkpqFXE03CcmCBX3msLm/GtgqD6iSq
MEJdYyxLBFHG35E8tZ2VfbW6Up149+OH6Gv7EEAtghuSTw3gaCuxiKxazTZfURe1
Mpi7OBDDGHerHCMh1MHAvnzZKiksUrrcYZ6c1zq1k3G9FSWbpv7t+3oFQbry3z/6
LN2rcfYBEvs8HQ0ybmwt8/pi5Z+uqjPUd5ZIUU0ioRqja+9XuQpVWNwfbjQTN0zG
tTEUYIHf21i7E1jyotI98B5+XplGcLlpv/+QtEaorVVx57cUpUI2yL8EshCJHm16
kryg0CV01WtYVijgBJCHyLxHFHsR2D7Gctn4J+VQvPTagf3pxLcaoJrYQ+0taby9
CaMLJ9fm8Eps8Tji1Yv8950EZn0ZpmwmaqGySy3KZnlcDkwb9gIyA4M2HqXFIyEa
gMvYadtzkuhVDLvPu5jOoNKl0iNfrB9qwS2HIz3rdk6WD2eAdgnhBh8D6GnlV/CG
mP2dFq8WoZsTp5vgIn0UP1v51rM//nzdbQYe7fu9Plq3Z6b9ZWiHecIiwKyrhYtR
1BukdQaQEM26ZOOavQ+UGFeBs4wAGBBHvCVcmbKqIR+O2n8sKdq34UfLEfbZhS2Q
oOKtwfq4RCsj7xycc0BALpmYkDjIVm57o8tOk44OVZelfFI59XbEdYJZIlng/QIA
TSGjdh8fIg4nqKTrPMtDrGgOtKPZR/LUHGPwsf0AMHR9xQQU9U0kEzlMh2IyV1NV
e7EoRHWxTetKiLpyAbB5rDaVpSJlm0nYPzVIuKPQHYPc1XnuDJPcxnsR1FgJRoW/
4/yJNVcmXJED3xYnvfvqxsOAzpWjIkO7AloW9TIPiIFao8R96Z6f73DN9wtq+BK0
nOCQ7zI4eIPOtIoeTSgzrsq32aRhCEQz2adxIMdX2jss1Qp6CUtz5Rxl735K6mpd
OwcltHDaN1HTcn4Nqqi4r4795wH3YZoK7pi+2PvvakACB/6MApFRULD5rnEdLP1Q
ttjKpWwtGuzl49wx5G7T6B2vkdxoG/D/+0zZV2UNfjWc2mZGGlzFgD9j6k8G4voQ
B2CwMQL3w/Pj3fp9PcyUBtSRef75zSlnR+bKgFFJUuGiUJzfu2kKdVgHynnCh6M2
kUNRbcUzjd8bWYAR1ayyyNTD2Ejwjy3djdOGP/9loVU0a+qSxJZ9wupsIedCXZEI
ctFMkRJVxWSC0fClqmvlKsuIvCMbC0NyQnHAqI1n55XWNTbk5hkaj7nU5PiQXuaS
5NEcKWsWj7iUKEf/nzV3HikiOR34OydPlsSppAcEu6mPx07aQ2xd8MYEyyqVBMZf
VJ4BFMvt1a5e/h4iTHPZ4uaA70KMOuy7n+j0rk246QNU9SmyIwsIJp+Iq6sO6+sv
4/cmkcF4qbAds2iDIlwYqNhaOc9LV9Ve7LwsLjSUNbiMsdBXPB+rOvteG65xD4tn
YilbHuD1Mje5wk3bgO9bfkp4EWgLXhGVzXvMgF2UI9o8WZ3Z5SVoOBXD3yApWt++
qMsXHJuZG9Y+z0EwMVjFRqkMPkZSMf3o3pFrqRs+Sw+MN18v+iWYizVZV8sWAGc5
EEFtfzKfdBP6RwxiESUaYpLv4Z+1biV5Ol2VuV2PObQSyub6hdijZjhvZ2jSHpjw
I7gcZqhH4GW9opjFZvU7P5wyXbtIMOxOXt1Y3y4SQyF8aw20698OjkLP/i36fEj+
wUiqWJm64vEJewRMUyZyVAlyFP4pO/wkmdPMEP0L/HCAb/ZL3x9f/YfG7+SzVdQY
u2yqtFPRmotK+SgEo5Bj2Aig3t+5GKy581pwQHWyC2IcX3uNLKFdZ5LSxvbxwZgY
F9STvF1atZi6Ob2JzkXQarclZMq89fD6W8fQYR1WA2iI3E7dT8n0AAz02i86Gg2w
PJ52rnCziBtZN+8RktE4HqAx0IqIGNByM3VpH9K2aOvld/V+x0sbRc49TwU4hEGa
dSKbARN8q2DOLbbFGK8S8T/lWvTaW4R3QryZ9W+QtTnz0bOvckWDmmr1Zk9PDDPm
BOS396Xq/5iDI1kLlJU6p33ax4za8cjT5OPWkRedGdMnIk4k1KKNygNiIUqAzxJ7
5Z11pacAyq9b+AQ/pAujD4jKM/5jWY0IIHq1hlfaRk/Hc75kgOT3oh7xWQuVJPBa
Rs4JLhBpyrVTkRos9tvQv0tAaVggQmtIVF+rvg1RVaoSVOtZETsN6gx0jBTbupAF
L2PryFcex8YnKKdazgs70/lfbbK1UrEISiGMDZcLIrvDBhYHtXR2d6PKam1wBa0w
fg5fs8XolSNcLSZhQxXvv5RmX+mYAg2tZkdh+RINA6rtRX6lSifks/EB8WDjLRhF
NdvCAoGTbaXcZljSAbG27AWMbtRf6uAN0T5Lb9pSgYP+1ysvqRHcIR/ktIReg09i
JRc+FtD4sC/Aum4r1rz3qX/B+tNw2QfUhQDh/Xr0rwrdSZIo3B1iF/Pp66ZNFx4q
ByY+ntDhSk3jAiPXdZ36gM54tHx2MP81EIJK7Yku0r1UKqK0nnIdSeCi9+d79xcE
m1n3B+J1r80lV/SUBN8Q7gtmIirIXbaA0Ijzk+Hkofq1lLErdhrPfy59wqmJFnVt
PlIn7w9tyG+fIyi18O6LhFkkb+znFy2OjRbfYUoEF8enKx6oQ1KE2gSrGTBNDNRH
7x3IQc6CzOiJmp06S/9ylOaLmOKXKufFY54wIHrT3V2Vbdcw4x0cDkFRHjahBbSD
32+JHEhigjT8gaw4PnbHSrQ6V8pCPS+/s3zjhgU+MoQgOL39y9Mqrf8UEBxdk9h0
kFFZ0l3qt7NrY+xLhMLJxa3qXFaOHqzzSmaq9e1+5vmnYGgIpsdVSFTWwy6rlBMJ
NFKurBV2OhdoLKUeAc10GaKVB2W9Nfr/85WPcueuPiLqSo+/8H5zYX98b7y4aQig
nwNnG1TIsa31WUtR6oNbOIChPJcbRkHW4doF9+UvbKNv65FWCahnEtoia6WvoNGE
XMXU1ZPsC7K4zeqt2F4anoYtLx2ZCH12+IIh0IN0hMAE+opyD5dK/hwDAGWBTjm/
4kSvGal+nEEoR8JPQZl4pQOqffr5WWykY71oPR/QumKWfak6/LM6Zk1Xpnsah6do
i6uGckspFxeiLruaka2XfF6YtSjSDgZTo1JwT4cYvI1OK5afSy+plQ7+1GXKW5Z/
r0zDamZczG33vctxDZcRNL6LFqBMoz2Gg0fOTypxvbOKv6IKYr2fZ4riJNNcsrZp
VdpD2fb59KWb6EF2w9QWanZCM6I8NGckQJiGKFj+bSISSvwEm361lzQNvjzYhUf6
CfF2N7QouIKMoFDmLohCLN9m9VW8owCvGHsqfg0U8c3NwvrRWUKXwBKQN+LoTlyH
WmhGjniTB0iuWG4iFMHHaZwBhE7DUlWPvyhPkfBqqbKjthN1nSGOkb5tVsx3DgX7
qJimAditHi2vLWeXIE9eg7jPJ7T9R5TFxF0uKSSu+RfIETF7UgjF6yE2UVKQIJ1T
QJ4O9hn8WejYaWd6cstWT/+NG6yV5ez7OD+cwogJllFd1Ifd2TIsWSy+MofmbYkw
EM4Ov/FiwW9fXGTPNHgOGnrK8FcyxDSH7TKfbD5rousfFhrKIZ+vJIiHNc9zsqGZ
NFKZLN6jueDCyUIaqcOzACbRC0s1a6AA8SKNg1TtqEOT6WiVNf90e09e9QfqfYrD
klLFq5daJqhB5au4pfz0VcpT0ifMYl7nMRUMZAc0YAdBcBxOm2h2YmuDYC/6z1jU
Smb5ZcDJtDJEJ4EL96FvQPSVVmvXdNYlGEm+NW7PEhyuRj2eJZP/kM+PALkS0OLs
9u4BY+aryaDOg7GrMQPpAvkS4+6mC+7JEMnkRXTVF0anddjX/cxJtTjcjnzuNO2B
59JvONftruQFZaF6DJ6gMT4u5J8CbSvugCC4Te5t8bAhp4A44lZii9yrM18i4zdV
0CEhW9n0EczA8nhqYMDdCYvoqyIfHHgkWwT5z/UmU43qboViFE27ADghm+85qrX0
3vJVn6dM4N6lwdB4r00hvEqGmFtOVBU35n4cdMPmHs9aDSJZkynAbGScRU/xr+19
AmV3TeIQ5ln/dlx1GJPFQOyNIZefLNn3WaTq8fjVD65j+RSzOiCNxf4J/5NZk4kR
k+hVCzu0glmdx7RhNkZh544VORuL2MNuYtY+r/o9qtzgPtm/ifwXLkdgEXg92znU
7kv7v77tT7j9xu1H25QjR818/vSPw0p1Rdh7qW8VUBJTo2X+5dV4OcPFSqDvM4+B
o5vH76RoHvAZLD5wukMwA7q++gJ5xgl6o7ZjdAXqv/+v4MX4xc8phwX+Hk3xXuW9
pE0Rt9At3Adkg/e68uvDutGllFl5PUF3b9p63+YewrXQk/rAnpoULJsJ6pvalXmN
N3ZIfQTClPghxwHCAi1hi2m7A0VaWgO092EGeF8dwzTh5ED0LNO9GXJf7Ta44X7m
N2ayMLuU70nDLBP9Z5H2Sdo2/9KA0ODMbyx+t3cl+EcJvY2DbJBs6QgovjokCDef
jr82IfZfva5jyC5HRfzHCGaVudYeJWZSYGxeWvxDnyG3ReIN+r/ItfrPmnq0yx71
AFkv2WQdq48k9wNgdYZ0qgCvu5kC957by+PYqZHVltsxLqmUVpPJ71VFgiZeuQ7B
KQ1FnwDIVMCmb51XCExgNKLRwWlaZDfJgNGMjtQj6F/TRPz1VSdxjmgkFuccpsA1
kGBjDdaJdDJfCUY82ihw1thn//s8YeQ1XxO9wzHB75tT2Ir/jwHhpTVUl9wBUARH
JSOQ/GD9oUEgjt+5pxhDIP4+f0mloFe5ZHiVaNCR4XIr3iIa9AECwYlElE7reKXv
oawsLAkQEM7aktklPyCHoYVC+Rpe14eBzsFNndfAuWZXwFacRI5rau0oKTzQGbOL
/4au/i/pEOaqRLpqomYVCe57HD+/i92GClzcvxnHcJ3PqGuZogpsFoikzcw5YWIK
TLf5Qn6SfXaYBgU2jEqvfBfPdfAXccnWZKRkGQxEmqzsz8B5+B56EMhCDn6UuVHS
oyMAcMHp0XHz2a/GBtHuvk/2Rt5Ijm1eTzeXNrH4/RC5TRcviAnSvcpUn8RoXkxx
m/SpjaoeJN8bg1WDa0mnxXWrKhIAJctiOFU+TlEqzEN9yb/6YBesfZMHJlShQEKy
i+hewtCGw29UCY8EVeSJUpIF7Tj1z0nNW2p8OvSt04+064sL03jNGKyu8B9eRuH8
x1eXmj4/X3S5Mdg/j6a57GFxVXyIl/FrB9/cYlACvM5M4WhV17bLZe/ZLh2GUWDe
dDCFUSEh9MtaxGgT4yis2sYEjRzaIDnXhIcv+mE8FTXCt5YT10tIr/G4e4FRpaTK
zjR4HtLjcZKaU8WnyMb7H7nKMgZZnyap7rzUtGcjZdWtfe7FR+qyV1Hm60nf0T4I
qvdw1nBk6fseH8zqzDUEudnyq6xIRfzj32MUByLDqp4r7rO96Jc4u8uNrASAF3Nq
zoa+DRMp8W6EVBgM6uQ5IiD0UiG6ObYlebV2U+tPEPpYBQYFbqfzYaeAKe1VH2Y6
1nB+PHkCq2RXGue3aUhqE7K8J3GdfkJu97KgakPERKYCG9KTxSWF4k8/D07eLnyA
awVDhS6fxywtCmcQ970ylt6Fm3ni0eh2U5LwS8Z3fYK0bzmNZIRZH+y4LZrvlBeG
R60dR/7P27GRkOGy2IqNCyWBYiF5UDpLMF8SQUdcwyPCCe+nhPDp5Vh4KuqnzIBB
i5bgC4YXy8Sq5BnvoYymXpO7hltIfxnuLegKwvo76mV60f0gpkwbXim/C1KZMmBK
Zv4Y7JbopQ+3MthV4CW2N1095KEqtFyIXwIYODm1HKM7TGfxhT1YIN3NvuPWJ5UR
zf1/qHT/cDC15tfViZnh9WnDpSrgBARrSB9LOw5gc7EGDNLNFtHKpMsTXb3tV64s
E5rhan3p7WhaReDV6CHx9scR9yFo7oeWc8Eb/3u8ZaCMnYuPVRcwhxavRZ7L2iW8
rBTjK9Ebw3eqmhXhzq8ed+oN8aR/OPT2kVE9KPTp/Cla4w8UoW6U0BDmCxm/Rhe2
l5jws6NNuzZpt/QKIFCOolRY/ttJgR7u2N5cbucRx3FwMNR5ffb+1FBwP5w7vrks
C213XkEEM4q5AlMOEez++Gxwj68GP1sAoOWvsMMfGZpBM6NGoyrckf4yWzeeXeAQ
qom7qPdIrIicJTMGcCq4828BY/8Cc8eVPVUEkEQp22/fGqQGGpOlVhrpC9TT4oZa
vcc8Yq4I0YGAtDcFdxt28g5QdfTx5iF4CMOADta3+G4jOppQi1VDdsPvVOLYbW2U
XD0cWfB8nGsZJiLOisG2TYYO0aCLmXPcA178ViQEtVpbBWK1j7jbyli9y1M2Cb9C
CQsApfgFhDq0ntrs5N6pJ+4Uuo/D19JgZKFXjizROqLi37y/i1DSFYSymkMG3c/u
HyPcUrPaZR9YsX6CvlhWfwWXfNYH+ce3hvZHsxfFZU9S9ev3vCJF9JnOe3RN3JOr
eZc8s+30ntV8lxrYwfamJFW8fuVEeN9f2he4JM/9P259coa6fyKDeQnC6mzQBnqZ
VyZ8fYOGKabnIGSNIAlet179mLI84H9OWuN+Gt2bJpTliPVVbQFmwOGvhGNe4SHS
9eKQCRH8rOKm/Hxdvl4QzPYk9xfw9hPokX2n+zmv5qNwEtFWn0GkcByr6e1KZpwM
jSab315WVOukgNWGejUIE+20XjTqtOQfQG9aVVdvTMyOWJPhVvUWM5Wjgi9VrAEQ
oc2nt2dG92/IvImCcLGvsCzdBgsKn2egYzvw/0GH1MndiK93f5CJYNVgjBjPQDxQ
PfDnUA1d0jkd4bTOw0o15QWVuKtrS6TkVTctaYUBWYWxVuk9tx5saX6Onv+pnbpw
/fS1raPhlYDFbct12DqmufUcsvOBST0dZADr1GAvjtHViEv2s7a1MjiS+I7XQiqr
eF26GyJL1U2afQlq86Qm7KCYK1KQ3zSTR7zKWzIoXHWBWrii6LA9ehn8yfoYNz/A
5NYEWo37kAwSdBLUK95E2VzOq/EeJJm5no9iYRv1WSLiuPzp75Lz6GjJ+PZZkUqe
c69+8VS5i/82/YjiDj2D6O5GnNnShX1UtTz9LRTwTM+oYAtxala2FCiVQm9L2KEU
pxqXuq4W6T+kr0SrU2aGUwxUHQA+2szR16Oaek958WCaweDx4nszUbrKna3q5QQP
0ZlsTgk+x2Tu5pr/h6NKWHenTPgFNORAglvF01Bq7Kffg4ud7udFgaPyCRnzSpFy
fHukSKZycqrlVwaGgWpp9D3/Vi7zL5Qo10GMFzvHplSPFxy1E4pHWAP/PXfh9FX6
1EO7lg9J8TVaHnIRB1WW29ZiKEHgKTfiJmJIztxk4WwAzCX7XCoFc4uV6uW08tJ4
irBMIakAyQz69Pnkwt72F81xeQq9k4kb/WDwA2cGiMl0Rhv9q/SleAU+SYyEZaAW
UebXeZvpqyGJ08Pc3RqzVXvM3ZFbxzgk6HkTtcbCeuP1Y7vvbDovXFo2nynM3vwR
VStFAPKKyHHLmp62IcNgoLh2Dd+vkCoAuaVODDm/ekjVNbowPo7grju9pvkqV7Ui
Nvz08lWcbczxSbQB//gFywP/nuf7cUnD/9ciC7Ttzwm3Cds0dGW7oZJQLbFbQ4Go
/5Bp0Q5IL5aTeZL6PVF6LBklcvpDPo/psc+E3H8mUa6zQEC6/iyep4FQ40Aa8/rR
o9NPJKBQ5MMoeoYzkWCk1ETCTkuygIcD1yikwySIQO7RVOD899XwZchqn07GOJtO
DojE4sRgMgpu3NlcSHQyrwVDdNq2rmDlY2KKrhygqjG6f2e1R/fVY7TPPQ+uPhDA
sCO6liGRC9IXJBKceg5mS7KGir9B+laF+em5W5Ucqf5Lgp2iUvFoMBzwcAm1OzwZ
su/rFpCQl4jsBEPip8lsHN7PmVoistRr+KoKT7+t5t22lFq7I5NA+LrhJqBpJ4RQ
kH1blIwEitnx4lKpaDOtAElrN1wQCos7upzW9pp1+KHKZ28LsItHIFOwZkQq774Q
BbGrBOVmRV4a50Q7/Nvg3hWMrLR0gUTawVgUZ44qkFoA/w8J/m/nHgI2zk7WSAlx
BXeR9R3NBWDV54qdf9cE75APgpXx7xadzrg0ZO1pZmrsM1OiAbQfVjcpvbpz8gPw
cReB0zq+CSp714B+g2jdBCAjMqo4CuL1K5X49+oMrGxH1TVAaPB9KXKoN8FELf7W
fq5JdsNyJMM4wNZrgaqRkFp7qsthjnt/TbQk8sYjjO7NaL2R/foZS8eLltj++ySr
PCvKReyTTlVTZuzhBGKErrZNcPZ1kclbR8846b/uCANhz0FIvCB42pO+6QUuYW51
upJrd4vZFJBNPUrhJQTwfPNBzw7yXgL6q+8jX0gb+BbiHenajQVnO0FHlKHX1jRF
xuG003v/ccNiC2DXB/fAgmrgvuT+SM1CwWjAqmf/FakikOzwYw8XwE6JFYhabu0D
e4Q4J3qlO303qHUj9HtwVtdaFfFOT6zjXyx7rxfdJCyzbprI2cF4Z2Wu4udgRbXo
mzlIh7VKUcTJc2YhJ6JxBv/0XD+a+ELnvu04q0sfPzccUTvuiAUjvm6AcTX5aN1T
26mUg0OfYQ7kjbloB8eURQka5WhfhzZopKo/JWYWev/FMSjaIYqlCFChC0QB4BkH
stZjid68WMMOK2I9ZkUlUBpl5A+Ct1XdvkdVm2xCluISa7+bFVJR2pCJn61Au5kg
DqcbkANlkF9FOj6WFBPxltDdh42ymiGqcZq8KMzOHmf0ZvPYPyaaAcpQlELaQxit
eIK/jffUo7F85EyIb0t4Lt67x6XqMKx3BTos0ceEAkKvHBcbunJ68CGws9s+iTIS
1RuQPq7kt7zHJfiSE5stZJ6AoL61xClEY2VFre0BITd2hV/F2iFzPe39hPWQqUTb
2qSI9V4J8fHAs559BjR5ZxA3Yejqa2x+YOiCovqORMLgvoURZLfW8sEZsVDDuE6M
zzrQSzji4L/THHbSkuEwbmgOEzr0lPLaLkPy2lDXb9aW9vIWL4WEiUaJBTmUZLT7
cWAoRc3woq4UC1C/0B6LczA0szNKmW/DoOeceryiUzeSxD6oAFS51KF0uJNKOSQv
XT+cqNODxaNkH9UDg3jdCSpUrESsz6HafgTHEIemrQsB4VS6ISLajes9GyJPE4Y1
4xZ2o/g7ylSh0AOMf8539ibVN2o1FHU2x7cs7kW7wK3PAscKGcH+/J8mwvnnfvcQ
73lMHoeJrByiuzmLNZj93mqnHnbePaDTyk8NtWu+7jtJ7me22GhZ1gsz6PPFvA9x
/MoiKSIhlcgyTsCUA4pSkHcw0r4bCJWnjWf2vo5f6q3VJAIvA1IHcXGlxzygSRwT
b9uldch77cG12OASBqCeDipIoUyiCQ8VpJDzqQKj9LI2ildXEC/kZjGFHZa23Y/i
lICfJt8mwdJTexHKKgO2o32h5pRcqw4Ht5QVIfkdtFKsVlSQCzgrgwO9QNVH+28h
5AdvIrZfrBQOZ9wwtpzYefnAKmeQvsi8iyh5C1mGqnMN6QD8Hhn9l/rUCk3cAiQ4
7AbUxw+73fD84q1kvC+rD4LLft7a1xgxb1m6aMyfv3zLxfb8PS6M2HAR3N28z3Rf
mdWr/g95P1HZ3ugyKqjproHsNqXM2MT2pcsHUav+c/Bn3KjdeaLFnD3n1K2ulhik
qMreowmOuRGWItpDu1I/xP2PK/80R98YzMek1so1+u6XXVCVoM5b/bfiLfUWs0vX
yV8ci/jYmxPIK7Y1Hpsduho6J4NhzEc7xsiJ/6KcySEtxYIKphjlXExZPVUWku9S
ZLcV3JJQAV4qY4Tfc/uXCDyR4qn9vCp6wPzcpWA+QWfwVps40qlEw2nnhqLEz7vI
OwJgFGtppOrM2WFIxmo4Y5PJOHPcNxCkyHTrWRALDMV2emfwf+7iognO17LzdzFH
Bq5u9EAUEnA7UX8znGR5FqqfudCMBb/n3L2F+sVZem16x9kyC+n4iF6EItD4D0/p
0U4/OCUc61lUm4JVF/7pP0fAlp+5aunJUCkPztIp47C/RJCPJ0eEEOjHsGC24cEA
LTASSFRvNkAZByu9PNeH4SakH9t9BO4/uUBnCXrPTolEWKoYald2Dal93Ap96snA
WGd1UicCnkC0WVMCla7XrZxseMsSoZCbdzC2lyR5MqJX99HyeaXYLzvk3Yy6YHac
iMuIIOXtl7XOTIgW+M8bMdgn9s/qmWSY1FefOkii9DCGf5G2Ar8kIrKhLgvWsPIe
9wAj73o27cZBBHdGx5+uVsFWVWd80Ido5Bhqp6SeO3RNS3HAEDLZhnvA9H9h0RbQ
Xswyt5ei+S6vdrVeLDpI2XLwNexetUrwjnx6Hdm8w6irQMRLV9c9q5G7E+P6YcQ+
xfIN+01F0XLvwY7wRQRaGPb02aQV5nIg5DokjhtAMNGK3YUKcwb7a53gXEJeC6CH
tzYBtJ7Vbkrg4PqAlVT9toe6VEHDYWoQmNnm5TG2pfMIq8SaikF9aY6HJXzyB4vx
egzdoWi/sgpfp7ZsLksCRQ5bhL3LCEaqQL7kHCaFCmbjq+eKMOp1urwSreBPBJ/X
Y4UMw1G9y+RRDXpsmiZunyq+Ibk7BBl+il6NnIH3ovFVtqO3/aS8vDH132UD/Hc5
mG2An5XVRSmEJTfNzBWgZRWn3wRJ4sFEFqt3H3XyffQjARzTLI+rtSxFsfd3rZPc
hyMFl9sdEe8XWsF5UybULYCLtGfwsTttoxexaaDPtJuA1Rdp/bWBJbfmge14GYp1
5XLtv1vVklGf2S3kw1JUDVzq4+OG8IoH9t8rGkcktlXNLKwk6If+Xns0S3n6rpBv
fCJAR1KzPHXLKO2DkT9jSS5371pkfNdjpJ1q5knm35i/7SL3q7X+TA2R61ca0Eiu
uG/juJzHBtR9fU6Qy7vzz3mgvKBYY57uluAO7WPIdrDj39awoGoHE3T6TnU9pF5V
w6zCJtNUInWGhxT0PLYBBD+jxBUjBa0OFR3iITuH+VudV3k61/D8huRDMpEFU0Mu
04XqJvUP9hCoD/Si2rM+2732G1yr9V0G9Voe2TgltXUA+547OW87K6Noopf/Ig9Q
S6GL9ZKHCA+xEBjEKXK0X7uJvVJEqJM6ho5xM+7CprKu9AqaxNO9gAO5k7x8SA/u
Yh5lxkpL93PJ9yFdQmFtZvvvM1xdBPZsfrAQbpXGjGUAR14R5jN1eAAX2oYJmX15
HN3VbPCZwK3FIFVGHAnrwtIid+rxx6/KWjxCIPS5CpafULup/z7DiF2a29EXJue/
TemhvOB1QJoWc8cN+wjEmvq9dPEYzp9HMSojtMiumzjtyXmqP702kRSas72LWM3C
SkP/erLVCc+pEIe2a/a6vgz1VZ+4eg5W7CjTUUZ/Tbp6izLK68faw5gqHG0W0+6u
2MZk9nwFmyI5F/TmT5/9S6HhCpQcUMLokFY3rLcB4kh7szdwlixM1VOXhQ8+/vJR
jcyXGyZjbs9Scl0objotRJy2hg9RnEo/c9CRVj19cI/CEQQl9Fmg/48yRSEeH4xQ
lejzHbC2P/yujPXyuRkifYdLUR7Sh/Bcf6kopfvukfogi3Jg9EhD0HInxtm88mFg
YjGXoWQokMvAo53ugau4/Q5CqIDDQ0x0MPPMsDI8a6ud4ECmk4ozSZpRgGyu0hJP
fmz60vHMCAVrk0TY+6Tv/CwGqFt8R29ub8PkBCZmPy/Y9ZH4DhH1MvrodLHHcI2S
kkMZHIwzgElXe3QiJOFEGBwJ94yyxzDhCMcDUV09EoBpdLDh7mrNVkdaYZyhq8Uf
t1C5F+untvtzCHiH8G8jesMGdETmFlfDnLafBQnaJbB0HKzhvw5Oiq08YAldM6hr
HiLzpfEtlPFC1NdcjrE8ODovQ4JPAHSBHuNoe69G3oi1cjDXtLcPL+L1tWm7tPiP
OyydEsuneMarWu5eXeC1YKh4BZ8P/UHje2LHlV77i28B4F/Y5QJVSorQooOSuvJ8
9VPv8Tlur8HVTuBZYke57N+bgVl+TfcEdj6/QKDV/N6BYi8pIuA/KmNdDZj7e/MY
A2T2f8eo2C4Eg71iV7qz8ElCQhWGTardtsYDWlfEz96pF8S2XNdVkBsQw3rKXPd8
PPTO6lE1adIFQKpZuylfzxX50KbHE2nyEfkTrBMfpx5Su4PCPnYeuklR+ZLuWWgd
NhsiDNZBAhKB5E+fBBWeAcGgDeAQ7PhwafemUzcUVqhIz83+qQkaj+PQKAzZdzjG
DKFmJ2YtPmatR2etqJLs88F3e4xZ0lGyE6FAVZRzFRIKEQgOIIfIhBuoXBVgYZjI
S1mVkeHR4Zcqtp+VJJSfiKuqhA+QqQOAssOM/p5Bh6wH+fyMVPbAq16YPjEjJOlr
TJhpDxt9wf8tILkhJs+EDkS1nrDWRSPu8Put/bOKOB9LlYsG/wv/bIH19pdp6rdj
ViKNwrfYDMqEWW/mcMl9yEbrxKdOPAdfKXQANIlsGwuYIM5kSog4i1wH4e3RylSW
/nePqeoeriQzbmilvYvP2EwZ/KXFjvmLYT1WXi/jdfuxMbA2DFTdNFPxaS2wcUOZ
Deb8rqWxg9dUTQq3EFKfTb/jXJ2uzciA8bcwwUAtJEibZnDvyFSDY7D529ajJXMl
fkq1yvBqrUkiY+UqRbwj/Pnjzi7fWftFGpymJMGcMH67C1vOpsMY8im+vTXAph0y
z1Ljilb7QoMXiM8qrjpjOWKhHFF0eNN1NHVuAVbjdlnxPBvOXPHO66onz4dHlh2j
T2Z++jeXGik4paZm02UM3MUPns4iBTz/LsnzGFazJaCsgb1S8n4Y8IYzMDqVtI0P
/7oF6Wc/4njQ8ZvayJnEAKgqqlPQ122hxKC/TMR7Qd/2H6R2YVdwagKaIGsZCPgf
Putq7xGQfjTTcNs+cJ/JX1SGp6dPC84m9x2I+bjh523KlDPzSBfF81VZjhY2ulFw
ycgQs9p2qHaTVlYtgT4JDgFRUZflkdJ7Nr8sCMjnrOG51KzC7kQ1mIhKxxcqmnlp
bSIvId4YniARoGD6LwP4g9argfUNljRKP9JNALwWPEcBfFSE7ZDszgIiq6N7SxpM
vstcAkN/7EQmehsfgf2lKAvcnmi06DnNQXUQoenUDYNBqsLXwYl4jxte+AGoW2NA
1a4N+ODUjr5sUzP0tCWB8PRbfMvTuSUSLLLAcUmtTzq9NY2rb7YB9MxFwKWeU2Ig
vUrFC/sxbbjeoZRCuQ7NNWxURoNeltf4qJJY/zzAaenxISUswtBLEep8TcpENGyB
us6RrDyZU5qOVvy4TccuxE6HZ5/S+yY86EqvpfbDhBBA1FY1LoiMdcy2tgrLWm4k
DYatbPZvNTYE5744azyAvCQgyUPhEpW/f4LshVuMWpszaO2p/igRbLskKedGKSkd
s4LK6guVv9jEPnp2fUAsK1TxdPg68H7qVAVGR+SORT7PUbAlCYcOqtoVGytIL4Co
fzpH1+IqLZmFwxe4nCp/FGOS/4N8pROc9BrMm1woPI72KZae/G4JOqNfNLNNkr+B
/TGIL2nwu6ec+pKjo2M/+ddSeCgkQiEI+Z+wZXBeET7XrqkvmK/fn6CFwzDYoio7
h/Ek00tmwLNGDbCyz4QKUcVIAeplrkNYq44LaKauWyGCrzdKPb8ac0LOV/fF52i+
diC/owenuTQzqRyBsZEo7WmQ1eVosPVWzJrnXW93pKJQuUBH1G7yD/R9yTkUJIvF
XbQe+jRMSoYENwj6jYiVrLj4+GEDdcEk83Druk36DeT9+Y88inMmy7jP1j/KbvQj
V9zDjc0F4Tn/I6ZlXeyz5lxCaezWancpxSbY2o4w6D6vmb21hRsPB2M0ePQM3avy
ldc6YLrvb/vlwjZUANuIEKckOeCwKWcfms79XNvQO5VPzXYKAVKFoPRp1WGrZmod
JCgNtPta84O95gZ4kiA0YQbBKJbEZz/Fktac2wDIyzhJV4OJPq6VVu4Y+bfvviGz
Gm18E/o4fm7JJLcQ6HtJZ2TmORuZCToBBGPlpP/H5mSi+0qcXepvlJUlnQQsU1bn
igZWV771BiGUBz8hAxSudkoZa7eIA6MWFesYdVlVheoIU+8aYCx/P+i849ls/pmw
RNSBFuAV126EVonHDfNBKjWELdUrwq1DYX7Y7EKlwK6qeLVvfeRxnoAQyqfwgCYF
xmIUNF02FG0TT7twubsj+dTIAfSMefsunBq396ddR8jX+jn3oh49+GF6qNYnKZAb
HU6Gdixi66REjiXwlhjYejBtSB5cYLGH4cu9AA8jVWkltd0P2QOB4Bd9Gq3Uk7Va
IDdKmX4zEZUl4MU4dmGfo7sVlglFk3d3eaPSXGExdU8bXdVq5VjvmK3TtNTPxmup
c5hmwQMp84EjwzlUjHjMMMa4mEdxnTyyTW7XoW55OiwO61J8A1StZMOWb4DNrFhY
t/AJkxUYDIF/RZrDeSwIDA5UnnrzpDZCcxbzYAr3WKVzEYq1Ym9eFl3xPsL2pOwS
yyIhbUXEfHEIvjyBU63uoEGF3wKoftey+hO4gbaHMxa5f3A+5UVJwMYs66VN5YTE
AmNuCX/yIFWSuY7Dx87ZmS9opCMUrGKpVowGAm2sccmIPI7Q8rfZEEUnJNWP6j8b
tzOmJ0b1f9nMXuJ0PrTw/kr6FMyHz0z7TEgtOtG9TqxMCV3paoWnCgs1sGy/n1x9
6s4FLCOQA2+OvayugR5JIu6gWVKrcwc9nF6AlyfOGjJlcyTN8roEjWK4NbitQoiQ
yVYB3k8Y0bE5y5BarwMM5z4GSBnMhGEQguGdbuz22Ou/+P8PvaFaJJinfh4CC4ko
wCnIcEWQ1YCinyVy+0EZrt8gZR2PhKveho4jf/qSAzqbqGGjzDY0KOexSIrdVy57
vL2am4x0m/phxIiNlu7h1AhNg9x5XvlXdcpOSGs3vM5za22uEpbwaFNnEtZzyoY8
28hMJ+cWA4l1AmTOBbkSwGfNJtb3KyvGsxdxIIgNWfESF1nQD9KAqKNC8vW66sOC
LgUnRiIPdDqN/8T4uA3Y4lpee2te7vnVQw9Dth8rrFtaADApJZqBOYnVtgHZozFJ
CdZYQeppnkuvNN3jCf7Dwy+90rpy0KqoNfjI8h4gBK+YjG0QuC9WlA37WFiATpfx
9TK0OTTUCpWnygLJF4VlKK/airZ4GuMK/ygk9p7gftaJFmzIM+ec43upA+P3xA7f
g30kX6wjrLXOBtTXv6RDbF4tiHaW50yz7BulTTMcJ4AOxzqV5tyUxK4Hf+YJXZNA
67zJw5vbkehvZVoTLCJiIY8jzGVYHKVtgVWUq6F9ZzJHEpXbQ68S2zbMQmJBQwpp
Iy0znUs4KEdMGx+uRXrM9qgTShRzzhTEIylgqqQS8GWTDMf/ERA2vDE429AlUzwr
H7Vw2vs5TaHRCOV04cAQV2ZR7JA4mCvamMCs5wBsmprj6J1Hj+3xIW9MLke6V9ZJ
87Q68qNx5Cs0ChYtOyxOC7RYYaWTE04GjBPMjGarabsYSzj11MM4yT/M22vpiSje
8PLb4th1TDI8+T2HlMPNyOe+MJ95cHIzWs06zTUy1gTxg6s5zt6AAbsonGYjvtxx
DPvLkSVBlN8HvYk8kCS1XSWcw12HpzK1xpRu0ZCWK1jwyOx0RH8JTo4/LEYQW4ez
kimsK+giVeH6u/LAGScoR0Tnv4ISD5uIY/Aew8fZZfhxlNrMhQc6+zpxGX78eALE
CeTaqt3LLeuzF7G0S8PyqHS5UD7kmVGXpH6CTL3QUKiawiIUmw6mc/tZ1+hI+kHv
7mT46G29DPBYXMZwcablC1D9L+00RsRU3YVs+Ej4QMdKDVUi06aUSe4taMe5oO6J
W8YvAnPpfj5izz8T5BR6knPSMIHZc0n3aKD+6ErcmNdF/3e54Q18ft6iVTDyeaZP
RZs0nRjijwjuDLQUJetqwp06GZ5l9qlpUr9bdfRLQWVnaXzW7r4s6e+makcQYjoL
iYgsbQ+ITOs0i6dLqWTi/Dsi/RduRQyiMP/tOAMj5SOZtWJvsQu6UVL2MtOpDVl5
RRpH7i8tRetHJAejEB3pzRBaujw+/SxAdFOA1+4yiT2Dw9eC55lk8/8Amh2E8u+c
+ZeqRcimbtophFwU/NxFU00IFhQp/kRzI+Jd+pfCIZHZwtNwN09KoeUJqO8n5Q0c
Ky/IRfg6iO/WTgdDJP8eEzITRvUydytnIzqQF0m/lGXhJlvSrU0ilbiM7rPysSzi
/WeCHlonRKfrZwDIndUJyMovS2ojhTPt78WK4iMiUZsaDPuhScZXNCuHf9vIzPFM
vEJUBU4g+ooq4KGLqTELPCPOxs0PyrXVvAzYEL1y9ILzqohXP2x0hozdxzBK52yl
kI+sxwojffwxgjlPDaHTtvnvCKpWA1w8nOspoqqZqwpyrtGLhaDCu3Lf4E/ov5j4
q0bpdfDJKXK5+scu8RWvWVy04VWI1zdQrumw33ANCiXijCUOLxq1DwKVrg3Z7u85
ORGcV3ErhjZLc2TqsNqcyFj+xNKaYLyHQiD6DaBqkiQyRdn7l5ja2K43E5JujTO1
8DA8cT1Vj234gZkee7tfPENFSN0QlMxwSThAZN4bj2o8dqER2ugq/P3MNXNoMtiV
Tq4pijl3bH52RHJOHAJVya4n1FMpOExwK8AKE96aTb3dXE7YCdv2PQRhwLv4HySZ
NqDgk2tz8K0nn5rIqgdQD95No4qFkxKXVr9kKDB3+yi1uYNJz0YcFsJ4E/vafREK
7JOZ/n+9cg3n0P63MPmMSNeNwwU/pf08GC70luXevy3IX6ls6bQcjlbdJWNvig+z
O/4+LgqOFshxfQDIEtij7baWhZuqUJyK2lhXewg/RKQ+V0JJeLFwxS7f/epUXk7Q
X9iHjL5WsoGp2kCuNKxzo8yvXxiFSDG8amRiUzFXZoQASk2pEgxD2l4JTMLgctl7
OM5CNslnN0Ok/UapOEubPD7240MVq/GU95EnIpzIw/Y+sbzdG0uFNLsEjJI5dAhT
e7eZVvRa8ZvIqv6IKVIEj0/SHbHQirC7HmLUImX4kU0c/MDtygWldzBYPU7FrLu4
wV1xTYFPmbZoydTiYD78JbAfPtqhdeAmhXyBg1sSIRUqkea4hTqoznq9DTgSQSwI
8bdLRdAiLORCj8tSfs38epFZha8a1pKMGPFa/gZ0hh+nId5tks8QqqXFcQil8Tff
16gFg0DJRJavnFJn5nbYgzXmHTsmNobQqsvnDySemyYHaidOWGSQq9X6tKb+stDm
Z+vGDfQcngNjkXkHslJyR4H26p54fYnmfL0dzCbk0zscdEgJT9NL9G3+RdFcpazS
Vhy9DTMYIyQu4aX3inyxONsy0KW5kh5vyxfbMs5lMXl+15LOOgTySnYIyhRqVkmC
Lyb3MUxfNLQD+ruCuOYyEW8ZtPMS1J+Bw/3m9JbzvnqC6+u+OqI7ceLnSoDUrzC6
K0gS/bsK8KyonfLqosBKKHSh3CxLQ2NW7U5cikb/CVec+omV9UcMxhgAhKQEryHB
cJQZ9EtMWA1936DOHhc4WRSclWGxqPgWy2tWJSgfPBbLj8QjGSeUu/UKED/nNmaW
NHdVmpJxoegJ35k47AwWvwddYZxikr2nx03KnND2CawYDcjbQRh4k5u/072ntwG1
Zam2soB9xzA637Mz/wjZrW+fxSMQosmdUT0MRE2d7uNnj4kZh9ZT3iTLYIF+2BY2
XUUtIaPte84Q+7fZu6TbCEGFJeTRF+tZZ6L4mebsLoMo2bn5zlpYlRjSjrlKAd6k
v+o6ch/GwnigxuUBDepEkRbrWJ4T7aEddMsMmHIxoeiulMY5FUvWgYyO9mKeRawd
4F99Q44CMDtFyOJ7dCOlM6Ztzis5CjCc8w0nxrfEqOYAINUDWMg4K+kwnm8oJETW
mo1amgskV1wBcohzBC/yH0iFQyrtelALgZE/0xC5KMO2lfgxTMPOZ/shQcgY6ui1
y0+k51COnYz7AZrmrLx4iMM8FK1nK6epyWdH/dtOwpBNswnuLxmO8R0LzbBTEveV
Udgl5Pnoy8eqfzoVbe4WptHuEk5gB5ZeBRgmo1rmCJ/8fipkAV9fBK3OLUJLXj3m
aKUXrvfAO4AUL2oX+X1NPsjZ77g+aLErtcJXZR6csFX9Zd7D3IT3cz6uiG8Yd805
b/uRUs78pmRoAjvAaSrr99i6Iy6KfDx8ZNpzDLZimt/L8ZnBG5VA8bVnOm96wtmk
6uIaZlTnhPIWcUyDwvKfTQBCLn4WIF/ClLtrmH4RErq68xGyz45RX6GxmAcQxLbP
u9Xz9nE4oKKoWP0x1BgziHunITiMkdreBFx/5k+QSAAzmh5GhOcja/GNs7EIAbL2
B1/0i5e6UIySDPp1hTscKlILOe4Qsrkw7DncKEL3VV/U67G6Kxy7cr9GLYQT6JDr
i7jMtyQhVGa4+Ug9fSpYdDLnzrKjDybvj2IKnqVbFxGRUph99ZSRgefP8k/lU4Tg
iAaRtXn1rE+jEFLmnxX4GtyOV616MtKyteHeTMTtm8ZsuK1Vyh8gWR02bNoCzpGl
0G3s96sbr9+rSHRqwqMXfOc+/YPWLX+EirPQgWnFcF/RuMNIs9kOd5pKZPZ+V10N
2zYauhQz8dBynIbkO+vAzBxbeGeKlrAkX8u9onC4yM7oTIPUSB1ExuW5edmeTk1M
yoGt8pPTxAPkHfEyEkZZmOe98lPIkl42KHblRsnIDxYPyRQWbJSJBlRYrxp4oxK6
dDRpqkmp7+uWBvzkPGYdp/pUxcQ86QZPMqdBVzIotMVUiPsW5niWDdxVSU/EfpAX
HfbiRT5rk+kyNMRuKUV1YI/MZ/a4RcctFJ7vC6PjRCC4hkZKDayPakmMCoLGJxFa
VHhpWLyEChJ5/9Jxcu2pahU1hdaq1KlLjctN+w18C/P+LjVZ0mgCovxbhFJSEFLd
sWAB9KQT+zymidwQHqSjJLzF0fLDCrKkLGC5VMVjoMf+fV3dMYiwt6GqOj/0XM/2
GqHzmJbFTIXlh5DtQeI348EugHUueyyeAvI7/0hXmHVDwCyc4K7bCFzKRkAWLZjC
mUvavdyOu3ncd1BGOWkap+ymKh9EoV6gNVD/Aa9EZJbxEMSXpXv+RQg3fnotNuNw
65wBkV8TjennIZ0Uvde8o7uo8kCdKN2/j/Op5aWGzFH17Zta2f+4RlDrIDk4LzO6
MsxnH5daP0cVMoO0gLDY7Y6cDl84e8mqty1BZyWaxWYp5NaOoD7okzrb1ctuzxMk
6M1uDZibX76gtkLDjOcNiJ5CJBxKc2dpXK9vrM4ZX8WRKOwDBvaRtipQkwTuNbZO
hca1hfbFNPpth3ldbEJeBp/T/LYwR+IRrJ8jggiVQ6n4NB89hZvgLgcEECtLgy3i
15I/rNyGUtH4kAoTaim/gWdwc8GBjVbaVcHjafIeTBz9pxi1iZxU/G2YmVAVHMlI
LhN0eQ32kv2zlnPHXiomBAKysNMce18FkIET+5lgFPCGocSg9bVjx2x2Vn/wp1r8
8nLZu3Fyg1ENpdD/d4qynInblCPoyP1ec/lEn4efpn/ZOJKfNt2de9sulZI6EQ2T
6Lqv2McgYcyNMfCnf8EFDbxfZJtvSQAhHJlGjIx7ULYOEw7mTguJamYXJhQ98yrh
fvb9cjPW70wzOYCGgHWBAENQVbQe29iYnDkwMA8ToBiCmUhaNgXAaz1OyU5VNadK
xZI5a6cLNujSDFVCDxiugp7izDBjXG9/6uBJIMz87PbYgodhuqnUxqM1qq3s/1Bk
nameU4hCvIs5dBWzyMZb9xeOmEGh4+585qERXTLIp3p++rrUmyt/rjnXBZWVK21I
zmx9LG//15s0JfS80MPQrbj9jYILT2iDRYZHX1YDAJATHmME0BhCyypkJuE1vC8l
Nh/X82QLRh5iHQMrMqN76lPfzSy0YppZZJaDPbLJR8Oav86Ee8FFT1Y7H2bRrPop
p12HpQLXGZCsFiG9v1Kd031JgABZbeSQVYLzzF8vzSgkmcZemVfY1xXeyxQ7VJDs
wTN476twLsgj1F34foDBThx5+TpObEAH86G0XIi+vL38dd8q1l+tBHtX0iS3l6An
tsUhMzO8XuJMtkUaSnpo7doW2bNSR5uxNe82uKkJQ+5HtNFCLKFnE8JtNNu1LcFi
g4QH1YcdRkBkDPwC+G1i5V2RonN2olyRrByiEgTtctaC/Vgvv7x1pF+ZQNWY5eKC
OgoP7d98anQ09dQYoVFeu8BNqjsDdVnSvNZPqx360wTND8o0BnL+5W4GgdcaBJFN
1BTReXkuz4bLlFa5GWGjoxHnlfWo5aoEzOdyFGf9MRTyg/j0+AgsA5szHfOyY4n/
eLqtURKucvOwIRLLHlc8Co1a1xEFnyjgdMSugkMuQBzR+GH0kqtAZRyRa+mOXXqi
q6M7Uu1HszBrFIzop9FTtqqj+b8cbIdP7Sxox692ku6TZnInLyCMiAdxsW4faSwz
JtrXZcoXE4fj0NeABDMGHAeLksMYIfNKEGoUFNbJ6HULuADlRL85AKsrO8Tjm8kX
x/8RZkkuKysEVJ7BOkW9++kn9mt9fXI5fsrbh6cNp+z3ffU1sF7/VVOrqAXKHxM1
76+z8JKCneuPj9HizVOntGgqXiz6zJt5MsPz4DnGlSs3KyB4RnwnWnlxKijxm2Bs
pm2w7p7eUVzcNey10zK6pZsQGnx1jdQs1cVECPcZdjtprqft716o8UVjtuzPi/0G
YzdPjnm0ESknw8vTHIWsTg7T7z1M7kTxI/OT3NXzETuu9CSh1isJ+xJ1k2BbvjV+
XvZLyshcbgBaNMNbIMqXQOXqzhcKKZZ9fA0BuE0FXkwtJf5yDdMnN4TGVouf8Hs/
flyNfIZyoFAQweLJeE+lbbLoI4s8ZrxwYSE1Mq9h9b6zQ+JqCM+Y2DljcIhX9r9C
Z5fqhVqQnGY7BMZ8+LUFb9n+aXS91vspYB71tQGwaeT+q3RXT4CxYJWTAfhRhNKC
4LEa1hY1A+cWYGW0rpAyx0dhFmVXYwNauTS8zwM+/EmNMXSC7IqpOqWhr9jkH5uq
Totb6pem+A9wdNntBNY7C8JMk6DDr2oLQ3qXP8Az5N18MF/+eR2jG6V9BDog4cw2
Z12AXHtbmg84G21S0uHaHT36BuH7jB1l+ugQagPw+O3poHTEk74i22KEXCWXNY2x
kaeAea7bYFmluWci+CiZTUdEJsYMLK8yl7ICkQaN5HIgjCtvHIlIl3QXqdOXqgA4
7MMzhBgofvrQICVPJfWoGgIAH91ZOx1m1seUya1EnlG/LEU7hamAiz3RdvScePBR
HEor82xIAXeTn3N/dpu6CdKRhC7cZLN0p0P7ABhkO6i8B58aqoWVnFrZCDC+TaQU
0kkOFhruzTvQfvEzyoRSucoCbw9RgKI32Jfci6Bb8P5KsorzAeuybPj0IWktoZ2w
H8uD2mMh3YQTd3TUjGs/4TrW5q8F092OnW32lI6vMKAocy9oEBlbRsmL5TUY6wb7
1a5Z4b1xUXWXCR955R+s90NPvSvyHWY8eq7mq4nZ/N6KclkAy5lUVQYaZzQhxCaN
eYbXUvFVVKDf4pRmpjUaskVA5CiO3w4ViSP00hjBsL64OHqafNvouwPnA/grB3da
5ao4l8dGaJJIwXO8sBeJYMIQTJg/gAfqZszGP5WmLOUspA99eE0bx80gb5jxtA4o
MgUpJuLcxwOKRqxpqWkym/A6fS8TVDXbgbe6Uq/kEjwALyM7wXc8UWt3F3vREMoh
+aUooP0kzTL4+MpD7vVDqRcPM+3EI3V4zFMlSmP1gA0IuwlgXRuVSdh35AXJHq/U
kmIxDpQcAHm+MqYow5p06N0XfWJtpXJDxhLOS8Oc/57PoFG2bfejmw0BoX7ZaRTh
fdCaNl8sz3QKp5nr66A0U//j0qYcJYpIq7lo3l/ZTQH12CwOkgUNrqus00z2oxyf
t6zQTOhb58mf/DqM18hRe2Lr4f/baw+ykG3y6iweMqc33TyTVZtPixusAD2ZVOYr
AsRadOoknfFCAgcPveRTyaWU58rddSulJ3aHm//bmNfjJ0OSykaYdMMyrXb2cuPB
T66SifRB1ACzVST0Koaq/DdwUdp5CJNADumnxdrh9L++ARMp+yr924LZxAZI+nqb
lkHbv3yTA/mm5RILHQnfY7GSaqwLW28VrDRzW7Z+ESwLzjkXD2bbqau7ASEZEbt6
pD+G9rmdZeiib+VbYw4BBrU6t5yo53kdKUSKELZjWa39fYwddvJ+m9AqLhry4oXP
5fVfzoPuHkl0IgI4yiq1sZfMcY3DvXfvJC7TkSMcH4DCuDurFAqplcCLA466zEd/
sbfLCtvbORO1mHJn+XgKsKQc7VcFXre7l5kCIlFr30YLu0tmxk5LmABa8wcW51vU
o0wVse/Av93k1vDcb02y8Bhvzf3QSbcEmZZEWjZblSLrP9N87UYpFyPM9CtaNWMe
hGerm3dhDOujahNYjl8wdWlzd9+nnIVREHjcwFIpbAn9UhwQIspCvS+FCMGH7M8c
qV1hK3tIJrfE+uRISKrHJx3xYhSb3i2XfGBs3bIUYIDN/8ONskOQ+4fiIgQZp7j7
O113oJdMEetEyN10eQRDc14pTyzRtHXlUeJ0UeKLcRYBnAR8Oxd4EOcBVPyZghRQ
j9fLX42zeDbTEhUPxaC4MORxKeH+B4xyw/Dbdqbb7V2POPD6U31KiIV2e6osfeRU
VcpHyDZbqEKkgeJ813DtSMF2484VR3fAsKOVzt+hYdi1dIyJ06QpAhXoQP/S/T7R
pPc2VBcTj1vgY06e/tDKdlyj5xtok9MYbq4oI7BzsFtLRs5Pw8YbSOTQYb91ipMD
p+H8LV62NEF5GualtBEO8tjvRZJ0Kcfc2HHrRDJTMVFAUekZGMvfkeKeD9XegY0i
Hz7nM+1H/Twf+OFDkMsURNu/V3pClPm7iUOubaWBEjC9on+2oS0Yro7yHHt9a9+g
b63AVFD96Kr+IbU4DuMUx+FGOfnLsx9uCU8bGigVtRk/1ziXW/yBsZDs/zhHch6+
WLl3q3AnKLR8U+3tyKTYkbKasvYamSpKBcVabBIF4+ztfaidb53bB8zaXnzgJ8hN
UTsMwVN09bicuS2AT7vejqridDaQ4KKhQYJw9LUbLlIdeBgCM6Jk2Hq/XcwaVtDP
/lseD9w8DPlkrRCiPY0+JvTuB6Ayhb0v22atR2SdSIfJC0dTBpZsX6LOdz1AThDN
iPmuzFLYRbwD+rUngdEnv6Zsivt31tfGVgI7f8YCpiP68TCgBOBLNOjbYkXeKhTM
EjEUfwjuq4mfSO4kv7VMWz3eh+TY84YDgZiISrARzD2OTxFKUOL4XHnw4dRXqSSM
F2ygtA3u0lKEMw6yCkjIonbazigqykNxme4yXMAmvGPISjf1ZWe045K9iSUlR3BC
HNmbCwVghcoNRTKocX3voElNxxNdaF41lSBlOZL64LQjc0cmM7iRQaL054P9ks2F
+CXA7Yq2296bVH2FQmVcJGJXuW0YCodM3IP9QyNaOtasQTiFV/aPbSFvKnbNoTJ2
ZPAkCQKDnnv6NR/Ie7CT1SDeNlB/czrRypaJExCBciGr2LaQ9P+0wIZO2nCiAAoL
e5OMpkigvJs04+L8ux0HCThpTWi/6Fn/SbSR7e4iudJfgmgcMBhcjRQzAk+B1CIC
zoOXbfX8MaHZC8BF6kTtFNxZs1iTrBK0ViKbe/JzhrgndsEDMGXPtKuS0x8gsRZ8
nYUa+VZJm/s8rltKaSYA+xD3/Rt2UNy1xT2UdEtG7aK3B143wI82K6J2EA+pFmIo
/OMQjRZFfocpl5xngEhRSkGkiz/xYjw9rphYMfkmnMGkxWbrROPKz8G+OhAcrtEI
9GbC16XSv/pmGGZI8zsqr0crfowuFSdZBIhIEfFhSFFXgiZwK7rUzJ7n2Auk+AKq
TV5XAWFmCI1T5gaENCvFNXfVD6ibQyuuhq8PfU1bPxA7lziL795ThiDSQXqf4k+b
uUM3iuW/DZRBa3uCuvf6U5Nhuof70XYl4UdOBUVMdIzfAafiLAQoorfs8ep2U/YY
Q/WrydEXcoB305BrAlOetGZ+Qki8QYBOCwqgzK9Zztf8iKuz1rL7KcBp0rZSad6E
Ekw7Qi+PjlZs4TfZK/RLGOfJnxF3/e5LNVIXDsMfP3ooSkoyrQBE/KHRPnXRlQtZ
HDUctFVvHLyZvqCHh/Hd4AiSjJb1L8D3HNMdv5/q99Bxltmxb5PRDPHnRxXM4h1m
0TVaKF4mUYTIHJg0pbPwB3gzL9hgVFCyA1yQCHyCO3hYRIjlSoi6zNi0P9q0kr13
z+SMldTnLOdSVBM1UGIwRr+EHKPNZmVX9pjbIAuLwbYxatFmbGQM8op9R+9iwJAB
zB8ifF9aZuhEd8zNbA+/Oy6bCSPPPRnxC07Y9AQeIxps9qqs/RdlAMbAdj2uoCOr
4xzc9IAx96WL1F8uJYCzfon5cTIw738lOSqXh7HFPNb6+HlNME1O8qF3VHlQYmtK
b8MXcMeyExr2KumLS7GF3n9qgun3tmEbsHSL/Tl5qCOcfFYfLQc6nTbXcwBXxWFG
vyCkmtF88kVidq5+Tvc9LKf17Gt3Lxu709UVwMULlLZo0Yb/1iEpDjBZ3n7d2uJ7
8UG6JLPI7wedAa2b5mdg1Ssm1YOQRH7MM9QGvthuNxqkYIE7YNibngMsqEA6w2mE
800MZ1mTTZMFSimpkg1Mb080IxJd5AXdJEhIClOmOxgQvKo/PyHVxP/pjXCu1mOS
s/3IOe9YYepTqeDOnH8HXd9IpOL1mJ2LeL5Ivo+gb8U9p2ag4WPk3nqIK20/+CiJ
hyoy++uC5DAIL0eIVTujwu1CY+9ygUjcvGeLB7WsHTJDdaH/RJUIPAynmcZVM9bu
boPHhXU5b0D9DME37nDXzS4sr6wP64onXNYMlCOFAruVH0ce1q3sKd85lA6ioJhW
5G+XtGspvmoJKtt5LU2RjdlVBcQaC8CrfzgjaqyqXK51P15A4b97K4M7ep/T+73L
FB40oAakT0ncF1JwkUFRzBBt6xhO8d1Hy35RCyCd7xcgcdeM7jZsD5vlfYYoEqZF
KfsrMwcQ9fje1UZ5IB4+whVo+Vl5olmpi1hGf27gxnXC8Yy0f1+TcqvkUv4hC2nK
X3zLdrdeIvzFrxRvKTCb6Y11c5UOx9IdgbQjvQXeJFFDokO/9Kc8+Cr1atyWabuv
zWfaGvaZXvXY1l0I3HlF7CI1zVokRThWjWfe4t+m9oYSDNo87kcW1XCHgLmpLLCl
jHMMLtvPd5of/aIUQQ5v3orkMcb0eas4pHED6QABt9VODJKPRrkDIFXthyiMyyL7
uBIzgcd1v9zKB0sYT4dkwSTDMjzoWZfou1MsDB1rlnzlWtLCsIRES3fcxPZMAm75
rH8+PYPczXzeIhYEyBWB+XsDosFjspM3kYBRSAqyt/DDw2hslniWEpO/BsvXloJR
mHQu6tCtxUT1r+FumffEez6fShiTLdw5E1Z5TVRsckLUNU4PhmbcXCvX1e0wk3wu
A1c9GA8L4FDNQACYWkxbBnxVE1yvIP8Twr+m5juQGZqkvnv+C0H/Cjnf1mOwT9EG
I13s+FzpdwAE2Yv8f9dmdLY259rklnbjY15aUMmocSO+hEq0U0Rvt4tjeVzEkghV
ThocHloifSQuY3V00COGC2gJ9gnmJG9kKsUDeY2Pjah4l89FqIiZ2jFf8SSZpC0P
jBCPziel2IjA1TrxH7B/HQhe0JkyqyJXVgFhnnHE6PJ52jnBWhfMENxPass4204Y
6WamVaY5crYTtJ8V9H79wPFdA2nI0SJii7hCZO+QIMs4z1kI3do7c0seZigJv8FS
PvLJ/qCrwQXGyxRbgNNJZaK7C1mFwNcujPhlsejWDEfmcQEbnoSPBvNJJZKOXy4h
tLhe4jbVypfR5gUB/5cTAsqbNfdqFgw7JZMZs089XHy5WhtETTRIr1vkxkEuYecc
ge+pkoNHMJZmlM2KTbxaQvyBoHqHkga4iECB4ku4YwX9QcC6PNIGXi1KUh5BqxO4
iTlosoluEqFIahfF9tXDDMubF0Gq8OqnW0Sq4aHK5JnE4/WRTauXneLGV3f9LwAn
KrhIDPrwDeePqSPn28m7zddpiUhgs+5UnIP1QN1O0ilfixR/PvX5MwBYLwFgE+5G
wOed7iMb/vTTx2qEcIqts9Lwy3PTmpCAdZNVJkKiY4eaf8his4Bchtyla147vd9H
Ciddv00nT/ybcmK+W8L0BxFqkF7/bclCn4fePrM0gCrkyrL3fCwUe2TPXjdZPRfF
BNY9qxw76mE21FVuw3nY2YuvLfQwkMKozJW+n2TOnXRc3YXhkpBC0Z8iQ0ZLkG17
akfAEVrI9Url0ODhyewJtXsSpI2fzMa1G6gTHKcbuyFOoRl5s7VL2e5derPLP3BR
tYcoX96l+AHbxcEMFC2+mRod7nf56sFnVjR+ffxK8TuYiQVD/3YPaXXMV4P2rxRY
P0NLG87v5jlUi42a461YNLDYBd+/j7Vua43xkLwq2nLFIvsxs220jxXKdsLkP+0W
P/nc/bqMxVCDkD3qBtdKr6FYiku4mIprMflWputx/z+GJ1xyolz8Bt5qwdOppEOk
PLoA2XHxIfG0o4qbbbukjDXaFZl8/opGcVIpydzkD2wyWr311M6nIziPW4GDc+VI
u1gn26N+GAmrOE3rKTIl5sNfZ+CpvY3PPR8xTigWL8P7fptySyFjgILT3iPSVbMy
5aD6GJsTrn+OmHO3qBo/GUhUS8M+pP2ATCId+XbffeVMB1JAd4zShDHENXOdu40i
RBu5lcH3MINJDQ0uKVQG8pvc0FYRPKVr9ig/nckJapBm304S+mQ6E4QXe+GU/k8M
kfFPx2LFiKEWuO/i/PAf85xhcJg96vdHIKGzOrSfke+r7EKqo8B7U9tqoqmT/oO1
2Vn19bKr5V+xDkMoD6Ul4hE4xuxgKK14Dt2nszrVt+cZUq5RSnx95WDdKKKS/gLc
8vMLxyXoGRzbUuGpjoTne/h6h97K6nrdF51A7RWK62EXtINX4LvLqNrjyohTQ5+5
/xCR7iT5CI/J3rSPIerGfcZoM6664LsLIZOv78qYH7Vjw/GWLI5BuhGDg7u74YuW
GLtSSm/BOiAFpP77y/xZZC2+mCXEvcdLyKoNfacx7dK2Iknz7WTQKR9V5cfezxgk
cqKs/ZjAgsfR1m2D4b7wWUZPW5LXI2xCkGU3ehygFN6UHOuy75T7HSG2w5vYlVp4
bvFi8YXU1hXSLB6nh1sjgs3WsfvVlDL37dSm+BgKMRIenQ4Gd53pHl61z+tguWMw
rLYGDh9CuN5y0HSG6ZOcHx4HHJgPRNxN8MUY+m7t6NWgaVQJzGhEfOA7grCOVxss
YTSdnupo/nJLP1iFIihs6GW0pRKdK0KFsqACf3z3mrzk98X6SnxxtQLf9SejBCad
wH9kVrJMwF47vVyp2l//kMnpo3iir0RNbzjD8WpL80ku91BI9tMel+qwdxb3oho/
krbIBXcFFk684n94ZvBINOWH+tiiQ1VIzYczli5h/HqW4Ssrg9sL3E0uqm4M2+vp
jtk0IQhsq5dGyNejDbLEARWNS2tFfUoqtR/gGGtjYgnXimzfTk/tFgsmDRIgVCE5
xYvuvXgJ3ogpoHDeF+qmClanDwz721TNcISY7omeJ3KeaKchdvia9v6qdNM4tz31
IJrI7em5+SQHggifli79R5YmtN+FVIi9aDrDl+qOlpXrS6Y66hJKokYsqwXkZH56
myYdg1l0mIiYB5md+40W4DV8ttgP7y+X7Wugmqpbv8IOLp0+xAZGzJMBBRljfkT3
H/XEAgehzod+p190J4cabVpsTwqzuHEVu97gq7Jt1vc+OY4aJ1lP38HJVOtvvJ2r
VJYZ3jHYrQJ0lChexpOPd8/h6n3y8gTFG1L+OkXYNgQR5ecs/XfhE93OkLtfA+Zz
FXC31cNpxwi31wSpp1iiLA/hQPAfJe7sZZkL8uaVtSLr+OgUD3qqX1bWsLmUe/fx
z7YKr4aCTGqIgc1Ez+gVBztbtgtpiaHMRDVVfZPwcDzNpvAlJiu5/awS77mdJRt0
AFR9TtI+tGjh7BtG71Huy5w8tF66IxX7Uu8uvXtTaJOqJ0keavSWiP4tp+zz7wir
0+Pe3XQZ2njxCuLqb7xp5dZj6rAgGdhTfo/B/FVqCWBM8C817bacuDw7fW1SguMB
0TRhwdBw4iU2QAWxsmTvN+WQoZpt5lpwFdoCmh1Nr34n17Q2pVDxuiE2CUDU9pCH
kQ4eJHLPhqNPK8JeyNvxiWg3NQaiRE8wkdJYonGbe6OwNuLqVFQv6OgUikPYMd3N
jfR6cYDScxvmvV2F1D0nPICnfd40trxq7NKa3AdDNaLmk5Mj0CWvPrSf+DTARWJA
0C8TCIBnEQGKu8lSBw5aDU6RYoCEcVabh05uk16q5ixtVmi1qK91mZUmHPTfFuoq
5y85cfEFyMY1zIWOPUKpoloVk3VKqoVJPE1olx28EOVgc5Bh3tBeBKGvAwivmjwk
NubiXWeG/FRjyxTal4SsJQXN7HZGP/ZtGrdO6kLnnUludS9iABSRqLVYmpfNd5DI
u+jLniucew174SO6ZjigPH078+GRiED3KkbxSlTwk/xK4hSWhx7dlqmbHYWigmWe
+OwTy6MTiNSdsOmhjtUBidPRCF4Ur6UoFikYkQT8tU5QenLTvHC1zOa4uIq3VVpD
xAORekog1Xgt5VIGVWrOyhG4pJ5eCim/qgsaUmYBdXoAIbYbzpLOCk2KgCtsinZm
8ZBDBj2d7jv7RUfSsxDQY7OSJseWlvNRcz6uM2XLVLA7bKU/2OKtrMe+GrJQ47Uk
Pc4j4uGKiKPmvHqeVpL+mM9ufQwoB9cf5ldOL6wCAbADx7aYkKoSCTsXNe9RaaOP
C0p1p4TnLVt0CipgzA0fWmFcG9DwqELL7hXGNRlUpSZuyPq2uMZDzzMIClLa3KYW
p8I0M9zHnY1+dYTtJPZgSGM/He9eyazP3T432pNkimv9/i0Uc1EsCX4z9TjIexwC
IKG6PSpGpmScY86Yh75ewsaA4nSWI/9bGJujJ8aPZLs7ECW+KO00SusNsn7afjLF
wmdHshTlW7ui4dnD3rk9I+G3cF1+YCeTZFVM3fNJyMIt27c5tSgy7epBuwrycVU6
Osgek8xtfnPvZhNfn5OVpNaPbsKMl0IeuGYL2E5l4r2AL5yGXx/nGjPMiP11P7Hj
fnr11Yzy+Bd9fL/W5qF2dPxZRqFyTGSEv9qF+4NaZmOEyu16yGKhXtkmiXynxHHg
j44KO/tL+L2PT/yPSdyA2QjJSSgGuuOQZtJSnmafRmWnW9H9SOUaH/kmtBfC4mmH
ltrq1DKdSEZJe1nK873Md5Q79Ci8jLB/5wto5AOhREPMWpPhfYPbpPNjsDMzEmCK
XxWMDaaYwAv94oqTb/n+FNVxbo0JJZt+RwP+CXjQ7vGzY4DqOMzfz+U+iNYS1P+F
vxGPOgm3Az94xJWpNZ1LUO3LuPitGMOB6o/gCfxzr+FoR/u9tq87q1d57eKDcXfr
BUkdD6Ni3REx/huLbj71pFEvvcPOhjMerHf/EUxh9sqhLgQqK1E5VtudEz6pqF0P
Z2iSmb43V/U+MNqV3wfJ8r3nf9z1AlK7iRlh1O9O3SZnD1Us6LEbJ1WyEEjQjBJ1
qD46llLFuSoniYBZdCxQU/yKRatQloZMv8b9D6LjhiY18EPwIsjipHPKOVzHEnmz
bv7tflLP6gwwnMt5wCVMkRUZ77rAHpHegAkW4haTKyRPPE6636C0MSCeF5JJJNe0
bgoeXRJJOAiU5A1RLXwh0so8wUnehxH8VECM6rSBncY471bgnOW2facokE4KuWDL
ywGr5FZVXf/e8rjEHxBuvfNp+WerJmKYFg/tXhA+5O/vEidBp4ujeDbsvBdHntmS
Imht/DqICW+ldxDRtl1BRu8nHi6+OEEjHrR/618yAUtzkiMOV1FzLMBNFlWyCXGZ
bSXsGiCsNHHtUnNwzsHQKuhgITllbg9HC76kZdlw8yPU5idv5MDQqMIJakE5csO+
XqKfbkIuItXXQA+etiCtdKe5whKJl1p+NYCMlir8/2NDJlSCwLL0gG3CuvGcUHod
bwneCnFm6sKPSnFgL16gXYgsu/J1V6Inwh4HgJCV8rxvJCmdn/NylJyOdyx++wOY
f84jn4R/zuQuLhM4LRTrq0CSb8YBZwbgiMvvlhGOI7e0EyG8cYt+vZ6HIsDUJM4o
zzZ6jF7dWGtP+fDOCxsZM7lSeenWJ37SO3aN0kRqepq076p4WK+USWP4k31hPNvs
1Z3zI2B2A8Hq7KaXvcOUPRfXXn1lUYFYk+Zx/ISlJ8QJI4dg1a4tyq/nCUYkPNS9
l8jgLhKjliBeSyN0T6RcnjUIv8QAUCEtfjDQr+QS5VikVW6rXv73GFgY16p5qM/A
VWH4KD3WlJB2QkqUJG/QALrnNKUNIHR0jgSf7jJClPnLyNKpA0eEqYDs5nV/hMJL
bmCfTLa1oBqC3woqY1/zSTWHHK5d06+BkU153G0PA0MpPFoqqDvSGV/k57VU0VXL
lc6w86428FH6SKOlX4NzkF4x0319MirjD8diN7gat6s/0B8H7T0TKv+2Xxupp5Dl
G8aR2oYw/lsEU/JA84JYKky6CwnfsqgDxcMZCqeZfMP9NDTF9kgtpxpn/5j4UhPS
Oq3P5qh3lTr2YUMCcV6GhKL3+yirr4PQpr3f0PcijVi9rovNrXn5vBrmmcW/nVIi
K+kVNgIYYB64i1cLY9J83/VAplqWqbvISjhgTC9VV8f8ldTnMDUPxP44ocfIU9Fk
PkVfcQOjlvltAewfSKiroODhsuH2W6WL5CYKv14at/vZ268EmVF43Dumo+8xT5Gt
QUByUrrMepuCrPhxpfrUSN3U4Dc9W1v2/6M+TqrCS75JDmJ/9Ny6rdAWBcZBJudV
O3eKfv1bMnV9/qbonpxg040d/+7Mz1DjGQK8jvyJOLQloC6ggtCQPY4svCUt6hwC
DPZUw7Jv758ULmo8evmTVcikBPnmguNG4SyM8OAf8suEcqQfmYLzOXEYCA9tK5PJ
kUZoCsF0G2yiMqzjqh6ojiZHGxeZ4QhK1La+Q0DSYZknEqcfLwJ+FD/7GZjWrS8D
0N4v/eSyiZPXCJgQkYWup2m0exVU/QSQSkkfD7pheYAmB/pAVqe/Lc2iH0zqj+z1
Sf6lEPUW9N4plXOcQ/eaw2BExFJJExvP90nqm+kBxNH+z9QH4B7MHixV3s3ucRgd
0iVGsn9UX24RfyTxhJfSj2pbSKMYSQtA0Y726OSZpYz1dZx70kAtZMW9NmlkRL9T
Bv3DAtdi8nNK2u8E6M48wigNuWjUy8uEUa37rz41He15HOXMxccjGI4S79XwpuXj
56pc2OKDcKuEYbFC4tjhOYiR1z/APLyWKqHXHClRGJHUEdFGQfs0VVn5BEz4ZKYV
`pragma protect end_protected
