// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:09 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZdiWxcS6I154Uuu30uB9uv2KD0a5irVdCLvPf0xo8ju0BtxMnG2f7U0exBBClVCq
PoA6ws1Yrss14fkQO4CI+8+hmJbW9QoeK8FrUNdjTL77v1o5RGi7vl4P1AhEAR03
3ktn9NLIA12IwTkNw98lTUxgSpVQ3FnOATNxTDkQ3/A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4208)
2W66pKpbIEfPpJ5mhyWL3WvpczmlnJip06NSg77UVBhZ+6e7WdxFOQpo9I5Nb5La
LxFhAYO+nESsYRY0rI0ebNfGMlx5pGlbOCH+V/bqFWE19zuH1lScBFnp4kFJcSaB
3boaqZv5NR4cjFow81VM8sqLM3M4OLqU50rCrOZf+Afso1QZPbtX2R/7mfu62hBe
yOpBZyvueYdeQif8ZjuVlJPLItMPaAeupvm60x4Dnj+ltN9cBp4MeenWyiagN9v6
GjPfthhjWJuImZ9Zf0hihYKpyatR8d9BuJ1ZgYMmGnJvzvyI4BH9WYWZFJPYfZ2n
INGhKM0wb262XTXQg7tQS/lL6CHW9FZPBgeiSazCN9gyELcIWBpWIiiDa1pl3Pe9
FqdRI1xSjJvWlE0KRCxGvBgMRud4UbB9p8Zqk5ZPLVDBbcq28EgeNOMNPm21rqN1
TH8BkYav6me6J+31x1PHxoXQ5QFDnoFQzgq1+Hn3btpxdVbsUfDMm66CUjYmDIZz
+8xPQdFUAxCFJyUG95JNO3f36B/j2LcYJIAEOxFZ9bPtRlvv7Sfr/rJ/T7Y+zfG4
UzOVh5x3hVn22nUaaEiJBlaCXexU2lbJHmxPsuePiIrlfW5Cjb6JSiTeiLz1rZp5
1XYPNCRq9sx5SfDINnshBHSIq2ArCNxJhfikkaAyT6la9e1jFeCzanzPPQT6w3Vm
8ZOkl1leMMRP1rzWJbq2lMPjco81Zy3vQ6dUGTq7dqar08h66TnKnlAX4IK88ZC8
0FLGaBn2+tZHns/V/IDpFi8YcISfebLWhP1YO59PlkITLymrnrSFdEQgf7taAMN7
M4Xv2jqi7CrwMOztR10u16a4AxbzCavWKxeznxY2ZBQsTQ0+4PTWu92/8mQ+3DwD
aX92PikvLBvGq+1SQvUkDj7mM8akQ/ChdUVYwLnDcKpQyAkpcA7JDYzgICygukyu
dlHosnCCtxMIfx51j1CvYkINwjnaFaVM3Nb50HHVbw9C9hUHE4zTd+2avJ/USd1n
3s6uTbnAPomdRMqo68c2hsNeRM7qaS93693gahCTYPIXz9ab6cw24ZZmm5NIdinC
XcY0oj1o/15hNcefjKhveaEeR61wCDda+OtgPndLx7VHwsYCvJ+kMRdQtpWmrDin
L4EAntmgBRbJgDjCiJIOomajrpGWmMfzsNdtA4WWGQf/HS6g9Svef/9aGZs+nxy8
pQRViGnfFmT3btg0e1dt5xq/plWWHSjsSzCtXRNoZNb2jzpuHjdGhEqpvc3yIgAb
f+1EptHlMd7HPTWUV3CFFCWIkNsBdkqdAwZhjEec+tvjtiSfMHn6Z5X3v2qL05BI
pMkH74eeocAl7GAT8hAvvwSUfXfW33T/qBowOKnX7D9gu4Vn1OnkbHeg3AeSmmh0
j6M2Iy/QLgA64cfGAP05tbHeMtauDjgccNnHsdnATeZYEKwdquLYrqcsJdEq2CzC
HY5Rm4+bvLf6p1LrFwpeFu3BiX8KtU9XcaJm6hum7ZwiiD8afxa4eFy46zRAl4mx
LeFgJASW8pHRmSYgGfazi9KYwSyrzebpiJSpu0gELvgkwiaoYuoLiGxXu1oQyFdP
JY7m2B0DUHDFTHHkmOYQ5zTCQtNFPU3H4VGsY6JzZWTy6PRs3xsSP2osi2HxUZ/t
31EPoE9AiTDXG/WY1+H94cQjU8NnjE6vAWNR+tF2cudEUuZh4WgdC7Q5uxnnx4df
+HrmIzMWnXgPpkbGgUOk7fWHKQ/4AQ1DXq3H7jsYr3d1zwZrzfchg1FZCYVIAGQI
iYQ8RmVBPvW0BmbDcgeOJQllahoSzu+XRuFVIVCn4Do3Lr/2uhzofpT0hBWOptJt
7Fh4iNZOY2ssm0eW391BI6/QN7nQEbK/lU8r0PE2eVqURoV16lb1MSpwCHuOel1R
7MualTHLrELRPdUnj8Vi42NGXxAglwnurXD59Z9bbd1HjvacW+6lV5elxBgEISjS
iU2b7rnuDtwIQ4VOz9livio1rkuIJnIXEWtRhlYWK3Bz9AjkUJbFMC4pJ9X79BAo
Bbn9mjrtxLwUVkMK4EWmCEMt7HzoE71Zr6KggGO6sMgwVt0iE2jkvXMmRJOUE7KG
TSQ5bujiLPyoM09LpZ4D3JseCq9hl9522rdglzJEKBcHDmH0bJ+QGeK+hntaWGcL
PGY/akqi41VmOlxkoSHaiCZ7nCshk1r1UrxKnl8+PggJ2KvxowrItcsDBJKa7tSk
vLCIvii6707vXnM8mTIroxG+5R/EsHFF2ydAzcEvre0N27Uz57kNfsSivPqNLeu6
yYkdAX5Vu6fFa4RPlWDb7gZXGk1tyHhB5pq+UHWqbSCHc/SrqSxgLvAoxo65De8q
t4MUgST6Ca9YznrYJVbFo9Uob+z2nU4cQ0yDAzDyXdFupNQhItn5vZzwkie9ejJi
OSp7EYXbeNY74muiuYp2WZ65r6KaaeLrBYbaPjgfFalwplYhDydvr5Bhdt+kqYHm
5d1BJ7Vi4S94FQj7UKApOIRU9XQDbF6cdlWQN3vkrtU/C/b+qoq12JcRuk5ZCwx1
w4KQcw74X8KZnJE1XcjO595bPuRFhcQEjJAX1TQzb55Ay2HHflW/6ixcSfsM9kCH
SsW1a7kIjep+OzyqGxfEY80E3k7wq2/EEi2saJ1+At3u3qUmejE4KlQn1UIyst8A
vta2HzjsoMsB2UxlJi6PlRAiRvCHw2msW3XB4nnnds7EOJuEaM0LKn1Aws0x8Pyl
qY1H5XdIpg7kDhu9eu4nfY7WG7TMY5MagRaEfZtSCu0dYcO2RbtBs1cb59SWtMPV
OvflUP1r1UT/l8xuEqdtnOpDDzOfB8dopn+R2cwUS40u1lrEn0GT+DkMh/tTb9e+
hxw7P7cDxhPfE7T0IhwKXnz3Xd1As9Ofu1DXNOiKsEFeOEmQZjFq4CkP3CTLd8M/
ziUJo0kvqgNM4aH0htUc/Kb7Ts2V/ydczNddGseh+Cr4BZJ9jSPJlAvT4ujlNIrU
QxFsAlVLezPYtJZe4IIO3GZ7oMQtdK+FKk5NMD+jSAgxeydeS7X+isSwKY8F8SwQ
2V7I1p1TpN8ZceWo6cTB9wCi0KkV+Iln9mwnNOCOVUuQFIx7Zec+6YzwcN5xZpra
VzVrq1DzsrOP5+76V1+Lzbc9KTR7Eh9kyjvCSSudM8Mj+jVlTqEvYPhJ1VxGssMi
6jvCHCPW9HFvPqasm6jdTiunj3iEUl+KFwd6xIgE9jbFZsI6vUmMevTF/Kzr2SUH
siyp9PvTweki+FvrNpfRB8iCgiuQMovuK6aAslYjpmoU0bIFZSXEXMvCaivG7VUh
KSWP7d/IuPH++w9w1LkcD41mIb/OkbzXVSz9HV/jNTP3+8N7s+SI4QSLuae6RGwI
3jA+k0tMrndZ5hKgqBXzS5EB3LK4kGq4hJabJBJzfTxKtO6fTIl7EwH9ccETKfzH
kwCaq2cPhKS0AYar/f6trfIAdm7P+6dokybMesrop4SWIg+5U6s2Xr/JUFNNXftJ
PbZLxPlLGXZN9HxBTw0XX7eo0ucB/jTpC9hLVfHJDsyiYOOXSaGdwxNM9071Y93z
bvSzoCH8ooXvMRrhbpN5B4v+OuSL1MyccxqAEZsz35+FE+iQoV+H0hkgxAVC+tFZ
4EvKkBIr8pljOOlb9GQWJ+foxkpEEo8rPEhiL/IW0f4OYlcA2b6pAtroeeif3bMn
k152DQkylBQceahQPpvH8a6Ovj1dlRVuy7pklyEQS13BB5V2Qkr645FczKH69k3f
GzbuuXk3kZqJTLft+YP2nuhFh/g7E4X2Z0ey3/02z74BvEBi3rcFKAuCUSsMaWwk
DaW7YgP3vmXJp6ca7prlICW8OTspDhUvULMFTerZBcBxlcM9L0feJpuzsjgNTVSX
aDsFx39Sbb0+KkCq0eh05nOffY7jqo+t2/nMJjEMlMtuVJdF4efQwbFAMfRRErQV
Su/Vwxv+Z8eY/2Ta63sdeNTu2dqEv+GAgkC/9ZCY9no9OZAEXgTTq14C2UZycAwZ
6/Dy0dC/TQRUMHz3TO7Adzf48FWBRnOawXpXa4uNexFhZa4d7YUbQsU1ZlMOzbjU
2+XZx3psWj7Ey+w7LaK9kn2XsIbOGMuHKGN7dIYl53jEQ/I4bmaeoABJdbXlbihQ
PtcBfnbM/XdT3686zJEimPOAMppIwlfj5bsX98FTz1w5/JjyDO09//Dinfi/Ak8J
iBdnMOdJbn9snGSJF+CsvLKFK2QNNWDbwzLvuAPj7eHigFMaU9On93rhB7hobCew
MiryBPmyv1iQ/DITXIgZ+nyx6UMIdtqWKCncflYUvPJIu9MTurhr1rHqUGeItk3v
EGp3rMes71B3iHFYqReqlA1RrlVxSxC28a/ag7pP+6yYvPzHAl39er9Gix5NHQFL
YlJhPnLaseSGczocHJIxe7r/PvwODMXnboFCXvcViezDK4P+rF0nvw7JD2s2tm0/
y0PWVt753paT4xipvg6TlPYiQVqQ+HIsKAumCWfihACn1Y3HRXw2Pg1tnA10agMn
IADbiCTRbUpwL5Lm9nf8HyGpyIDcAEObPeR5GR+saB/cNbrhXeFjY3JYLBJFiC4j
/0LPPZTZHx6ZVXj9p8yOnkUkxQqP3MHo5XJ+E1Ig8mdsA2AyAoSC4i/9QiHjr5eO
9szjv7rQOdOsK0R0n5zHlGxnyGTYBHkO5jQuF4879wpa1+0Oe0vVeh5EUX1nQ+nl
BcUxPmia+DlBYGw0+33Apf8A9JGMi88NpescWLcn6afgiTlJY7EZHS3sFZ5bbc4p
zst/5Gbf8nFAe+9HM1ivn4sxAD7A4WtV/GB9ZH/fhYnk3pXKUzlYu9c3QiCeu5iR
lYs26Br1/NjVK1POufL7c95v1r+ry6HYg9OER29KfGICHLqpQXb37QnK2kgMpRoc
vE9/818jn7IKqs3HrEz7F8zinJe3NjyUZbkF4h4G8O6YV0KbQUfskxoFwVs6P19Y
tqaqAZGURd/KPOhusms+u65SgJHyKPRwuh/pOjgsD48724oBCsUv4LlRVku73/9z
ZUwmJ3W1Ebrbh1Dz5qA1T8WfnmsMrR2YroWNrpD0ddHSU/obFQtI+wxchvdNLdYD
vJURjhYI91W0NJYsMZPlWDpfOSvJIyeuRdQu63OcpcEIY0M7IzA4yRRWcrUMG1dE
ilBbwXIq72OPS2YDfuf0wtaluTkqc5C+eVQEScnnpQohvgneifWf+c6yqmGKn2/M
pwQFUZJWBA15gxtKaFy2wVakhrbQ5Eppv2THdzEb41y/idQ9XlukjcmcVZd2RlCz
xmMo37ifF2oM6Wbi2POvHLrMrDxupxpplcQ2xq90gqPejau2pN4hj1ltmxXGNhjR
/4mRZAT/ysep5PRQWZ2dSjBZzV40ZbsnURzX0FtbPYQ5t5Mqm7fqKM+G/YIDh8OQ
ZGxpySEGxV63fs5X2rw0dQVSy/4xA6kPk7pyIjp5O5gBIvTJIvOMYFLgEPNwQnQu
LREPujOoLrqdmYQDwIoTk9iEfg0AL7SNTReappsQUyCqijwcgUrXpfwDJSB+q51L
bfQQ0ZpSeA6v3GwTMU41v0QHn99088Z5IVeEnxkyVoQ=
`pragma protect end_protected
