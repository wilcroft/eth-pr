// eth4to1.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module eth4to1 (
		input  wire        clk_clk,                      //             clk.clk
		output wire        clk_312_out_clk_clk,          // clk_312_out_clk.clk
		output wire [63:0] eth_in_mux_out_data,          //  eth_in_mux_out.data
		output wire        eth_in_mux_out_valid,         //                .valid
		input  wire        eth_in_mux_out_ready,         //                .ready
		output wire        eth_in_mux_out_startofpacket, //                .startofpacket
		output wire        eth_in_mux_out_endofpacket,   //                .endofpacket
		output wire [2:0]  eth_in_mux_out_empty,         //                .empty
		output wire [7:0]  eth_in_mux_out_channel,       //                .channel
		input  wire [9:0]  ethpack_tagin_data,           //   ethpack_tagin.data
		input  wire        ethpack_tagin_valid,          //                .valid
		output wire        ethpack_tagin_ready,          //                .ready
		input  wire        reset_reset_n,                //           reset.reset_n
		input  wire [71:0] xgmii_rx_data_0_data,         // xgmii_rx_data_0.data
		input  wire [71:0] xgmii_rx_data_1_data,         // xgmii_rx_data_1.data
		input  wire [71:0] xgmii_rx_data_2_data,         // xgmii_rx_data_2.data
		input  wire [71:0] xgmii_rx_data_3_data,         // xgmii_rx_data_3.data
		output wire [71:0] xgmii_tx_data_0_data,         // xgmii_tx_data_0.data
		output wire [71:0] xgmii_tx_data_1_data,         // xgmii_tx_data_1.data
		output wire [71:0] xgmii_tx_data_2_data,         // xgmii_tx_data_2.data
		output wire [71:0] xgmii_tx_data_3_data          // xgmii_tx_data_3.data
	);

	wire         ethpack_packetout0_valid;                  // ethpack:packetout_0_valid -> avalon_st_adapter:in_0_valid
	wire  [63:0] ethpack_packetout0_data;                   // ethpack:packetout_0_data -> avalon_st_adapter:in_0_data
	wire         ethpack_packetout0_ready;                  // avalon_st_adapter:in_0_ready -> ethpack:packetout_0_ready
	wire   [5:0] ethpack_packetout0_channel;                // ethpack:packetout_0_channel -> avalon_st_adapter:in_0_channel
	wire         ethpack_packetout0_startofpacket;          // ethpack:packetout_0_sop -> avalon_st_adapter:in_0_startofpacket
	wire         ethpack_packetout0_endofpacket;            // ethpack:packetout_0_eop -> avalon_st_adapter:in_0_endofpacket
	wire         avalon_st_adapter_out_0_valid;             // avalon_st_adapter:out_0_valid -> eth_in_mux:in0_valid
	wire  [63:0] avalon_st_adapter_out_0_data;              // avalon_st_adapter:out_0_data -> eth_in_mux:in0_data
	wire         avalon_st_adapter_out_0_ready;             // eth_in_mux:in0_ready -> avalon_st_adapter:out_0_ready
	wire   [5:0] avalon_st_adapter_out_0_channel;           // avalon_st_adapter:out_0_channel -> eth_in_mux:in0_channel
	wire         avalon_st_adapter_out_0_startofpacket;     // avalon_st_adapter:out_0_startofpacket -> eth_in_mux:in0_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;       // avalon_st_adapter:out_0_endofpacket -> eth_in_mux:in0_endofpacket
	wire   [2:0] avalon_st_adapter_out_0_empty;             // avalon_st_adapter:out_0_empty -> eth_in_mux:in0_empty
	wire         ethpack_packetout1_valid;                  // ethpack:packetout_1_valid -> avalon_st_adapter_001:in_0_valid
	wire  [63:0] ethpack_packetout1_data;                   // ethpack:packetout_1_data -> avalon_st_adapter_001:in_0_data
	wire         ethpack_packetout1_ready;                  // avalon_st_adapter_001:in_0_ready -> ethpack:packetout_1_ready
	wire   [5:0] ethpack_packetout1_channel;                // ethpack:packetout_1_channel -> avalon_st_adapter_001:in_0_channel
	wire         ethpack_packetout1_startofpacket;          // ethpack:packetout_1_sop -> avalon_st_adapter_001:in_0_startofpacket
	wire         ethpack_packetout1_endofpacket;            // ethpack:packetout_1_eop -> avalon_st_adapter_001:in_0_endofpacket
	wire         avalon_st_adapter_001_out_0_valid;         // avalon_st_adapter_001:out_0_valid -> eth_in_mux:in1_valid
	wire  [63:0] avalon_st_adapter_001_out_0_data;          // avalon_st_adapter_001:out_0_data -> eth_in_mux:in1_data
	wire         avalon_st_adapter_001_out_0_ready;         // eth_in_mux:in1_ready -> avalon_st_adapter_001:out_0_ready
	wire   [5:0] avalon_st_adapter_001_out_0_channel;       // avalon_st_adapter_001:out_0_channel -> eth_in_mux:in1_channel
	wire         avalon_st_adapter_001_out_0_startofpacket; // avalon_st_adapter_001:out_0_startofpacket -> eth_in_mux:in1_startofpacket
	wire         avalon_st_adapter_001_out_0_endofpacket;   // avalon_st_adapter_001:out_0_endofpacket -> eth_in_mux:in1_endofpacket
	wire   [2:0] avalon_st_adapter_001_out_0_empty;         // avalon_st_adapter_001:out_0_empty -> eth_in_mux:in1_empty
	wire         ethpack_packetout2_valid;                  // ethpack:packetout_2_valid -> avalon_st_adapter_002:in_0_valid
	wire  [63:0] ethpack_packetout2_data;                   // ethpack:packetout_2_data -> avalon_st_adapter_002:in_0_data
	wire         ethpack_packetout2_ready;                  // avalon_st_adapter_002:in_0_ready -> ethpack:packetout_2_ready
	wire   [5:0] ethpack_packetout2_channel;                // ethpack:packetout_2_channel -> avalon_st_adapter_002:in_0_channel
	wire         ethpack_packetout2_startofpacket;          // ethpack:packetout_2_sop -> avalon_st_adapter_002:in_0_startofpacket
	wire         ethpack_packetout2_endofpacket;            // ethpack:packetout_2_eop -> avalon_st_adapter_002:in_0_endofpacket
	wire         avalon_st_adapter_002_out_0_valid;         // avalon_st_adapter_002:out_0_valid -> eth_in_mux:in2_valid
	wire  [63:0] avalon_st_adapter_002_out_0_data;          // avalon_st_adapter_002:out_0_data -> eth_in_mux:in2_data
	wire         avalon_st_adapter_002_out_0_ready;         // eth_in_mux:in2_ready -> avalon_st_adapter_002:out_0_ready
	wire   [5:0] avalon_st_adapter_002_out_0_channel;       // avalon_st_adapter_002:out_0_channel -> eth_in_mux:in2_channel
	wire         avalon_st_adapter_002_out_0_startofpacket; // avalon_st_adapter_002:out_0_startofpacket -> eth_in_mux:in2_startofpacket
	wire         avalon_st_adapter_002_out_0_endofpacket;   // avalon_st_adapter_002:out_0_endofpacket -> eth_in_mux:in2_endofpacket
	wire   [2:0] avalon_st_adapter_002_out_0_empty;         // avalon_st_adapter_002:out_0_empty -> eth_in_mux:in2_empty
	wire         ethpack_packetout3_valid;                  // ethpack:packetout_3_valid -> avalon_st_adapter_003:in_0_valid
	wire  [63:0] ethpack_packetout3_data;                   // ethpack:packetout_3_data -> avalon_st_adapter_003:in_0_data
	wire         ethpack_packetout3_ready;                  // avalon_st_adapter_003:in_0_ready -> ethpack:packetout_3_ready
	wire   [5:0] ethpack_packetout3_channel;                // ethpack:packetout_3_channel -> avalon_st_adapter_003:in_0_channel
	wire         ethpack_packetout3_startofpacket;          // ethpack:packetout_3_sop -> avalon_st_adapter_003:in_0_startofpacket
	wire         ethpack_packetout3_endofpacket;            // ethpack:packetout_3_eop -> avalon_st_adapter_003:in_0_endofpacket
	wire         avalon_st_adapter_003_out_0_valid;         // avalon_st_adapter_003:out_0_valid -> eth_in_mux:in3_valid
	wire  [63:0] avalon_st_adapter_003_out_0_data;          // avalon_st_adapter_003:out_0_data -> eth_in_mux:in3_data
	wire         avalon_st_adapter_003_out_0_ready;         // eth_in_mux:in3_ready -> avalon_st_adapter_003:out_0_ready
	wire   [5:0] avalon_st_adapter_003_out_0_channel;       // avalon_st_adapter_003:out_0_channel -> eth_in_mux:in3_channel
	wire         avalon_st_adapter_003_out_0_startofpacket; // avalon_st_adapter_003:out_0_startofpacket -> eth_in_mux:in3_startofpacket
	wire         avalon_st_adapter_003_out_0_endofpacket;   // avalon_st_adapter_003:out_0_endofpacket -> eth_in_mux:in3_endofpacket
	wire   [2:0] avalon_st_adapter_003_out_0_empty;         // avalon_st_adapter_003:out_0_empty -> eth_in_mux:in3_empty
	wire         mac_0_rx_st_fifo_out_valid;                // mac_0:rx_st_fifo_out_valid -> avalon_st_adapter_004:in_0_valid
	wire  [63:0] mac_0_rx_st_fifo_out_data;                 // mac_0:rx_st_fifo_out_data -> avalon_st_adapter_004:in_0_data
	wire         mac_0_rx_st_fifo_out_ready;                // avalon_st_adapter_004:in_0_ready -> mac_0:rx_st_fifo_out_ready
	wire         mac_0_rx_st_fifo_out_startofpacket;        // mac_0:rx_st_fifo_out_startofpacket -> avalon_st_adapter_004:in_0_startofpacket
	wire         mac_0_rx_st_fifo_out_endofpacket;          // mac_0:rx_st_fifo_out_endofpacket -> avalon_st_adapter_004:in_0_endofpacket
	wire   [5:0] mac_0_rx_st_fifo_out_error;                // mac_0:rx_st_fifo_out_error -> avalon_st_adapter_004:in_0_error
	wire   [2:0] mac_0_rx_st_fifo_out_empty;                // mac_0:rx_st_fifo_out_empty -> avalon_st_adapter_004:in_0_empty
	wire         avalon_st_adapter_004_out_0_valid;         // avalon_st_adapter_004:out_0_valid -> ethpack:packetin_0_valid
	wire  [63:0] avalon_st_adapter_004_out_0_data;          // avalon_st_adapter_004:out_0_data -> ethpack:packetin_0_data
	wire         avalon_st_adapter_004_out_0_ready;         // ethpack:packetin_0_ready -> avalon_st_adapter_004:out_0_ready
	wire         avalon_st_adapter_004_out_0_startofpacket; // avalon_st_adapter_004:out_0_startofpacket -> ethpack:packetin_0_sop
	wire         avalon_st_adapter_004_out_0_endofpacket;   // avalon_st_adapter_004:out_0_endofpacket -> ethpack:packetin_0_eop
	wire         mac_1_rx_st_fifo_out_valid;                // mac_1:rx_st_fifo_out_valid -> avalon_st_adapter_005:in_0_valid
	wire  [63:0] mac_1_rx_st_fifo_out_data;                 // mac_1:rx_st_fifo_out_data -> avalon_st_adapter_005:in_0_data
	wire         mac_1_rx_st_fifo_out_ready;                // avalon_st_adapter_005:in_0_ready -> mac_1:rx_st_fifo_out_ready
	wire         mac_1_rx_st_fifo_out_startofpacket;        // mac_1:rx_st_fifo_out_startofpacket -> avalon_st_adapter_005:in_0_startofpacket
	wire         mac_1_rx_st_fifo_out_endofpacket;          // mac_1:rx_st_fifo_out_endofpacket -> avalon_st_adapter_005:in_0_endofpacket
	wire   [5:0] mac_1_rx_st_fifo_out_error;                // mac_1:rx_st_fifo_out_error -> avalon_st_adapter_005:in_0_error
	wire   [2:0] mac_1_rx_st_fifo_out_empty;                // mac_1:rx_st_fifo_out_empty -> avalon_st_adapter_005:in_0_empty
	wire         avalon_st_adapter_005_out_0_valid;         // avalon_st_adapter_005:out_0_valid -> ethpack:packetin_1_valid
	wire  [63:0] avalon_st_adapter_005_out_0_data;          // avalon_st_adapter_005:out_0_data -> ethpack:packetin_1_data
	wire         avalon_st_adapter_005_out_0_ready;         // ethpack:packetin_1_ready -> avalon_st_adapter_005:out_0_ready
	wire         avalon_st_adapter_005_out_0_startofpacket; // avalon_st_adapter_005:out_0_startofpacket -> ethpack:packetin_1_sop
	wire         avalon_st_adapter_005_out_0_endofpacket;   // avalon_st_adapter_005:out_0_endofpacket -> ethpack:packetin_1_eop
	wire         mac_2_rx_st_fifo_out_valid;                // mac_2:rx_st_fifo_out_valid -> avalon_st_adapter_006:in_0_valid
	wire  [63:0] mac_2_rx_st_fifo_out_data;                 // mac_2:rx_st_fifo_out_data -> avalon_st_adapter_006:in_0_data
	wire         mac_2_rx_st_fifo_out_ready;                // avalon_st_adapter_006:in_0_ready -> mac_2:rx_st_fifo_out_ready
	wire         mac_2_rx_st_fifo_out_startofpacket;        // mac_2:rx_st_fifo_out_startofpacket -> avalon_st_adapter_006:in_0_startofpacket
	wire         mac_2_rx_st_fifo_out_endofpacket;          // mac_2:rx_st_fifo_out_endofpacket -> avalon_st_adapter_006:in_0_endofpacket
	wire   [5:0] mac_2_rx_st_fifo_out_error;                // mac_2:rx_st_fifo_out_error -> avalon_st_adapter_006:in_0_error
	wire   [2:0] mac_2_rx_st_fifo_out_empty;                // mac_2:rx_st_fifo_out_empty -> avalon_st_adapter_006:in_0_empty
	wire         avalon_st_adapter_006_out_0_valid;         // avalon_st_adapter_006:out_0_valid -> ethpack:packetin_2_valid
	wire  [63:0] avalon_st_adapter_006_out_0_data;          // avalon_st_adapter_006:out_0_data -> ethpack:packetin_2_data
	wire         avalon_st_adapter_006_out_0_ready;         // ethpack:packetin_2_ready -> avalon_st_adapter_006:out_0_ready
	wire         avalon_st_adapter_006_out_0_startofpacket; // avalon_st_adapter_006:out_0_startofpacket -> ethpack:packetin_2_sop
	wire         avalon_st_adapter_006_out_0_endofpacket;   // avalon_st_adapter_006:out_0_endofpacket -> ethpack:packetin_2_eop
	wire         mac_3_rx_st_fifo_out_valid;                // mac_3:rx_st_fifo_out_valid -> avalon_st_adapter_007:in_0_valid
	wire  [63:0] mac_3_rx_st_fifo_out_data;                 // mac_3:rx_st_fifo_out_data -> avalon_st_adapter_007:in_0_data
	wire         mac_3_rx_st_fifo_out_ready;                // avalon_st_adapter_007:in_0_ready -> mac_3:rx_st_fifo_out_ready
	wire         mac_3_rx_st_fifo_out_startofpacket;        // mac_3:rx_st_fifo_out_startofpacket -> avalon_st_adapter_007:in_0_startofpacket
	wire         mac_3_rx_st_fifo_out_endofpacket;          // mac_3:rx_st_fifo_out_endofpacket -> avalon_st_adapter_007:in_0_endofpacket
	wire   [5:0] mac_3_rx_st_fifo_out_error;                // mac_3:rx_st_fifo_out_error -> avalon_st_adapter_007:in_0_error
	wire   [2:0] mac_3_rx_st_fifo_out_empty;                // mac_3:rx_st_fifo_out_empty -> avalon_st_adapter_007:in_0_empty
	wire         avalon_st_adapter_007_out_0_valid;         // avalon_st_adapter_007:out_0_valid -> ethpack:packetin_3_valid
	wire  [63:0] avalon_st_adapter_007_out_0_data;          // avalon_st_adapter_007:out_0_data -> ethpack:packetin_3_data
	wire         avalon_st_adapter_007_out_0_ready;         // ethpack:packetin_3_ready -> avalon_st_adapter_007:out_0_ready
	wire         avalon_st_adapter_007_out_0_startofpacket; // avalon_st_adapter_007:out_0_startofpacket -> ethpack:packetin_3_sop
	wire         avalon_st_adapter_007_out_0_endofpacket;   // avalon_st_adapter_007:out_0_endofpacket -> ethpack:packetin_3_eop
	wire         ethpack_transmitout0_valid;                // ethpack:transmitout_0_valid -> avalon_st_adapter_008:in_0_valid
	wire  [63:0] ethpack_transmitout0_data;                 // ethpack:transmitout_0_data -> avalon_st_adapter_008:in_0_data
	wire         ethpack_transmitout0_ready;                // avalon_st_adapter_008:in_0_ready -> ethpack:transmitout_0_ready
	wire         ethpack_transmitout0_startofpacket;        // ethpack:transmitout_0_sop -> avalon_st_adapter_008:in_0_startofpacket
	wire         ethpack_transmitout0_endofpacket;          // ethpack:transmitout_0_eop -> avalon_st_adapter_008:in_0_endofpacket
	wire         avalon_st_adapter_008_out_0_valid;         // avalon_st_adapter_008:out_0_valid -> mac_0:tx_st_fifo_in_valid
	wire  [63:0] avalon_st_adapter_008_out_0_data;          // avalon_st_adapter_008:out_0_data -> mac_0:tx_st_fifo_in_data
	wire         avalon_st_adapter_008_out_0_ready;         // mac_0:tx_st_fifo_in_ready -> avalon_st_adapter_008:out_0_ready
	wire         avalon_st_adapter_008_out_0_startofpacket; // avalon_st_adapter_008:out_0_startofpacket -> mac_0:tx_st_fifo_in_startofpacket
	wire         avalon_st_adapter_008_out_0_endofpacket;   // avalon_st_adapter_008:out_0_endofpacket -> mac_0:tx_st_fifo_in_endofpacket
	wire   [0:0] avalon_st_adapter_008_out_0_error;         // avalon_st_adapter_008:out_0_error -> mac_0:tx_st_fifo_in_error
	wire   [2:0] avalon_st_adapter_008_out_0_empty;         // avalon_st_adapter_008:out_0_empty -> mac_0:tx_st_fifo_in_empty
	wire         ethpack_transmitout1_valid;                // ethpack:transmitout_1_valid -> avalon_st_adapter_009:in_0_valid
	wire  [63:0] ethpack_transmitout1_data;                 // ethpack:transmitout_1_data -> avalon_st_adapter_009:in_0_data
	wire         ethpack_transmitout1_ready;                // avalon_st_adapter_009:in_0_ready -> ethpack:transmitout_1_ready
	wire         ethpack_transmitout1_startofpacket;        // ethpack:transmitout_1_sop -> avalon_st_adapter_009:in_0_startofpacket
	wire         ethpack_transmitout1_endofpacket;          // ethpack:transmitout_1_eop -> avalon_st_adapter_009:in_0_endofpacket
	wire         avalon_st_adapter_009_out_0_valid;         // avalon_st_adapter_009:out_0_valid -> mac_1:tx_st_fifo_in_valid
	wire  [63:0] avalon_st_adapter_009_out_0_data;          // avalon_st_adapter_009:out_0_data -> mac_1:tx_st_fifo_in_data
	wire         avalon_st_adapter_009_out_0_ready;         // mac_1:tx_st_fifo_in_ready -> avalon_st_adapter_009:out_0_ready
	wire         avalon_st_adapter_009_out_0_startofpacket; // avalon_st_adapter_009:out_0_startofpacket -> mac_1:tx_st_fifo_in_startofpacket
	wire         avalon_st_adapter_009_out_0_endofpacket;   // avalon_st_adapter_009:out_0_endofpacket -> mac_1:tx_st_fifo_in_endofpacket
	wire   [0:0] avalon_st_adapter_009_out_0_error;         // avalon_st_adapter_009:out_0_error -> mac_1:tx_st_fifo_in_error
	wire   [2:0] avalon_st_adapter_009_out_0_empty;         // avalon_st_adapter_009:out_0_empty -> mac_1:tx_st_fifo_in_empty
	wire         ethpack_transmitout2_valid;                // ethpack:transmitout_2_valid -> avalon_st_adapter_010:in_0_valid
	wire  [63:0] ethpack_transmitout2_data;                 // ethpack:transmitout_2_data -> avalon_st_adapter_010:in_0_data
	wire         ethpack_transmitout2_ready;                // avalon_st_adapter_010:in_0_ready -> ethpack:transmitout_2_ready
	wire         ethpack_transmitout2_startofpacket;        // ethpack:transmitout_2_sop -> avalon_st_adapter_010:in_0_startofpacket
	wire         ethpack_transmitout2_endofpacket;          // ethpack:transmitout_2_eop -> avalon_st_adapter_010:in_0_endofpacket
	wire         avalon_st_adapter_010_out_0_valid;         // avalon_st_adapter_010:out_0_valid -> mac_2:tx_st_fifo_in_valid
	wire  [63:0] avalon_st_adapter_010_out_0_data;          // avalon_st_adapter_010:out_0_data -> mac_2:tx_st_fifo_in_data
	wire         avalon_st_adapter_010_out_0_ready;         // mac_2:tx_st_fifo_in_ready -> avalon_st_adapter_010:out_0_ready
	wire         avalon_st_adapter_010_out_0_startofpacket; // avalon_st_adapter_010:out_0_startofpacket -> mac_2:tx_st_fifo_in_startofpacket
	wire         avalon_st_adapter_010_out_0_endofpacket;   // avalon_st_adapter_010:out_0_endofpacket -> mac_2:tx_st_fifo_in_endofpacket
	wire   [0:0] avalon_st_adapter_010_out_0_error;         // avalon_st_adapter_010:out_0_error -> mac_2:tx_st_fifo_in_error
	wire   [2:0] avalon_st_adapter_010_out_0_empty;         // avalon_st_adapter_010:out_0_empty -> mac_2:tx_st_fifo_in_empty
	wire         ethpack_transmitout3_valid;                // ethpack:transmitout_3_valid -> avalon_st_adapter_011:in_0_valid
	wire  [63:0] ethpack_transmitout3_data;                 // ethpack:transmitout_3_data -> avalon_st_adapter_011:in_0_data
	wire         ethpack_transmitout3_ready;                // avalon_st_adapter_011:in_0_ready -> ethpack:transmitout_3_ready
	wire         ethpack_transmitout3_startofpacket;        // ethpack:transmitout_3_sop -> avalon_st_adapter_011:in_0_startofpacket
	wire         ethpack_transmitout3_endofpacket;          // ethpack:transmitout_3_eop -> avalon_st_adapter_011:in_0_endofpacket
	wire         avalon_st_adapter_011_out_0_valid;         // avalon_st_adapter_011:out_0_valid -> mac_3:tx_st_fifo_in_valid
	wire  [63:0] avalon_st_adapter_011_out_0_data;          // avalon_st_adapter_011:out_0_data -> mac_3:tx_st_fifo_in_data
	wire         avalon_st_adapter_011_out_0_ready;         // mac_3:tx_st_fifo_in_ready -> avalon_st_adapter_011:out_0_ready
	wire         avalon_st_adapter_011_out_0_startofpacket; // avalon_st_adapter_011:out_0_startofpacket -> mac_3:tx_st_fifo_in_startofpacket
	wire         avalon_st_adapter_011_out_0_endofpacket;   // avalon_st_adapter_011:out_0_endofpacket -> mac_3:tx_st_fifo_in_endofpacket
	wire   [0:0] avalon_st_adapter_011_out_0_error;         // avalon_st_adapter_011:out_0_error -> mac_3:tx_st_fifo_in_error
	wire   [2:0] avalon_st_adapter_011_out_0_empty;         // avalon_st_adapter_011:out_0_empty -> mac_3:tx_st_fifo_in_empty
	wire         rst_controller_reset_out_reset;            // rst_controller:reset_out -> [avalon_st_adapter:in_rst_0_reset, avalon_st_adapter_001:in_rst_0_reset, avalon_st_adapter_002:in_rst_0_reset, avalon_st_adapter_003:in_rst_0_reset, avalon_st_adapter_004:in_rst_0_reset, avalon_st_adapter_005:in_rst_0_reset, avalon_st_adapter_006:in_rst_0_reset, avalon_st_adapter_007:in_rst_0_reset, avalon_st_adapter_008:in_rst_0_reset, avalon_st_adapter_009:in_rst_0_reset, avalon_st_adapter_010:in_rst_0_reset, avalon_st_adapter_011:in_rst_0_reset, eth_in_mux:reset_n, ethpack:reset]
	wire         rst_controller_001_reset_out_reset;        // rst_controller_001:reset_out -> [mac_0:rst_in_reset_reset, mac_1:rst_in_reset_reset, mac_2:rst_in_reset_reset, mac_3:rst_in_reset_reset]

	eth4to1_eth_in_mux eth_in_mux (
		.clk               (clk_312_out_clk_clk),                       //   clk.clk
		.reset_n           (~rst_controller_reset_out_reset),           // reset.reset_n
		.out_data          (eth_in_mux_out_data),                       //   out.data
		.out_valid         (eth_in_mux_out_valid),                      //      .valid
		.out_ready         (eth_in_mux_out_ready),                      //      .ready
		.out_startofpacket (eth_in_mux_out_startofpacket),              //      .startofpacket
		.out_endofpacket   (eth_in_mux_out_endofpacket),                //      .endofpacket
		.out_empty         (eth_in_mux_out_empty),                      //      .empty
		.out_channel       (eth_in_mux_out_channel),                    //      .channel
		.in0_data          (avalon_st_adapter_out_0_data),              //   in0.data
		.in0_valid         (avalon_st_adapter_out_0_valid),             //      .valid
		.in0_ready         (avalon_st_adapter_out_0_ready),             //      .ready
		.in0_startofpacket (avalon_st_adapter_out_0_startofpacket),     //      .startofpacket
		.in0_endofpacket   (avalon_st_adapter_out_0_endofpacket),       //      .endofpacket
		.in0_empty         (avalon_st_adapter_out_0_empty),             //      .empty
		.in0_channel       (avalon_st_adapter_out_0_channel),           //      .channel
		.in1_data          (avalon_st_adapter_001_out_0_data),          //   in1.data
		.in1_valid         (avalon_st_adapter_001_out_0_valid),         //      .valid
		.in1_ready         (avalon_st_adapter_001_out_0_ready),         //      .ready
		.in1_startofpacket (avalon_st_adapter_001_out_0_startofpacket), //      .startofpacket
		.in1_endofpacket   (avalon_st_adapter_001_out_0_endofpacket),   //      .endofpacket
		.in1_empty         (avalon_st_adapter_001_out_0_empty),         //      .empty
		.in1_channel       (avalon_st_adapter_001_out_0_channel),       //      .channel
		.in2_data          (avalon_st_adapter_002_out_0_data),          //   in2.data
		.in2_valid         (avalon_st_adapter_002_out_0_valid),         //      .valid
		.in2_ready         (avalon_st_adapter_002_out_0_ready),         //      .ready
		.in2_startofpacket (avalon_st_adapter_002_out_0_startofpacket), //      .startofpacket
		.in2_endofpacket   (avalon_st_adapter_002_out_0_endofpacket),   //      .endofpacket
		.in2_empty         (avalon_st_adapter_002_out_0_empty),         //      .empty
		.in2_channel       (avalon_st_adapter_002_out_0_channel),       //      .channel
		.in3_data          (avalon_st_adapter_003_out_0_data),          //   in3.data
		.in3_valid         (avalon_st_adapter_003_out_0_valid),         //      .valid
		.in3_ready         (avalon_st_adapter_003_out_0_ready),         //      .ready
		.in3_startofpacket (avalon_st_adapter_003_out_0_startofpacket), //      .startofpacket
		.in3_endofpacket   (avalon_st_adapter_003_out_0_endofpacket),   //      .endofpacket
		.in3_empty         (avalon_st_adapter_003_out_0_empty),         //      .empty
		.in3_channel       (avalon_st_adapter_003_out_0_channel)        //      .channel
	);

	pmem_group_wrap ethpack (
		.clock               (clk_312_out_clk_clk),                       //        clock.clk
		.reset               (rst_controller_reset_out_reset),            //        reset.reset
		.packetin_0_data     (avalon_st_adapter_004_out_0_data),          //    packetin0.data
		.packetin_0_sop      (avalon_st_adapter_004_out_0_startofpacket), //             .startofpacket
		.packetin_0_eop      (avalon_st_adapter_004_out_0_endofpacket),   //             .endofpacket
		.packetin_0_valid    (avalon_st_adapter_004_out_0_valid),         //             .valid
		.packetin_0_ready    (avalon_st_adapter_004_out_0_ready),         //             .ready
		.packetin_1_data     (avalon_st_adapter_005_out_0_data),          //    packetin1.data
		.packetin_1_sop      (avalon_st_adapter_005_out_0_startofpacket), //             .startofpacket
		.packetin_1_eop      (avalon_st_adapter_005_out_0_endofpacket),   //             .endofpacket
		.packetin_1_valid    (avalon_st_adapter_005_out_0_valid),         //             .valid
		.packetin_1_ready    (avalon_st_adapter_005_out_0_ready),         //             .ready
		.packetin_2_data     (avalon_st_adapter_006_out_0_data),          //    packetin2.data
		.packetin_2_sop      (avalon_st_adapter_006_out_0_startofpacket), //             .startofpacket
		.packetin_2_eop      (avalon_st_adapter_006_out_0_endofpacket),   //             .endofpacket
		.packetin_2_valid    (avalon_st_adapter_006_out_0_valid),         //             .valid
		.packetin_2_ready    (avalon_st_adapter_006_out_0_ready),         //             .ready
		.packetin_3_data     (avalon_st_adapter_007_out_0_data),          //    packetin3.data
		.packetin_3_sop      (avalon_st_adapter_007_out_0_startofpacket), //             .startofpacket
		.packetin_3_eop      (avalon_st_adapter_007_out_0_endofpacket),   //             .endofpacket
		.packetin_3_valid    (avalon_st_adapter_007_out_0_valid),         //             .valid
		.packetin_3_ready    (avalon_st_adapter_007_out_0_ready),         //             .ready
		.packetout_0_sop     (ethpack_packetout0_startofpacket),          //   packetout0.startofpacket
		.packetout_0_eop     (ethpack_packetout0_endofpacket),            //             .endofpacket
		.packetout_0_data    (ethpack_packetout0_data),                   //             .data
		.packetout_0_channel (ethpack_packetout0_channel),                //             .channel
		.packetout_0_valid   (ethpack_packetout0_valid),                  //             .valid
		.packetout_0_ready   (ethpack_packetout0_ready),                  //             .ready
		.packetout_1_sop     (ethpack_packetout1_startofpacket),          //   packetout1.startofpacket
		.packetout_1_eop     (ethpack_packetout1_endofpacket),            //             .endofpacket
		.packetout_1_data    (ethpack_packetout1_data),                   //             .data
		.packetout_1_channel (ethpack_packetout1_channel),                //             .channel
		.packetout_1_valid   (ethpack_packetout1_valid),                  //             .valid
		.packetout_1_ready   (ethpack_packetout1_ready),                  //             .ready
		.packetout_2_sop     (ethpack_packetout2_startofpacket),          //   packetout2.startofpacket
		.packetout_2_eop     (ethpack_packetout2_endofpacket),            //             .endofpacket
		.packetout_2_data    (ethpack_packetout2_data),                   //             .data
		.packetout_2_channel (ethpack_packetout2_channel),                //             .channel
		.packetout_2_valid   (ethpack_packetout2_valid),                  //             .valid
		.packetout_2_ready   (ethpack_packetout2_ready),                  //             .ready
		.packetout_3_sop     (ethpack_packetout3_startofpacket),          //   packetout3.startofpacket
		.packetout_3_eop     (ethpack_packetout3_endofpacket),            //             .endofpacket
		.packetout_3_data    (ethpack_packetout3_data),                   //             .data
		.packetout_3_channel (ethpack_packetout3_channel),                //             .channel
		.packetout_3_valid   (ethpack_packetout3_valid),                  //             .valid
		.packetout_3_ready   (ethpack_packetout3_ready),                  //             .ready
		.tagin_data          (ethpack_tagin_data),                        //        tagin.data
		.tagin_valid         (ethpack_tagin_valid),                       //             .valid
		.tagin_ready         (ethpack_tagin_ready),                       //             .ready
		.transmitout_0_data  (ethpack_transmitout0_data),                 // transmitout0.data
		.transmitout_0_valid (ethpack_transmitout0_valid),                //             .valid
		.transmitout_0_ready (ethpack_transmitout0_ready),                //             .ready
		.transmitout_0_sop   (ethpack_transmitout0_startofpacket),        //             .startofpacket
		.transmitout_0_eop   (ethpack_transmitout0_endofpacket),          //             .endofpacket
		.transmitout_1_data  (ethpack_transmitout1_data),                 // transmitout1.data
		.transmitout_1_valid (ethpack_transmitout1_valid),                //             .valid
		.transmitout_1_ready (ethpack_transmitout1_ready),                //             .ready
		.transmitout_1_sop   (ethpack_transmitout1_startofpacket),        //             .startofpacket
		.transmitout_1_eop   (ethpack_transmitout1_endofpacket),          //             .endofpacket
		.transmitout_2_data  (ethpack_transmitout2_data),                 // transmitout2.data
		.transmitout_2_valid (ethpack_transmitout2_valid),                //             .valid
		.transmitout_2_ready (ethpack_transmitout2_ready),                //             .ready
		.transmitout_2_sop   (ethpack_transmitout2_startofpacket),        //             .startofpacket
		.transmitout_2_eop   (ethpack_transmitout2_endofpacket),          //             .endofpacket
		.transmitout_3_data  (ethpack_transmitout3_data),                 // transmitout3.data
		.transmitout_3_valid (ethpack_transmitout3_valid),                //             .valid
		.transmitout_3_ready (ethpack_transmitout3_ready),                //             .ready
		.transmitout_3_sop   (ethpack_transmitout3_startofpacket),        //             .startofpacket
		.transmitout_3_eop   (ethpack_transmitout3_endofpacket)           //             .endofpacket
	);

	eth4to1_mac_0 mac_0 (
		.clk_156_in_clk_clk                     (clk_clk),                                   //                    clk_156_in_clk.clk
		.clk_312_in_clk_clk                     (clk_312_out_clk_clk),                       //                    clk_312_in_clk.clk
		.mac10g_avalon_st_pause_data            (),                                          //            mac10g_avalon_st_pause.data
		.mac10g_avalon_st_rxstatus_valid        (),                                          //         mac10g_avalon_st_rxstatus.valid
		.mac10g_avalon_st_rxstatus_data         (),                                          //                                  .data
		.mac10g_avalon_st_rxstatus_error        (),                                          //                                  .error
		.mac10g_avalon_st_txstatus_data         (),                                          //         mac10g_avalon_st_txstatus.data
		.mac10g_avalon_st_txstatus_valid        (),                                          //                                  .valid
		.mac10g_avalon_st_txstatus_error        (),                                          //                                  .error
		.mac10g_csr_address                     (),                                          //                        mac10g_csr.address
		.mac10g_csr_waitrequest                 (),                                          //                                  .waitrequest
		.mac10g_csr_read                        (),                                          //                                  .read
		.mac10g_csr_readdata                    (),                                          //                                  .readdata
		.mac10g_csr_write                       (),                                          //                                  .write
		.mac10g_csr_writedata                   (),                                          //                                  .writedata
		.mac10g_link_fault_status_xgmii_rx_data (),                                          // mac10g_link_fault_status_xgmii_rx.data
		.mac10g_xgmii_rx_data                   (xgmii_rx_data_0_data),                      //                   mac10g_xgmii_rx.data
		.mac10g_xgmii_tx_data                   (xgmii_tx_data_0_data),                      //                   mac10g_xgmii_tx.data
		.rst_in_reset_reset                     (rst_controller_001_reset_out_reset),        //                      rst_in_reset.reset
		.rx_st_fifo_out_data                    (mac_0_rx_st_fifo_out_data),                 //                    rx_st_fifo_out.data
		.rx_st_fifo_out_valid                   (mac_0_rx_st_fifo_out_valid),                //                                  .valid
		.rx_st_fifo_out_ready                   (mac_0_rx_st_fifo_out_ready),                //                                  .ready
		.rx_st_fifo_out_startofpacket           (mac_0_rx_st_fifo_out_startofpacket),        //                                  .startofpacket
		.rx_st_fifo_out_endofpacket             (mac_0_rx_st_fifo_out_endofpacket),          //                                  .endofpacket
		.rx_st_fifo_out_empty                   (mac_0_rx_st_fifo_out_empty),                //                                  .empty
		.rx_st_fifo_out_error                   (mac_0_rx_st_fifo_out_error),                //                                  .error
		.tx_st_fifo_in_data                     (avalon_st_adapter_008_out_0_data),          //                     tx_st_fifo_in.data
		.tx_st_fifo_in_valid                    (avalon_st_adapter_008_out_0_valid),         //                                  .valid
		.tx_st_fifo_in_ready                    (avalon_st_adapter_008_out_0_ready),         //                                  .ready
		.tx_st_fifo_in_startofpacket            (avalon_st_adapter_008_out_0_startofpacket), //                                  .startofpacket
		.tx_st_fifo_in_endofpacket              (avalon_st_adapter_008_out_0_endofpacket),   //                                  .endofpacket
		.tx_st_fifo_in_empty                    (avalon_st_adapter_008_out_0_empty),         //                                  .empty
		.tx_st_fifo_in_error                    (avalon_st_adapter_008_out_0_error)          //                                  .error
	);

	eth4to1_mac_1 mac_1 (
		.clk_156_in_clk_clk                     (clk_clk),                                   //                    clk_156_in_clk.clk
		.clk_312_in_clk_clk                     (clk_312_out_clk_clk),                       //                    clk_312_in_clk.clk
		.mac10g_avalon_st_pause_data            (),                                          //            mac10g_avalon_st_pause.data
		.mac10g_avalon_st_rxstatus_valid        (),                                          //         mac10g_avalon_st_rxstatus.valid
		.mac10g_avalon_st_rxstatus_data         (),                                          //                                  .data
		.mac10g_avalon_st_rxstatus_error        (),                                          //                                  .error
		.mac10g_avalon_st_txstatus_data         (),                                          //         mac10g_avalon_st_txstatus.data
		.mac10g_avalon_st_txstatus_valid        (),                                          //                                  .valid
		.mac10g_avalon_st_txstatus_error        (),                                          //                                  .error
		.mac10g_csr_address                     (),                                          //                        mac10g_csr.address
		.mac10g_csr_waitrequest                 (),                                          //                                  .waitrequest
		.mac10g_csr_read                        (),                                          //                                  .read
		.mac10g_csr_readdata                    (),                                          //                                  .readdata
		.mac10g_csr_write                       (),                                          //                                  .write
		.mac10g_csr_writedata                   (),                                          //                                  .writedata
		.mac10g_link_fault_status_xgmii_rx_data (),                                          // mac10g_link_fault_status_xgmii_rx.data
		.mac10g_xgmii_rx_data                   (xgmii_rx_data_1_data),                      //                   mac10g_xgmii_rx.data
		.mac10g_xgmii_tx_data                   (xgmii_tx_data_1_data),                      //                   mac10g_xgmii_tx.data
		.rst_in_reset_reset                     (rst_controller_001_reset_out_reset),        //                      rst_in_reset.reset
		.rx_st_fifo_out_data                    (mac_1_rx_st_fifo_out_data),                 //                    rx_st_fifo_out.data
		.rx_st_fifo_out_valid                   (mac_1_rx_st_fifo_out_valid),                //                                  .valid
		.rx_st_fifo_out_ready                   (mac_1_rx_st_fifo_out_ready),                //                                  .ready
		.rx_st_fifo_out_startofpacket           (mac_1_rx_st_fifo_out_startofpacket),        //                                  .startofpacket
		.rx_st_fifo_out_endofpacket             (mac_1_rx_st_fifo_out_endofpacket),          //                                  .endofpacket
		.rx_st_fifo_out_empty                   (mac_1_rx_st_fifo_out_empty),                //                                  .empty
		.rx_st_fifo_out_error                   (mac_1_rx_st_fifo_out_error),                //                                  .error
		.tx_st_fifo_in_data                     (avalon_st_adapter_009_out_0_data),          //                     tx_st_fifo_in.data
		.tx_st_fifo_in_valid                    (avalon_st_adapter_009_out_0_valid),         //                                  .valid
		.tx_st_fifo_in_ready                    (avalon_st_adapter_009_out_0_ready),         //                                  .ready
		.tx_st_fifo_in_startofpacket            (avalon_st_adapter_009_out_0_startofpacket), //                                  .startofpacket
		.tx_st_fifo_in_endofpacket              (avalon_st_adapter_009_out_0_endofpacket),   //                                  .endofpacket
		.tx_st_fifo_in_empty                    (avalon_st_adapter_009_out_0_empty),         //                                  .empty
		.tx_st_fifo_in_error                    (avalon_st_adapter_009_out_0_error)          //                                  .error
	);

	eth4to1_mac_2 mac_2 (
		.clk_156_in_clk_clk                     (clk_clk),                                   //                    clk_156_in_clk.clk
		.clk_312_in_clk_clk                     (clk_312_out_clk_clk),                       //                    clk_312_in_clk.clk
		.mac10g_avalon_st_pause_data            (),                                          //            mac10g_avalon_st_pause.data
		.mac10g_avalon_st_rxstatus_valid        (),                                          //         mac10g_avalon_st_rxstatus.valid
		.mac10g_avalon_st_rxstatus_data         (),                                          //                                  .data
		.mac10g_avalon_st_rxstatus_error        (),                                          //                                  .error
		.mac10g_avalon_st_txstatus_data         (),                                          //         mac10g_avalon_st_txstatus.data
		.mac10g_avalon_st_txstatus_valid        (),                                          //                                  .valid
		.mac10g_avalon_st_txstatus_error        (),                                          //                                  .error
		.mac10g_csr_address                     (),                                          //                        mac10g_csr.address
		.mac10g_csr_waitrequest                 (),                                          //                                  .waitrequest
		.mac10g_csr_read                        (),                                          //                                  .read
		.mac10g_csr_readdata                    (),                                          //                                  .readdata
		.mac10g_csr_write                       (),                                          //                                  .write
		.mac10g_csr_writedata                   (),                                          //                                  .writedata
		.mac10g_link_fault_status_xgmii_rx_data (),                                          // mac10g_link_fault_status_xgmii_rx.data
		.mac10g_xgmii_rx_data                   (xgmii_rx_data_2_data),                      //                   mac10g_xgmii_rx.data
		.mac10g_xgmii_tx_data                   (xgmii_tx_data_2_data),                      //                   mac10g_xgmii_tx.data
		.rst_in_reset_reset                     (rst_controller_001_reset_out_reset),        //                      rst_in_reset.reset
		.rx_st_fifo_out_data                    (mac_2_rx_st_fifo_out_data),                 //                    rx_st_fifo_out.data
		.rx_st_fifo_out_valid                   (mac_2_rx_st_fifo_out_valid),                //                                  .valid
		.rx_st_fifo_out_ready                   (mac_2_rx_st_fifo_out_ready),                //                                  .ready
		.rx_st_fifo_out_startofpacket           (mac_2_rx_st_fifo_out_startofpacket),        //                                  .startofpacket
		.rx_st_fifo_out_endofpacket             (mac_2_rx_st_fifo_out_endofpacket),          //                                  .endofpacket
		.rx_st_fifo_out_empty                   (mac_2_rx_st_fifo_out_empty),                //                                  .empty
		.rx_st_fifo_out_error                   (mac_2_rx_st_fifo_out_error),                //                                  .error
		.tx_st_fifo_in_data                     (avalon_st_adapter_010_out_0_data),          //                     tx_st_fifo_in.data
		.tx_st_fifo_in_valid                    (avalon_st_adapter_010_out_0_valid),         //                                  .valid
		.tx_st_fifo_in_ready                    (avalon_st_adapter_010_out_0_ready),         //                                  .ready
		.tx_st_fifo_in_startofpacket            (avalon_st_adapter_010_out_0_startofpacket), //                                  .startofpacket
		.tx_st_fifo_in_endofpacket              (avalon_st_adapter_010_out_0_endofpacket),   //                                  .endofpacket
		.tx_st_fifo_in_empty                    (avalon_st_adapter_010_out_0_empty),         //                                  .empty
		.tx_st_fifo_in_error                    (avalon_st_adapter_010_out_0_error)          //                                  .error
	);

	eth4to1_mac_3 mac_3 (
		.clk_156_in_clk_clk                     (clk_clk),                                   //                    clk_156_in_clk.clk
		.clk_312_in_clk_clk                     (clk_312_out_clk_clk),                       //                    clk_312_in_clk.clk
		.mac10g_avalon_st_pause_data            (),                                          //            mac10g_avalon_st_pause.data
		.mac10g_avalon_st_rxstatus_valid        (),                                          //         mac10g_avalon_st_rxstatus.valid
		.mac10g_avalon_st_rxstatus_data         (),                                          //                                  .data
		.mac10g_avalon_st_rxstatus_error        (),                                          //                                  .error
		.mac10g_avalon_st_txstatus_data         (),                                          //         mac10g_avalon_st_txstatus.data
		.mac10g_avalon_st_txstatus_valid        (),                                          //                                  .valid
		.mac10g_avalon_st_txstatus_error        (),                                          //                                  .error
		.mac10g_csr_address                     (),                                          //                        mac10g_csr.address
		.mac10g_csr_waitrequest                 (),                                          //                                  .waitrequest
		.mac10g_csr_read                        (),                                          //                                  .read
		.mac10g_csr_readdata                    (),                                          //                                  .readdata
		.mac10g_csr_write                       (),                                          //                                  .write
		.mac10g_csr_writedata                   (),                                          //                                  .writedata
		.mac10g_link_fault_status_xgmii_rx_data (),                                          // mac10g_link_fault_status_xgmii_rx.data
		.mac10g_xgmii_rx_data                   (xgmii_rx_data_3_data),                      //                   mac10g_xgmii_rx.data
		.mac10g_xgmii_tx_data                   (xgmii_tx_data_3_data),                      //                   mac10g_xgmii_tx.data
		.rst_in_reset_reset                     (rst_controller_001_reset_out_reset),        //                      rst_in_reset.reset
		.rx_st_fifo_out_data                    (mac_3_rx_st_fifo_out_data),                 //                    rx_st_fifo_out.data
		.rx_st_fifo_out_valid                   (mac_3_rx_st_fifo_out_valid),                //                                  .valid
		.rx_st_fifo_out_ready                   (mac_3_rx_st_fifo_out_ready),                //                                  .ready
		.rx_st_fifo_out_startofpacket           (mac_3_rx_st_fifo_out_startofpacket),        //                                  .startofpacket
		.rx_st_fifo_out_endofpacket             (mac_3_rx_st_fifo_out_endofpacket),          //                                  .endofpacket
		.rx_st_fifo_out_empty                   (mac_3_rx_st_fifo_out_empty),                //                                  .empty
		.rx_st_fifo_out_error                   (mac_3_rx_st_fifo_out_error),                //                                  .error
		.tx_st_fifo_in_data                     (avalon_st_adapter_011_out_0_data),          //                     tx_st_fifo_in.data
		.tx_st_fifo_in_valid                    (avalon_st_adapter_011_out_0_valid),         //                                  .valid
		.tx_st_fifo_in_ready                    (avalon_st_adapter_011_out_0_ready),         //                                  .ready
		.tx_st_fifo_in_startofpacket            (avalon_st_adapter_011_out_0_startofpacket), //                                  .startofpacket
		.tx_st_fifo_in_endofpacket              (avalon_st_adapter_011_out_0_endofpacket),   //                                  .endofpacket
		.tx_st_fifo_in_empty                    (avalon_st_adapter_011_out_0_empty),         //                                  .empty
		.tx_st_fifo_in_error                    (avalon_st_adapter_011_out_0_error)          //                                  .error
	);

	eth4to1_pll_0 pll_0 (
		.refclk   (clk_clk),             //  refclk.clk
		.rst      (~reset_reset_n),      //   reset.reset
		.outclk_0 (clk_312_out_clk_clk), // outclk0.clk
		.locked   ()                     // (terminated)
	);

	eth4to1_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (64),
		.inChannelWidth  (6),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (64),
		.outChannelWidth (6),
		.outErrorWidth   (0),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (clk_312_out_clk_clk),                   // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),        // in_rst_0.reset
		.in_0_data           (ethpack_packetout0_data),               //     in_0.data
		.in_0_valid          (ethpack_packetout0_valid),              //         .valid
		.in_0_ready          (ethpack_packetout0_ready),              //         .ready
		.in_0_startofpacket  (ethpack_packetout0_startofpacket),      //         .startofpacket
		.in_0_endofpacket    (ethpack_packetout0_endofpacket),        //         .endofpacket
		.in_0_channel        (ethpack_packetout0_channel),            //         .channel
		.out_0_data          (avalon_st_adapter_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_out_0_empty),         //         .empty
		.out_0_channel       (avalon_st_adapter_out_0_channel)        //         .channel
	);

	eth4to1_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (64),
		.inChannelWidth  (6),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (64),
		.outChannelWidth (6),
		.outErrorWidth   (0),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_001 (
		.in_clk_0_clk        (clk_312_out_clk_clk),                       // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),            // in_rst_0.reset
		.in_0_data           (ethpack_packetout1_data),                   //     in_0.data
		.in_0_valid          (ethpack_packetout1_valid),                  //         .valid
		.in_0_ready          (ethpack_packetout1_ready),                  //         .ready
		.in_0_startofpacket  (ethpack_packetout1_startofpacket),          //         .startofpacket
		.in_0_endofpacket    (ethpack_packetout1_endofpacket),            //         .endofpacket
		.in_0_channel        (ethpack_packetout1_channel),                //         .channel
		.out_0_data          (avalon_st_adapter_001_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_001_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_001_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_001_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_001_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_001_out_0_empty),         //         .empty
		.out_0_channel       (avalon_st_adapter_001_out_0_channel)        //         .channel
	);

	eth4to1_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (64),
		.inChannelWidth  (6),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (64),
		.outChannelWidth (6),
		.outErrorWidth   (0),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_002 (
		.in_clk_0_clk        (clk_312_out_clk_clk),                       // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),            // in_rst_0.reset
		.in_0_data           (ethpack_packetout2_data),                   //     in_0.data
		.in_0_valid          (ethpack_packetout2_valid),                  //         .valid
		.in_0_ready          (ethpack_packetout2_ready),                  //         .ready
		.in_0_startofpacket  (ethpack_packetout2_startofpacket),          //         .startofpacket
		.in_0_endofpacket    (ethpack_packetout2_endofpacket),            //         .endofpacket
		.in_0_channel        (ethpack_packetout2_channel),                //         .channel
		.out_0_data          (avalon_st_adapter_002_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_002_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_002_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_002_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_002_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_002_out_0_empty),         //         .empty
		.out_0_channel       (avalon_st_adapter_002_out_0_channel)        //         .channel
	);

	eth4to1_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (64),
		.inChannelWidth  (6),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (64),
		.outChannelWidth (6),
		.outErrorWidth   (0),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_003 (
		.in_clk_0_clk        (clk_312_out_clk_clk),                       // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),            // in_rst_0.reset
		.in_0_data           (ethpack_packetout3_data),                   //     in_0.data
		.in_0_valid          (ethpack_packetout3_valid),                  //         .valid
		.in_0_ready          (ethpack_packetout3_ready),                  //         .ready
		.in_0_startofpacket  (ethpack_packetout3_startofpacket),          //         .startofpacket
		.in_0_endofpacket    (ethpack_packetout3_endofpacket),            //         .endofpacket
		.in_0_channel        (ethpack_packetout3_channel),                //         .channel
		.out_0_data          (avalon_st_adapter_003_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_003_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_003_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_003_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_003_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_003_out_0_empty),         //         .empty
		.out_0_channel       (avalon_st_adapter_003_out_0_channel)        //         .channel
	);

	eth4to1_avalon_st_adapter_004 #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (64),
		.inChannelWidth  (0),
		.inErrorWidth    (6),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (64),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_004 (
		.in_clk_0_clk        (clk_312_out_clk_clk),                       // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),            // in_rst_0.reset
		.in_0_data           (mac_0_rx_st_fifo_out_data),                 //     in_0.data
		.in_0_valid          (mac_0_rx_st_fifo_out_valid),                //         .valid
		.in_0_ready          (mac_0_rx_st_fifo_out_ready),                //         .ready
		.in_0_startofpacket  (mac_0_rx_st_fifo_out_startofpacket),        //         .startofpacket
		.in_0_endofpacket    (mac_0_rx_st_fifo_out_endofpacket),          //         .endofpacket
		.in_0_empty          (mac_0_rx_st_fifo_out_empty),                //         .empty
		.in_0_error          (mac_0_rx_st_fifo_out_error),                //         .error
		.out_0_data          (avalon_st_adapter_004_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_004_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_004_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_004_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_004_out_0_endofpacket)    //         .endofpacket
	);

	eth4to1_avalon_st_adapter_004 #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (64),
		.inChannelWidth  (0),
		.inErrorWidth    (6),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (64),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_005 (
		.in_clk_0_clk        (clk_312_out_clk_clk),                       // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),            // in_rst_0.reset
		.in_0_data           (mac_1_rx_st_fifo_out_data),                 //     in_0.data
		.in_0_valid          (mac_1_rx_st_fifo_out_valid),                //         .valid
		.in_0_ready          (mac_1_rx_st_fifo_out_ready),                //         .ready
		.in_0_startofpacket  (mac_1_rx_st_fifo_out_startofpacket),        //         .startofpacket
		.in_0_endofpacket    (mac_1_rx_st_fifo_out_endofpacket),          //         .endofpacket
		.in_0_empty          (mac_1_rx_st_fifo_out_empty),                //         .empty
		.in_0_error          (mac_1_rx_st_fifo_out_error),                //         .error
		.out_0_data          (avalon_st_adapter_005_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_005_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_005_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_005_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_005_out_0_endofpacket)    //         .endofpacket
	);

	eth4to1_avalon_st_adapter_004 #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (64),
		.inChannelWidth  (0),
		.inErrorWidth    (6),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (64),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_006 (
		.in_clk_0_clk        (clk_312_out_clk_clk),                       // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),            // in_rst_0.reset
		.in_0_data           (mac_2_rx_st_fifo_out_data),                 //     in_0.data
		.in_0_valid          (mac_2_rx_st_fifo_out_valid),                //         .valid
		.in_0_ready          (mac_2_rx_st_fifo_out_ready),                //         .ready
		.in_0_startofpacket  (mac_2_rx_st_fifo_out_startofpacket),        //         .startofpacket
		.in_0_endofpacket    (mac_2_rx_st_fifo_out_endofpacket),          //         .endofpacket
		.in_0_empty          (mac_2_rx_st_fifo_out_empty),                //         .empty
		.in_0_error          (mac_2_rx_st_fifo_out_error),                //         .error
		.out_0_data          (avalon_st_adapter_006_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_006_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_006_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_006_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_006_out_0_endofpacket)    //         .endofpacket
	);

	eth4to1_avalon_st_adapter_004 #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (64),
		.inChannelWidth  (0),
		.inErrorWidth    (6),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (64),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_007 (
		.in_clk_0_clk        (clk_312_out_clk_clk),                       // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),            // in_rst_0.reset
		.in_0_data           (mac_3_rx_st_fifo_out_data),                 //     in_0.data
		.in_0_valid          (mac_3_rx_st_fifo_out_valid),                //         .valid
		.in_0_ready          (mac_3_rx_st_fifo_out_ready),                //         .ready
		.in_0_startofpacket  (mac_3_rx_st_fifo_out_startofpacket),        //         .startofpacket
		.in_0_endofpacket    (mac_3_rx_st_fifo_out_endofpacket),          //         .endofpacket
		.in_0_empty          (mac_3_rx_st_fifo_out_empty),                //         .empty
		.in_0_error          (mac_3_rx_st_fifo_out_error),                //         .error
		.out_0_data          (avalon_st_adapter_007_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_007_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_007_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_007_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_007_out_0_endofpacket)    //         .endofpacket
	);

	eth4to1_avalon_st_adapter_008 #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (64),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (64),
		.outChannelWidth (0),
		.outErrorWidth   (1),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_008 (
		.in_clk_0_clk        (clk_312_out_clk_clk),                       // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),            // in_rst_0.reset
		.in_0_data           (ethpack_transmitout0_data),                 //     in_0.data
		.in_0_valid          (ethpack_transmitout0_valid),                //         .valid
		.in_0_ready          (ethpack_transmitout0_ready),                //         .ready
		.in_0_startofpacket  (ethpack_transmitout0_startofpacket),        //         .startofpacket
		.in_0_endofpacket    (ethpack_transmitout0_endofpacket),          //         .endofpacket
		.out_0_data          (avalon_st_adapter_008_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_008_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_008_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_008_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_008_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_008_out_0_empty),         //         .empty
		.out_0_error         (avalon_st_adapter_008_out_0_error)          //         .error
	);

	eth4to1_avalon_st_adapter_008 #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (64),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (64),
		.outChannelWidth (0),
		.outErrorWidth   (1),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_009 (
		.in_clk_0_clk        (clk_312_out_clk_clk),                       // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),            // in_rst_0.reset
		.in_0_data           (ethpack_transmitout1_data),                 //     in_0.data
		.in_0_valid          (ethpack_transmitout1_valid),                //         .valid
		.in_0_ready          (ethpack_transmitout1_ready),                //         .ready
		.in_0_startofpacket  (ethpack_transmitout1_startofpacket),        //         .startofpacket
		.in_0_endofpacket    (ethpack_transmitout1_endofpacket),          //         .endofpacket
		.out_0_data          (avalon_st_adapter_009_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_009_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_009_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_009_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_009_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_009_out_0_empty),         //         .empty
		.out_0_error         (avalon_st_adapter_009_out_0_error)          //         .error
	);

	eth4to1_avalon_st_adapter_008 #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (64),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (64),
		.outChannelWidth (0),
		.outErrorWidth   (1),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_010 (
		.in_clk_0_clk        (clk_312_out_clk_clk),                       // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),            // in_rst_0.reset
		.in_0_data           (ethpack_transmitout2_data),                 //     in_0.data
		.in_0_valid          (ethpack_transmitout2_valid),                //         .valid
		.in_0_ready          (ethpack_transmitout2_ready),                //         .ready
		.in_0_startofpacket  (ethpack_transmitout2_startofpacket),        //         .startofpacket
		.in_0_endofpacket    (ethpack_transmitout2_endofpacket),          //         .endofpacket
		.out_0_data          (avalon_st_adapter_010_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_010_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_010_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_010_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_010_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_010_out_0_empty),         //         .empty
		.out_0_error         (avalon_st_adapter_010_out_0_error)          //         .error
	);

	eth4to1_avalon_st_adapter_008 #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (64),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (64),
		.outChannelWidth (0),
		.outErrorWidth   (1),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_011 (
		.in_clk_0_clk        (clk_312_out_clk_clk),                       // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),            // in_rst_0.reset
		.in_0_data           (ethpack_transmitout3_data),                 //     in_0.data
		.in_0_valid          (ethpack_transmitout3_valid),                //         .valid
		.in_0_ready          (ethpack_transmitout3_ready),                //         .ready
		.in_0_startofpacket  (ethpack_transmitout3_startofpacket),        //         .startofpacket
		.in_0_endofpacket    (ethpack_transmitout3_endofpacket),          //         .endofpacket
		.out_0_data          (avalon_st_adapter_011_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_011_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_011_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_011_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_011_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_011_out_0_empty),         //         .empty
		.out_0_error         (avalon_st_adapter_011_out_0_error)          //         .error
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_312_out_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
