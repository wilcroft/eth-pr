// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:08 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FXl1F2YG4/qe8BMT6bMzDmKGNMb7oOOroJqGY7heK+vnvhWL7YSIYGf5QAU9i1Lc
1DTB4ek3EBJXs3ov9/KWVhDxvlvdPDxySOx456XS6L6Uo84awqnJjZzAmfyQJqyF
G3Kra7x2K2kYmXeZ1leupSg5CZw/bQLhQmES2Cfjgzw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13344)
jMb3czLOouEH2z1bkz9KhRlZMTTFJM9ml53xw9a8fiLab34WyLtGhKknQ4in1xxA
ywH19shtrKdwwrUpLf+5R2JMQygS6slHz/0shbwdH0XTr4GUbqGFhYOk7SB2hDeo
7AAO8c7DJapi1Gw3KT8KeHOtAGh5k/Y3X8WBLFMv1mSnL0UdKZ/mSpsq2ZjpmU3L
ANhFBtAfScvJcZUcXdPxBCAnS/eWwXVoAJNBJUQjnx/zJuOQ9DYR3kVm2z28iatK
IdITxwxelWYS5Y8sN1tlKomwuV6SENkcIPkweMNEEHt2BG0mdp3m/SORqLC1aRWL
nc4+Mb4g9Q3JYyLEZA7XPPgIFZ0JGY/4WrBfpqUfPOh7jgmXN/KfSqLBEgmT5YEz
dt2AT5pxhw62nWudbAC/KHN2AGRgg4kzQ6mVTdi72E/91rdNFiKtk2gkKRL8s/xU
eF0gkNBoC2c7WVFljap+SRSDRtYl6/Gt9vPjnKDYaiiYq08OjPBpoal7wAGE2MLV
oCNzzZa2Qg+OvVH/2iGhR+Vl/aeN6Z9f5BRrwUlMpScoa43Imbg6k9pM10Wr3cbs
GNC2sTqX1ICGKfUu2MSfY9u0tGbf6JNkYgRFnltOY+CWVbCF13oMeqhIsBLPLhXE
1cKcfYOk92QCkfrMlPPnpYKK3M4K4WzZO97vT4/sWgtcKWBoEFe3dJ32Xcsmcecn
eEZHJTIivavnRLAngbkbnlIhdraRm+1cLpakCw4vazXjbxJA7nahKaA6Sm4kZ/Fi
0/kONX/NHuohAfwVCsBxIY4VYMTOO6ipLzRqLq646zEf/yjHtQDEIz2OjaX/anbd
fQ0vs9y51jvM01WcLpD95u5S13ck0QDolbgonbdkf50PCDuU1u3Eg7IObQCVCCrY
q1iNeW2GOMjU0MKtDzRFmaCh2dV/XFlobAdddwxOsIhQbyD98PHTzomEhXh0KpQN
zREJzSwDqBEEBahwzzOTKsok4L8Hlp+Nbwz+swrP/1/BiB9f7bRXQ2iMSrVF9B2J
rjomxZYTj6UyJ5Uxbe8xgKopgnxjvJ8tL1LLG2ucTi4EkFIuCczCv51xgBDp964J
jhDFeFCFQiKPRiND31jbEN5q6b95ELqUA/FxsYAFz+danC2zxBkUvzIN1iKVLW0z
dJ6SD8l6Jim3n5up6Ep1MOuRoGN6NUCyfg9lC8qia1hrK/XM3a/QdORJz66TXkSl
ACXSnwlpJCyX+1Z79LjAFPi4eSUJ4wB19wuVurnNSbgEzuEwY5K2GgUkVYwJCfs3
M7qCaFEsZwXxax1H/OIawGEiTHGqprcCV/nbVBq7U2CVTNjlL1oFFgRSqL9bUmRy
kd6dooBYoXiRdcKjZxwJRqZm/5/tswGZ/ij9oDKA/ICThetjF8put6YMX9QQydU1
q4dPuimnO/hMZqNZiX2DZ/wsqyzwHU7vqbWZmnPWeMRJUxzqhK19q5v6cwPkfyF/
ICERwmJxAChxhueKwc29qMmkjoNvDOWLFhjBrOKOSW4Qu7jUIcbxum0K6viV7mXY
Zj89fkVhppFJZqNJbwdRQ0wnDtfHU5EZWgKyfOYjK5h0ARdUasbDmBhriadspkGe
xFXPg2QVhvvAZozUt2Vy9euQloUnJAnmhcRSMGkCPDgA2aDcJnj/RsCHGDB28Oqi
NOjnj03B5h1LGRz8URrDrkftZQ3acmYErIODCw+TzwE2sR4Qb+dYitohxlJ2GjNc
K/iXU3W6wSryzq3H0IT8MfH/hAjhfiT5dGZne+OSfzBzkI4dSugzVSh39aGOZOeq
H5ypzE9Cc3pTHZCfm4mpUXwuoCo89hwy9BSBV91/lBwOyp4zLp6oJdXOwgJXa0VQ
8W3Vd93VUEcp5BuQNhOEgEcGQadHWvw1VPbVvsmbEnkmSSc7s+NIN2fJBIJS+HkR
AlUwrG9wWpKqAdV50f/1t3NV3WDmHo3CEsVqv/ZqIglbuyHlfgliwMqK3/uUEKZ4
WL6l7iyWJ+HoysZxGrtBdnJgrMMxvxVaKuY5ZlUJayde+d9FgtbWJIeA6af3cN3+
pYZXGqIlgE40rc+fcjedFXTM+srTqm9S/bIqSZhdW9xctucyqBfd0xLFtphRUJpc
25WahQsXTHLq6F3gzXk1ac4BhLDaZQIRYSPssNTrRw1Y5WRTkJ4eWBXc/YTRfRbU
RxaANH+//i2jNJxDsBGi9nTo8X5jahub/srzmsws5bTe9/L2qYysRbXJnAyKpX9s
ySfFNXJeNmOT+V3JL3RrIumnC6yl2/mchkEkCdDiu+p27uACULp3LuWTdKt9DPHT
3HDjEzOux8awt58P08Ffa+gsnJz9U86feeEPE/x4bdVeTFvmHqTbG2vNUj5So1UD
Z1yozIOXN23P/JZ+wnbHsSNbyMnPsYVOGmWSZLfCH2qn0Gd49EK/CiRV68CqmQTN
OnlQ+ZdUi9eOdxiS64/StEOH3fUD3jzD88KdqcEdxSNyvW+QYSgZFlifb61aj3Ih
BDLWZJe+8GLkLMWPjVdg33SFx87B4EBNU0FX1My/CcHNfU9XfwRyNAsOdj6aUXNq
izRGUuxnoVEecfjdW6z7wT7kWD+TvHbqto+v0ka381hHmCisH0GebrPo8k3U3CWt
1kkawoGW8Jitnh8QKh+z4lG+6bGEcCzqO0sJ+kQh5kguUN1Y92p1+vpy3P1CFi1h
J8tAqHbceTMv4jLPbZ5QHwZf8kbxlA4Lj/95jNviHnu5ISGp74stnMYD5N/Tt5uw
VzeeEZ8115OCK/0uL9KaL4ele06/uBo4KTSn30BAdm0kRWAtgB2pR2aOGoreOIJ+
BXWNmHClf1MxJ9VQ6zhtKN51x55Gb8TKxALomzexM9ISp7mxXG2bmZ5cO0BL9t1p
xGSho5VBvbMTPbmps2ieUIpQ2+/w2bjL19mDtfkxTQPyw4enF6ixkBPqjuqmxG0g
LzayqIHVjE+Os9IEGQq+mOb4ghUKZe+FnOB5hgZgfARC4G/zIkl1MkGLe4Of7Iu8
Ew5mp6LCe88oXid0QlNi5uo7ERgGtwYBljc0ER78e9Q1gGdCoAo06XAhEy0phsy0
UCn0GoUsyYxY/Az1pKLGtvtuysUd7rLDdwXM730XU6edV5kpu6/IbgEmh2Vistvh
jSkUj40gEvWwtGL/qoXKi/pFe5XpSAU6OOV0kLhGbfSB30VbX/1HabiVx3934Yqo
0lQ9OlVZsZSWfowM+xTLipAAT1hcylGT2uhxwKpU0KmlgVXKhhyKYmNpsB/tlzYT
mhDLyQ1hP5HSnqqj5or6S+vlBKvVJAMr4MbAkxHN0XDolFvVkxZBARaacCoHu6KU
+Da6lYqcGeXuTdXZMozKXW3f0eW3Jptx8Xr62ekhGJhchOAnLjTvr8xf3b+ZmTiv
WpgX6EyCCzNJ8pNTylrk27EPOtvMEGw9va/12apaOmC0YQhTOc86k8b7rx3sGzr9
stAU+QTExX6RcZRRXbRAoHqsHyr+/XhFJJBaM6d7sNKy7SMi6IT9qUtPGjUXd61P
vFZtyHIaIbCsebHnujailZmXUUykQRAX983V43TzaorlOc3n669Mj3WoJbXY8RTy
EuR4WS8p+lOHs3iIdsZq/fNWPqSMlJdzdqVGi9+lOklOApx/MrDt82sg8h12vXry
XonaS9Ashm1sMeDecJpApIszfpihcWUEG2CjCrSwMoH9Fb6QPte1u00YgnbupCCx
VZ3uBjl1dwO2BYZ0VA5gMaU15rmKMMgh/C1gZnWhusc4qFU2sXVyZk4OilvnwKiH
IJ7PDSoD4CJHQez6pAaxEh3RBsRZz3lrxbVspo8WfWBi4KcCUVRDGQKp9KUnirdI
Q2GsFFAnb6wngjoqR9NIz8Ejzh/3bGgiRUM8+G7+hZwPePvhQNcC+OI0vLFZXhjr
WZDseDYlPcBK5ZVxfJ0Y1VAZDy5QXVohfN4RWXXkdnIOFfRTiLMQO5XhL+QatiUm
K+7FVXP5iQRPYloIjgTQ8I0aBqpgOV6tvEBsaoQLtIjVnOWZE9zC2XZ04YS7wiAu
FwoL/cvId9r7CsHd/somvzTDDFPdcF/sPNKyenjY2YE5TMh7Jcj3bZLwnlJ9uSn7
25DJIgjOOu4Y0RySRztRw0ILzOSG69PWeJP7mzLyGMk1bhO43f/S4RFWYpwvsaSZ
O4rS2W5D9rx7Q9zyj9OhnzSt6VbVq6ZsXk1I21J9kYtQpIn3XgOfp8a0SPD2YKHP
5IVnSi04Jy1EOY58rlrP6ZeEXg2rFJFgeTDDc2AWS24/0czbMz9VQrGgwl2y2nHP
/AGfOaso2/nbphexU5EkNiqXTRlvXR3ctCqjDcKC6OY15HcXM9vwiF3NuhIYV9JT
DE9mOw+UsdMIvPZuEK774WPLBezt2cm+ijhYZ8rQj5cvVxt2akCuTrWpbWx64CoA
YdCpIdhO/YY8g/y6GT0dGgDczP57a5UZqevF4GC7ru5qXHye2O1jo3qpgMilYw/t
xONeyUTyufoBD8iGZB72L7YQ8aaNR7DGoj6Cfa0vgaDPsXkZcSonIrLV6GbVNqgQ
TsyWRodxpCN/qHhdMdxVjPNslO9FT3nm71nqNPtTd03hdF8vqlU1ngkfVlFK+cou
CZDrfqfXHlirnqCIRgSynRYZ/vaW0bwNFsL83LebYHXqy/iPrrItdYxBdDSpyhcT
+v/uaR1xUNvh8fiyuuaN+9U+gbdvwI/xrzDwzRriFnUhiJuRDIER08K9QQO2CmWl
Cg+k1ishv3ciTMebZ2e1tO3uzu4wRFMdlDHUvRYvLHUacn0fWPzR9hpHwxURaZup
zbQEaKTAhS6YfJ2ypozE1KTuWya/Zl44iW1Ng2NQmAvfFWJ5sNVW4zvU8LItvRsq
Iv0/SYQtzApk+NinendtKkg6C4ggVwvQ9RHf11Qjg9Ruzs0rsdVU2HWH5GdiKy58
pbUqYjGIz2c1mp4IcELcEKMb3ffgNQdHBrJ7IPGRYlffNOQFjV+sf1AfWS8+6Mp/
uxL/Rp9R476aem8JbhRPwFQlaT+UgZY8shJrYaD+uN+N4UASQaXN3EP/pWmem5dk
4Pr72rlbw3/Z2d7V/BilpAx+QZSbS6mrrWRBzWl48x+LiOxK5/KBum2ae3hGrJbH
8ahORGxhWy02XioRRhoVdUqlwtJsBWAEjM7o5pd+1aPkmmdtfiA81+BwkFLHLsK9
2E3Is2+3XVWa7r13TKILJn5YGKSBia+/DIAJ9rlHhsvT29KX99+Rs5ByJef0iWgQ
fhgQ6TmMRm4jPk/tSDdRAlKoXyHF3IRwe3Tj15klVXQ4WMqMzOt8N4fA4wOFUkX8
IY7fW+Nm3xU8RRacKunvPlGNN7gPQRFG/F3RdLYJiM2fMLsMRd0OW0GrWDnuLbqH
sXj8FSoEiP3lPZ8ClBd2j9twc+H6fSfwcZkcHgF5EAfnZwMwCynO8wXzcyXyiTxI
xpjQlsfOJgcnTCrQeD9WhytzoE8DyfU1fOuH1kImAseECZGPtewj41Rb7zzQSVh4
oxIFh7igVePCv3E5USDHaLCYKKJ3af/ygsziY22Mj32X+b+cy6GSWkpnpRwIrHSd
ahuBp76Lc73aml0nkDbR3eA+8PtIMB1CF1FLY+M4ZhrOoqMcKhALagfZibO/UVVC
tZejk0btrnseTjfXfSnax0Pi3Igxcfxt0OGKczlKpmfDkE9/J2HuvzTZZMstGuRK
tmrQZGhyKxcv81dRhBVe1RExXIy9HC3BMab0UmlFmj3stEEvJsTnS/CTZVwCkLAb
Zun3SEbT+U9ecrQLZLn+N+sTI1TXdfvi4rxP2UMXUjT1dVdrKesjfmi6aC/g00ZA
vGmdLa6rYnJKowIpyjHRYVAAXnnKCxdsfhK9beqbXEnSWYfbOnUzUeukAzgYglwk
MhdY3iKtq8GU9hAohxq1V5WNeZS/LEVwGIY0vtekPYCTSj2X27SIvrIJCv1G2Whg
K6iWLXYpKlt6hgNVvhpuQgaMWaecnWfza3Gm8ZedhV2YDvopV9A7MTsrkoZn1PMy
PACUxJIlg1OlrbGIDJr1PEgrGOZPAxb5ziq1SIxmOuyGdINi/ljGMRjl454/JlT5
9u/9GkuTNnlfM/MvO9uNQrpn85jJmsDbI64fNfU32nLB+RoxPI4PRgHwuSNc8TpC
yJDslMJrm4PI5e0QViM1AddkHxISbRlgZoFk67vVbTXyU3ht9Yk9NngS4RaW8C8e
uEB+65e9lkz/YsdAPrc5G3u8NHHAZ0g4qxlhDFZf128s0ROtBjHyUuPCK7/fNbyR
PXd5B2zi6kFXHV4KL9sLuPxk0X9uX1b4K4pLs3FfSNvpe2qwurrWClnnpHs18+tt
c+lZ/TJIXjN+8X0oDhiUcw+YGzT+ZlsLUs+lWVaiOFTM40n8zdz1bHKw5ZnuIFyF
HjcMtKHw5++YiB7m0OaP/OxmPTsmWdSnwvjJt0lR4+q9UD2aHF8C11MU1LoCCaOu
Di49OuhjPcyiVcN+k9A3vDyG/qPN8cBub0tSnvtx+7440u8g88GYfxUhKgocRVHs
ntiSQQkBLgteBUdh+gYg7IuiTTitqu0a0ixOGQDrogfsffBCteP5kbO+G5ESrjOq
Y1C+kIh98K+zjSothoj+89MMSI5eRHpobBz/2IbOCKkIH4uGoa7G3hj/VucRfPwY
8LrartiNcPRYCCN0YvRBrB6ZTgFB6x+gzkUZhX2o6FCscQGI0Kg1bPfxW+/8cPmr
Rnr6suvaMbAXHITe/vEh3hpEy3rYqsDfVNBqUS2pj+DZkEuBx3dOSiQ8rygamChq
RZcSRMdozK3fqt41RN3Nu2M7SFWUnTiCuyssbbmCzdU/GLIR8XrU2wHwtG1MNI0s
7+rdk9T6zgbDiiLMukw8KIDDEh9cWrigjMgVR3SfRvZNCovAmxlRW73dF6BNl42w
YkzPOsktrClISprs3G3C8b3oohGD6zKjK10A33y4TJ1H2uCDSVp5sTDBZEGEYY+c
hAESWHsIUa+Ry1gFLPJQD5Nc7KxnI6KYpKkVY62v6udvqnMWU/1C43w5JSiPDMct
U88slQvJg37lYKKtcnxdQK6YvEjQpf7ISu0leB61UdWO9XtmN+V6DdLoBa8Ihlqg
9pOiriOw61iBHedDFRkPv7GeurW4WvaUvljgmPxJrvRhc+8JdBKGYmZWvJwDjF5z
P44qQxddjuviB9pLlJiQbLXyjacxbw/uIW4wQq+n7QxEisBzAxJDAvbsrOJe9DSf
dCaj0Z9bevEclLY3bDxuNWe5HFCzeSoZCogBz2rV725CvcR0uoFD972ZYiyssfTp
gVJspG4cgl+PR1yckhdAVSRNg+C/m/4FiyY19A3wPJjsID2kmsO4e+YbXElBW0pr
m0jShTjrUn1/QA6nG8IpYawiH+lPdNaJCVY5EiWkli22HzOyK7La0CTbBXzpW+Ij
rZYHXaeiJAuwb+UUkvgcteSfKEYRig1JqKIyUVcdQdg4pb0piku5GokyTd9hPLUw
K1YjGNavarjVKeMNWci66+uqmWLGkASR0iKeHXFlDJdybAcEi2QoROwLWLL88dJm
5z8pK/W/i+wPMhLika1owzP4epYs9mYXCr70BtxzBE+EYuO4PskLGchbbPwe1VTS
ZFKgMSq8VF1F1CQkxxb07r9j2INsuE+r95RX9DHi8QRiaRGxkl693hn28ENrh8uZ
QajO5PDFbRrs5KBqoIIOD/Rv1dS5wb9UvCnVJDycd13HvloWt3NRecEa+ZHPM0u7
RaYG/5luN4DUb4dSHZ8asGS12Bp5rAnLtr4fYlRunXY/t9grbeijNM9cKYiEEW21
JaUefxq9byxcZXggHzGQzAxHkW3w9xIE0JU+AFxxPjNvJ57s9TTa6HgwHIZ1fhOw
KvqrXmFPneaQQMwOCzXo2DY89/LLiIh7lKToloPjs8zr0rm/9eqAoTN3LB2DWzuo
qUXONrlGvr8y33sf6/WTWgQXeXr9Ju0JZOc8K6Jrme59N8plRS+oXsULHhe+81Q3
RoW4uO3NUnUrGj987dGKZBuvmZDMs9tJY1EvNvBUoV0eH4sNByLKAUwpL+fWXQxd
8uE36D+nrsbP8fnW5mc1yGlWFqfYF6wVT8HL6xBNdyU1zpb+afsJg5CPiCDIR1Bt
G5jAo/G31IfEbzBkJnayLNhMeTKTGLx0K3eWlfjDKLG9d/3Vsvx9sn9K9dcMXemo
ZMLExt8PeIzs0UvJ5gHw81dORSMigyvOMK0FhIS3nv/Jcx87HGidwHjXuFkYsUxx
955KD7CHUW7j02nwGLiMIgEHKAHziUkXkNVvCe2WKgAyfUk0HB1kdTF+Ve0nPVWn
arlaO7Na48fq/XeZMUa/t1ssrPjxSKRxFHMyFSOLuo0xj1+LVf5+fXxRU6uXQzuq
OnuSh95rinlxo7o0LnzU+I1cNih4Io5oCu5qriMF5aAkubFtucby8K3A03V0l1hP
O8vg4hD8o1x87YZJCXuXGY2jT/Yag4PwB1qCDP2EvC4L+/WsRdtuf4OEcvJgJNGD
jQTSZEOv7QB2HQZfNLtcpoC/OyaEMTjgHlFtNI6l28PHyTMZukRwYIvfbxeul3F7
9uA/DKLNwV0s0f8ATALvPAKXvTZc2zacMUA4kCeHjFtkmiMY2fHJ0jAAd9f5ZPdG
hMt3G/6sP+gDMkbRsKukLTb8mjSKJ9wwCj3v+WnWD4tLUHGT2ssNU4pLBgaBavhq
IT+bKMwn2IYoCpszf3l56j1Q6KhBwpz175HG7IqqpKLuQQpqUrfMQLRtdlQW8bbi
WRqpwb5SQ6zB5obI3NtHJt+n7mMKNQmZ7GslMt3J7sGTsjf5gB8s98IMQhL/4D3r
Qprg+ODssPz+92d92acwlfeU6leGtfRYwMrHDMIOpMLAoxatMR5NxxLNfa4ftRCr
FIVYe9LUN1LKvHUeOu4yJmzViNO1pPqABf6tTCN5ikjeUGe+BdPzkzeqMdlD7g/8
Bna0jYyrMO21wSTL638Lg2TZPfUeVTTT6BokuNUxHR6ceRb+g7ROHbvqeIZh2BcE
y42ryL8URth1jwqMN/kiPfiXVE0eEeBqSSVTE5q6eOt8QCbFCk0BsolTiGd/ARZ5
PPg+aaRf5NJYiOxB3JkGwl2PgFT1z5TcVYkgIbcC0csDgmP5Qfbrl8QppwP0mfX2
/YvnWd5/bEkrhC2d7ER2lbAsp17yOLlEsUXu7Wz/dD+Gk2VPdf2+VlwSz/3Tmbxr
kXbfKZtexiexHRm7hgj6rdbBqwam5NwWOtO/z/KbK1vKT1W0qNo4pIKUfV4njqbQ
F8DyFHVMMLGVDcMNlmTNu45zIdoKjWdiyEP4jDT9dfxvJGc0hXqn0slfHc/AD9iv
3WTH/pUcZHsqFia+IoEtu/rJIqTdSpLAQE53IvDUoBnr+XGkvA1v/mG0zDbS7ikp
e4Mg59jTyq3WRKT47HUJh7iuYL3DN/xKr0JCIUTmAz+wuJjd7iewYyAnzHNi5lGN
akSm8HsfA27yPdtKnw2zApOS32dUkAutdLuPUMMZKZL9S4LaewP85T13WxH22qu3
8WbbXkHtXCtvphvD1mDZgmTYR6JUZlbPhXOaVf5C+NbMmwPXsfaxDSW1TNubPupN
cluUyzTxbH2t2zIsQ6+ZIfiKHMmlF3kPXI7RR1w0l9NM0ltwu66Xgvc5Ij3dWTRS
M1kZmus20XALvjKj/ChnzlCg4ABFAkU3aHHaheB2rMQnGrGzJiNKdgpvq7n2K3YK
uxjPK7upW6YBPJz1Yj/9a3V9nRDrMehkOjnZaVjojTTb19OF7aukYeoBeh7x0Tn8
VKqoc4ZSDtkep87qTSqmW30rYPz3nDDQoR53iCBlqgx1+TK7gLHil55qklLTEUWH
FmTv1jbKBV80GdsWVVUo9l+hAyaINxutxJkbOEUkmjItlrR+14r0ED4TzIl/gt+v
TbK9Jut73ia993iRvl4XHSdpEugIW5k4pAxELXjx67dB1bEzECQQwwZQMHYDwEzW
v97jK6vfaO0j8zF0oV7WYwDaPjYAKK3MiLtZJyW8sRgEf2/eKS2K4M17YKEZvisk
sX1HMDlBLr/cZZl36WvnMMUExH8irh+/qw1MfLiOJ3PUalr4CDqf0VJxmhfGBveg
bmasQ+TQwzqHCZsOQtEwN9WmNM71y6sKAQiVXHrPMxsexYHFKH7HFoD6A0wWA6EN
m102qqJHGb5IMm2BXAjgcPrVbL+ZAZlX+kLzRfY83DRgnEvIiGxiWObJiuZzJ4XW
3lKOz8wTRFzGIZEfTu2Cd/AHkXzaZaPxkOTTEeQG7BBXJdl3GYLrEISXaECHDF2F
VmJ9Bkvjg2quO85yPRpw9NltYZBxS/gZg42Y5QWON6XntH88VNJ6D6zwMEMMCfDO
1YBPt9qgEl1OIUncxeP4bBnooV60yzhuhJQdXBSdI/sBCJ2i686DCfRax5f8BmoG
aksS4PcqMxsbZTTPKZmsJ6VpeiQieweqtSXxDJZOez3OZuvJEO06yY9MG6k8AZe/
WjDgTK7VFATWqUnmb1CnYyzH1DHcz6ihJbe7Z7bcfh3S4ZS9TH8HBdIznr3/Kkga
G8gzHiITE8c47f3B6oMwNVEevBQYkl+PZ65uHhxuHrHOl2GthivWPXGJFs20ZqTe
A4Hus22qX4LANLgEnSWoFfFTJG1Nu8lmhbdMayku6L2Pwg2YPRLGx+wHixdfbUDB
2ys8gAmV56uy5BxXttpLqZatsjcmHUGAJCcE4TkqIbmyEdz2LyKcWfMzbfzhFhrz
Soo1WE6bI0ztuDuOhBlTIxmJXq+lV30c/mfMto0M0HZKTKRAeooamexgNwRSYjZq
upjppiXEI/bxpUbPd4PUbFU2t0XIXR8LCB9HeUn4lzVYBQCOGI67tFD8Dih2X2iD
+5TzWzU48gsNsfblM0IelEEknk2yHFDuKpeodDJyk0bP9VcYwbyCZCfdbAO2rmia
fzm9Np7xV2sfvZi4USqv/d2+1mET/QFCXatkJB2hNx6CsidD9nGcb3NwD7+mcz2F
ekpLL6gluWiRIAhuW4zG5zASIcW4hQb2ylDM07+S5IvQ8Is889iPHVqhgZzqkopv
Cm+Ra0z83X8i2n6JuD8ruD18CmM4YePyVZV6B9bflZj3iAsCDR4Hvb8lLCp0PExV
XtTTG6xpVlfpsboAdxA7XwReWuu7eeFb0kMl209+3VuKhvfRSVwKvl1Ynn2RXJxl
wsNH7jgQswG4baCkjR+ZKWvHd/SEXRXmcIKG8Bte21lsm0mEU7ePrLl6NtjTZHlw
ywkqZz6ICavrj4BW42U30mGPoWePbn3Ri/Kinwo1YgjyQ1g8k9vuQKIRu6nmAk20
bbj4qKgFupfVnJYKbrntNNH4Z+aWKxhQlfB+Y8PvJGmKzDJSUsiJmX6tsiiTPrU4
sa0hPGaCFO1TepvcbzqQvspZ865V6mq/mXnsViIv2eVgn7cB/voIf6Hn2Qqxi41L
Ydl3QiufFmqc1+eB0R7pFymtRleKjM6CDNmPbSLmoB9nXxJ/K+2J0g54RwieT6Ms
NGKBc7njKqHf5At56PbYThkF9oQQ0UUrlSU05IN+JFuCM1nNsX3dfW15i2PcBGxj
d2NldDpJ3UW7iRQOeDjb83t+Y1mnq49ndXHEgfC9tsaQr/F6tute4LLcSjUtE8ok
s5znmrQ8F4nccyGOzpH6sDJqzbkSfQj6tOEameaOhwgjn8nFxRNFF6ytuoD8KO64
7hm3ykrI1xhFKkgVPpR2otFHC4f9Y1AEKPOvVQeq+JrkU1UiGF0LKD3ccF2gkV2t
9dYsM5okP+F70+NjF3SjmKZU1egHPdU19Fm168s1Uxb7grQZzf8YOgNYjhzN2opU
JMllYMPENcQOevMq9e3mDox2/KeY2E5hr9L8ciERU9P259EYQwC3AsdFxR/BkInz
Ew4UJ5mW1SE3aYUn6fYIsIK2erBmeJ2Hqe/x5gXjvBdLq2XeDTcGj250+eZg97wn
rRuNuTVTb5xYcOdqgHN2irCPNpv3ufqKacUBX/TqzJ8a+M498bknN41mM5CudYeB
C4XoO8pT+m8sW3fu7SApjwTTLAEYzVN8B6oxsXm7BaYBABsrG0B/AY84S5uCOfU1
1Snto98I4+DbAq8ecAvMmIDi/x/7DBTzfkSrW/Jq7qwrnfTaPkU9r9pV5zQKNnrL
jMTpceA1pXhHBY8foPWIXemjs8WVkV7oXOH3qFAQ9kUk8At34CnGqVf0HOBPQjb2
NvTGW5fNLxSKqMrCVNyjTzxLkBrcTqxvaxa/yl5gzKqwPvf3EsulAX+VUe9w3oXb
mDJLH/mVlbhiDuKOzGkl4SIwDgH0bqTqlkYslZuMzKQdBKtVtFtMqePnMaU6ptrh
qgPH5RQ4X8z/q4SNx/Rx0rFYpLJ0uCN302HaPb58b7CfBIGSzvxsaxC+hlRWujdQ
O0D0hm3h9G4HlP2a1+qHTuD12kyzkLn+lPBveHDfPTfUfIvwYRVHfA2Puytt03cu
RxZHawy5o/S6D9+qERuqDVpoQ0QIf4uVJ/Tt+vllcG35StyR0anyK7TRs48y/r/C
T8aH2kSMIKR2ehg+Xpr99dI4zFcHq8AzU7uhCQUjTR2JrMBvqSGYfqo3HyM4P/nj
7mMZhjgod9OBpMThMyfAHhhNAcJP77sltGVQKmtm31IamzY623ouIDaNwIIgevTc
73pf6TVtcEIxk0TQwjdIF7XCEeS5WHPIQJsXYRcO4JTaq26CvCxsbGplWdxqd2aF
9tCM/wWyS2dCTTBDHK8OcJKVNSYM1JV/FQOa3wab21BRt1aq/ZKRQXLqNaKAPKU0
gxWBJwsPyg9m4eHSFu+7Im08tVh9jdgpnbti9q6H0+Dc16ruf1pyiAZwMLYiUqcg
VQ8mDhyABn6l4WqFZNndOQI2aOg1x1krK2NrnEHaA+DEyTZAHJLu+tlNDIa9DRPY
WtpKZYVV0GY0JqOqTozHAYfVQOSyn3B0Ue3W1nLbXet2QL8uxeDFjDRxpcMiLAdL
UvHCCe2XnWvQl0RdUonVksFVnxvnQXMwBMsIemK8UfJzCL0YMMvlgxIm/jO9Eaqf
eOqepstPG8b3Dr3tXfzZGAH4IvewIVJ4FNxCtS1FZZorV0+FIOCYRu4t1NZb6ukw
Iq/3faR4OlMiZn9BaHRoZ/R3SWD6HWzwpmUZyFFeEOZh+YqKktmCP8h90IpTNeus
Qf8xswSqA/n4SLjTaY3Fw2TZ7+urunjiN9yMJRQ5i1Rle5RYhbVTct1n8qhDQVRI
cjhu2lgNwCuRhSqRk+LpIc1t1NitWwDvqHyHEQeC7VJzw8+OhfwI/mxHorfGZKY+
T8yAc8C0i/zKQnt123/h1gJSfid4LsbneP9rcFJKMHnbuXronV+uDj8VzCURZyd/
MAYPqDNjefogCIXgvPEUR6Csj5kW6YqJaprWxbUllH0FmmKUW/3DOf39vNhGD51A
3J7k3p2wWYQFQGiCXED4334ld6nLBazB1nOqjkZvq78R74QqeqPsXEPtzmqhKcjc
CwkMYYDn3FoJU0fXOANY4q3ccS5osFNGdZKaL8ciHNMyX2zeclDIhBMLPcdfijc/
UIg7PSlANYRzOogntbFcAdmD5A3g9wR7R874Lok2Mk485unIqe5IQ7VCjPnMqnJD
8gSv+rTxCQvGWl2TiwRvLp56xXVnGzB1gMzFbo9ZOAE/jCLgd4+au8tP0yEcRSS2
BEY+2JSd//+QQEB36GC3pzqb5HDq+NLpSsC/AFxCALYE0Xl4/kxSZHKgG85zZiV/
1IHJKIjpo5IjlC8blBbV+xa09jbn5BsCkdwhunAK3uX1VCNp0RKTIw8u2SNhR0Tt
dBoRidnfW8I4tY7FMDo+lwCXmYF2Nb9daOkus96F8MSBFVLSxe2yhTJZenTg34LO
E4jRNcL/5i44wdtng7FeZt3tyDck5qNJdCWDkrmST5Y/yR41t4xleNI2NWWG1hrb
bdl1tjWM2Sxo+wQYetmvyExTndHH7iq+imwmhGd4D1K7XehoCdLeWhxMjJOg8q6D
2tWf+B4J1r7k6VLDdxzhVZvQdwxdyX4CbJORyZjbWk1HB5LSBh5nQZOelL3sB2bW
VvPE0TMM2Jkr/q/ShR4NsKZ9KKc3ssipr/oaxl0pjG+s2kukPP82DIiwkZWMVPn3
NZFGSRl2+urtltSzUyJTBiARhgICNVuucE2b2FGRqka1aMvlc9wu5JaMBWReYM8+
zfJTiDAdSW2esi+jSh1Rfd38WtpOPOpIP5z6XJOkuNlY8lxaPSN945y5wtdrz8g7
XmuYrWVOosyEvzwkGIwbht3Fqe5kSiy3HbhURb6WH1gXFq1cLdg2QmcrH+8CNbWy
ebEOR2+9iObx7LUe9w0FV0ryuHJxhiodnlU3IQswS7yeukuCItuKtrg3jHQwHXjv
6KrUNJe9EVEEfIbS6jlpF+jx/0fx5gJxAf1yx7ZnVFYHtkflDMeWSyZJRAGKgP2H
YgPu7IG3dOUM/BTb2/Fc0a3zmngwO21HtcCCM96XFvGbraq9yFePRSW6xjOk527P
TwsrjlSM6mq6TYZcnGiyy0TIL8Qc6m7AhRPhEVUaT7k2B9g1VH4jxL5TRpjazyuH
ET7vjM2DA0vgggx3Oa1r2f5v04rY/jTwHmJVBSGowvm0nWGbA6PgNUDX73eW2loT
v2Om3hqd8Y1IQEsVNyB26DFg4Ro2QQ0DfK5ZhE2o1qskxN9noneGho6N37fbCYr9
YzA3XwyKuqzwjM6t+Jlf9Oqme3XSLF4uP1DT7vbpJtzz3h5feYPtb3CnAfDR+MpP
xiAdQ7DS6WCOujn7VWz1Gz2026SRyPDlP9hrDzWsvyJbTamW77ZQ5d5ykvP8lC4J
daZGV1h4EmkBJA8HIm6nnj4SpGENdHT5fxANvGlSqrpiYS3i2W65bhOUkl5n1jbv
8QEhortTOhNQ/YQdFMjXgeBTyZUkxcbFdnMQuFN3/UpIklDbOCGJNQe26DvV9mrz
e/TVs2cvpoX1dAV5AnGg/KbbDH/MV9FWf2jQWWcNHBFqBhsqn6YLforjijyEcEoi
eIsXAYirewV9VGImxT2Md//3VYLGdCZs8hP8A2arvX70NGCv+L0CMGilfNeEUCPv
rsqp4eSsHrVmwlXcDeoD57hjEcW0syIo4/uHcpvgbFHOLx0qA7jtHleauTwn5+cX
9ImFCcNJgZA9WrqI6bg5ydag45Q9FlHSd9nJSzszeX/DI2r48BfPVLtDYNQ8IeOY
g2GN4iCDbl3iauKLpNlg1citeUDCRl26Gpay6hyK2E7OeMyZp3HtyGZPFw9KITLI
QMRC6TyprRFynVCoy1qvIearSDegbDel7G2S4Eam5rqdWvKMVL07jKARDMRiR+8q
U7YuAVtNU7Gpj7qGffgd2uMTSMdhhMeX9sXVQ4PX7ViN+Dmy7g1XLKi+62bfpX2g
sCBRQjyDW2v/mAwwD8mqdXZ/MHHzmMW52eER+KKWp/pT1KXVjpktK2jWMizO56+R
3wySNHAzKxEig/F63V7DJ9K3s4QQ5mceM/Ydo9WUbKLFKZ/0D+TjwRruybbTd5D0
WT450saZdBJ4vPt5b4mKCg0FnY4gKUsbcSVRAUp5gyp/nsaI3HyuWLbF+HfdG142
DqljZ4EIE+BUvccI4clbqEvICsHXLfaoHsnEjaO4wLIwTKdZEdNxfMPABb3Hdu5J
mby7zTrVQcGIJuECpwgSuhIMluy6S/axCdjsCRADXbM8SB2vDf2fNtiJ2uVG976N
Cz4okQDNVLT9SNLt/u4mHfCs6x9eCuzgGCn2EBqrMilH/3Ngvrwqz/5kY/O1fx/F
mAiqKQeZse+2ORferiIzvEngaXUFobd1KuXectqp0kdFepq4fmrAEfMq50egIpLv
1W+aGHdjjUcthLWGjmdf9D1PZm0jk2pHw7+s/Pgp592TaMZgG+HnM2V/KyaOuCP2
yLuotCmok9kf5RHdQmC2z3LEXzNy1S3ntIAKhP7ZvWf0js8jqv93sfx0LmRIdQpH
a6xIU2bYAjHkroikCwghiO0a/hNBaPBRL3hCMFAOf50CdJPbvKsys+F40WSYSEA4
iHndbgjRHt8GB68twK2Wl00AbdkOqonalCF11pBNO+4I0TuvFVGmZB9uEeBZAa9e
oNj5L9y7FAodQ69iB/AOlmZ1u5nt2QPaxS/TIkw4t6O3iJm1EPtpDPdKUPX2ypTU
7M/OdJxIFFlo9gmU3YWDF9tfWKTnoCwcjN6w++PqCn4CAp0SjOYAHYKBLqNmD7/L
8n0uAdsnsT0RixfL9KQGXb3+RmlqlyAbn6cGdR5W8OBPe6x0M9731LeotBvBJI+L
/C02ecYUccenLuS/sgiMbF1cgc9RU8vQahoSzZSEdSgrS8Il7VOtWujb4HlV2eht
v9Q2igyTyVNISt6x42KDi7jUt25nRWg/TxP13/IdnVIlSPHGEsk9K7rgr6PXo4fm
k/u8poQdnbmriw5acyC+iU7a0md0dkxJamafgebQ05Hzef7iArnEkSzeBwvvcgFH
w4KkHKtTZZ1U+UkI5btHmoFNeLdSfINensgEHClABx8TZSCYk9PU8HsesyoDyPGE
ofa3rM2w2g6+9c4Zos5DP5TWBEh1WGfcWrrHVeB5Tm0GI22KGyOHdwUvHo8tG80S
taox1AV55dmNMKZAIBzzseINPX8KqL1mrdrja+7X9hEwMCrNKjCcWREeA1BwSsUt
OyOtBHQnvCj9rG1etLaR8ZO3FwSxg3PpNYXpZGpEsL1ttMgV++E7RP/lI50h49cl
YsBruqijEkwjSLkKAZRLq+c+Hf01N68xgbSsMfKCWmIxfSLOwDoobCJQmEOOUg5T
0aRJqdGgQolIeu6RtjO6sFZleLmI7xiDf9MHyWybt+qDBq/LY9teY7v7fQtY45f/
yrRDFxhfiVTfOaie7WDt9EhkoEy1jQWhczYqxAwW2PEEikjsyUrbfVSGuqV0NNPQ
3ixzT6knIpaT+qAfFbaszhT9tPrbKCgFW0PSzx23UKh44AIhsJQH2Dx+2DO9NFjh
sW8U6WAJ7KYpbQ6uavnCzsDYoKN82IGeSiXydATq7mjzVXRSJKON0T4lcwq2HwY2
qbeop/L0jH43gK3s4taf8URkxwf8/LtnnXYVcyJ3s2InQjOLgem1skMOZW4AP7tI
z6Adrl/Tlehva2lzCTY9Db3c8iEim9qy9KPHZcrltGfDQyi7MfeihVs7BxDSjOKO
ycsVgALp5pusy9HgyUgpkytp53gZv7LFGZnphnuR2HfuBixq24GijQb64Lp2/8Zn
eOv+Tk3PG3Z17Zi/T2OZfVHeE/RQpidOROosme7fcrjAhWww/gPNly4Dm7bvjeii
pLIsAlwlJ34TJHet5xLyVyk1PXIGX2OsIh6VCPszc4vMvgbOHfbvlnvxukaWBRyd
YHl9/7QAdQasSFNUgDNwVlRPDmbd0A+uzNc0ug/epUmmrWZEyod5EHdxMx7c5X4Q
cjmilThYzmVHh8OVTAAT3tHvBW2LPhjfLHs0FjTwGaRXRdINqoVnbz9LGRVl4yX9
RJrJkrUBoR8GSMKor7xtaaOk9pxq7sd2QBQmpH2a7MhDGNVhNgi99gcBVvCzaK4U
d97St9FeSL9zFILVDw4/0fW+nFVJolO0++0myqmKqef4mrM9Tzykk1iuhNLQFPcz
EWHXxw3nwBeojTOrzbgFmnewwsE7rwiVyWltVNfWx2GEkoctr30Xw0taWKdm2uJZ
dJGSOPpUUDJECKWy6078dvbXDH3+fhTX3GcP0FMWwRt8TYJNUNJOXdNfqRKy+CHw
`pragma protect end_protected
