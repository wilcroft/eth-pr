// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:14 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FprV022TJIxpYdtpqr0yxEOwjEZsm8DmKNX0CX4oLW+LivR+tYhwJT9Lcgm095ot
31y/jTrW1eEkkFjofUJeHvfpLnfNjqvgUxqQrtsvtLvc48MxxLwTTGfwDDXTjIPA
eFnZv709fZvN+fpv+ZBzXGAuulSIOwnZFjXm/HaPWPM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31024)
qG6ql3CUb924iZ9sD/Ix7tz7mZ7AmoFbm6fzA6GoGICARj8lIojx670+bbK0tOHw
eBaF2Ohxq/Ili4VT4eerqxG+3rEYebiX4trLZ42HFXEWUd1cNURvHjP4QOOwIa23
3g4eMWG8IZXA139S7HWAcIl/dQETEDv0znr9/u63QZa+huyeRkqOoi/gIEH0Gquc
Hrz7r+Y8BpngCfeVwMRLMHxXdLbGv78Xni+G8k7eeCCELNf5/LWbQqn+DewcpoRe
xC7AG+A6RYQfvQyaczpNPMAQI8ZVJUEG2RgVRYyq3uwD7eMv9+p+wzjalacjqnoI
7Xunp0JYnv3ymFRNNVjjuCmLtLqcD6TyU6OqvVz6cauDu3Qqcx+JyeiPsYUUuxY5
cbocdlT2JOank791I2dQ2nW4tsuITjkOCrHkFqvxRjAPgwNTb5PKlpu8xxZU5Ytd
yLy29FBros4s5kEKBbWif46guSkVOqhxmqISQi8yqvSNr+ElDaz+hwN4+bc0uOl+
fLVGFIDLRyK79tBBvHzrI+8JPqnpctdUmDFFdpNPTxlUawrqHz4IYLZHXTEUpiCJ
gnoXrDsRs0VOxF4pdM2gJmxQFT+O/KFSbnbRAfADat7egI2fbYDZAj/TEXbbmWaQ
qKY51dPSu3lHuB8l6MrG3Ec9T6FnfTcO3BSrEvbucsKMz9Q5iOXMZiZzeQN/HW1g
VpMX5ZH/06RMOHUNdy1Kh9mcJznPdM9fR+onjg792hAmGN9/HjTTC97XDPKPVznX
sCn680nvG9OtlR7IsR+oVF0/LViHWrxVpzk3NxjDozSzEjEowJ4yQKT49ewGyISU
S/jQIUOUPFRtG1olB8kGpTkcJY9j9cazEqClrBkzfStHc6sQl6F9qSzG67oT/QoA
XC5O5nP+M/esC7BdtBtevvlo/JDaF7VgXeIjP8QVWWLCjz78V6zNDILOoEGieDVK
Xsf9yyFg7m8NvYTXj4rEmA1nlIv73zen1A/E6jmEyXxmioPD8MN4B22Vmjb8DwNh
FieQ2VvAz0TYnIaekKXgLnknmC0OFE14mZvkDmJBG3pnpP2X9ONulilOu7qNXLVc
WdXXO/HxRYRbJZp3ESx+HvH9wGYr7Klua9D+Kt0FpqZSGuwbOtRad/LgVcFWUBbr
2ZerEDuMiLxV7dVYNNpXfPX+zqCsXwR0WAWvDnaNKRqI0PgLHh8k/ZjmHQ/9fjPp
kYLDOi7t7s3h3QuKtgiE5eKLr1MFWtkTOR3LhUEJRH+vrmQWLuM2cg4IaR+PdSkf
9kUXOODZ8dkzQBjf13wFLtFSxTLWhC/koz2XQsbYZdMKCZJH01TOiHgt+QfG7sz0
SoRSJhErrpXKggYkcHknvp7zMK1PAWdDTL+8ZXX+mSInBd7+AHfgI94Q3cwAOVVm
KdWHi3vEJDNLdMF3EZeYvGEKL0aTtoTHjIG0xlYqcdBA14xb8osih2STOfgqT1VO
9X4k8ZYVJDjLOWA/n0q0Zo2CwddpU2G+ZMwj/AT1IOTa1kLaPdjftOdL+RpsnoZB
rvooZc9i9leiyPUL2igNiC/daCZuRAtwLepedi6z7kYbY9ewIRkWySJxakhz7NN0
b3XzIuC/HBEs/BjiM58kryZ6/2apBiCTJVGwUEQM/YrDJcg0CkrlpIugPx0V6QtP
U0fGk0n/tNTywgtHw7+V6QN5OKO72dcR1ZWefUgMrUK8lT4p1ZqqXEzq3wk9GcWj
uc8pb9OYSN05FmfxyTvwRZvgaOs2OOyNw8gjznODXkg2A2R/G3wvQOKNsQz7RbKa
B+OGdCVsh91njYp4bKdWvm9UQGpKrg5ewO0/8k9eoy1QIW27CF/kp2ExIdeAZM/g
9i0s0jThmXlQR0hLLkQOWS0iKRLfiU9+CK+TAifRH1t/Hpk6GQ91PcNnPqtvmtkl
iM5fPEGZTKS7Aeocug/t98+1jarM/xGNlhncLA8st46GDaZ5DDfNeiQ8uPa0EMbL
ZL+oiVGtuBdPnbO2I9xd/FhBppA5lQLnI/QrHltP78Tt86K3SaehYSjNw75SjRKv
K1Bts9D0BptIwW9/P9Q4SSXh7XAXgOqRhUXoWKi2bYdn7w81Tb7Ymcgp0yTlHUfK
4mMO4BfxxAUEb2Gac73dpdaAUkayT+bAv8zEJSk/KXEVhVqVWZFyBwoulD4yYk+K
HM7sineSPVu7bU8Vy42ZbvQAx1LwlwhGckjI31Je5Amo2YA+VYSAUB/sL382MA/P
hVzLxraxlaGxAu9k2KxplpbYcRjK0FcC8WWqlPXIQ9QqCzyRl2EXlwJBG+FGwUMu
VPT8W5gMT/+DFWICRQ0dfmEkMa89V+39PqCeorFcV6lMp5mQl+bfYsO7Pb/yhTnf
CyoAJggMS06l0ddnC2uiA547Z7RII4E1y21yJeEHCqERfFmRU4J8VUj3EsG87rDl
E0jyQ+YU7PH+d6arWSfXXHigP/9lKdxIRgs3uIDZRNuHdJICo0SRPB/xnKVWfo1s
OsbuCrYIZHgwQTmk5vgz4KwrPB2Th9XV65e6Px60M3NN1ccG7LCcfcxHm1dlprhd
cn3We+pMnSKdFdHtoPbgyC2JTd05ctEIr0nIQMKtbnUSrtpj25AF/PJ2Xiq5bl4g
BXdgMRzET41kFkP9KhiLY5jgwuYaSXoM14Hsv1td1oU/h66laK2iXIJc4VKytHSj
ZTQKJbA/vMYshW+xtbenPFzio3oJRv2ouv/sAd4896WcG+MXHymfodfpM2rJH1Gs
GZcnYxanHRrWnzGib7Vvg2899xlbNOczQhF97G/BoC5/zl2V8g7d0e65Usnrpqj5
nOqeLqsLmI7teRbUQWefDJAuUt65SZhiA8BsMI8DE7GGS9Le0cjChimJWDNU0vS9
XUTySR+514XnTUeO0m0Dv7OdTgTTgFKHqG9iLdXw8S2uJ8bCdTTTwPIApmGLF/5Q
SrH7IJMJvLAelTXQfjysEzbkZFrP4DxsNGkyUWPLIqrO9WhrTfzLSdJe1G51vsQx
pcPL3M8MnD60B9t95X1S1AWHmJy2ZrZ4p0zLcxqld/eQc1USvZXd2bEsE+uv2/i1
sqc0U/oplQbVyajOBQBqoGRYdkgfQ/v41yIgqVIzIsnQsM2w34JYl6xVCICPKOU8
LJ6V5y2vpk6G1foWd7rV+eAbfz4WqVTrjs+eBMwVAQB4WK48m53eGNF0/h2d6EAO
SVzTs/r0AD0A+/413sNa6Tt3Bf0rY7xExcDipnSUir14t9NcpFxCVtci3XwsKNKW
2Ofz8+avkEXyZxbbUE7P1Ccu7U4BX4LrLCM2drUC7gh02cK5s68JjqlCNGxIHOG3
85Uy4sdO2CxjLlYQu9BQsb3FhJK8e2572ojQlvqGdSDxSYKVF+YXKba9LB/SNmiS
Xcj7A8fSVWMBhLn6K5B7hNXdCIhZiAvsY2sinKnXqr0iM8P3JMdTzCoyQRChChac
rEUxk+ky2LgFPPoyP+grWDYal9dNZb3EArZ51H4wg2rI0d2awphWsfpaM5962nRT
4C5tGV56Ggm8NQI1O+5Rm8Fg5/qV7LIqrRLg5GTV0tkRXHDi6ucWBcwspYeYIXja
dl19aXvdW2ttovL6mtlgFarPbimpROPERwWJPYM2ybgp7EziHaIzq9SWK1TCP8KB
yKk4u62g+tdo2Uiz8ppHDwUAhSVLqKTAaNUkZL1+un0PH4ywqhVLX72/A2lljFw2
6tBmuPRGA3d9WqDPjhMHBtyDzMFLQnlqBQmgIek2RlaaN4Ra14Kjpv3u+gX/siib
ZpF4aeMApz3ElT6zULpKf8Pes6vHpnGbF63SYFtyYr14Yalpc49W0i81+8kO+K4c
g1s5sGxkKujRUrKJu4X42JCffpqmQIybRDLYylT6Wr3sHetq4YCGhM6Za75JMKtH
ilR2PBnetAgxG4RoN8CDmj2LkHZez6GBxa8kZSZw18Fg3SXGQcI7jzOq9J0wZ3bM
Vy8viwjTLYPo2kvXG2rPM84AWjr1UNBgwxDyCi//VXUMMSDE9QtyS2WmGSPtkIeC
8uyY6E9Bcg5q1eRAvp2GsKZ/Hus1pOlTZaA8RoszWim2GdyI9XR7MYW4XVdEqbEO
FyjOADzOKQGpk/EODuEMmISdwaUiQoQ8LsWeC423DSnnMTxTBzNoDDvOYoFtelTL
fLW165uZnaKrd38CuiYOVdHWRqXidK/YptO7unyvnKOv73yMZjzRE3rDFnuK1Jwp
I993Ri48C1Wnw/x/iQEASW5jQmF4WxPkwlUmWk0a/9Z6EGI0ORkNZYuUnrVa86QB
XBHd3y772vTNGTsNMXVsw6GMI+AsPKQYX3I6MSeH9P0TvWkbYdlh0PNp2WrDYRR4
/LMGQGwagSw3l/ggvdu1w8P8Osl54PIK9wcb4a8oP0b6S9JND+ojpYzsOsJ9z/E1
FZRNLr84T0RvqpNrg4aQNam5qjgu+hKEp0TrmTt2K7PTO+ILltT+a27iuMof7i1U
AUjArs7LYB1dp0ABSTGq8mxWE1Mtbrha6O0IX18PR6NwJlNqQ4YCeLJpQN868F0k
MOq/ZHvNUqXTtVgPIeG4rg6c9IeqamDcCsUo1rcZttryH24y/yh6vjqMZdw/WjDs
RcMpO002D1gHMkcxrrskbW1X/jmgtL/6RzafaEZyAyUHYmFCMnhdJO2NyWt8YWPf
/jBe6JFneRCMy4dmYVdLpzkDid+SSJu9Fom24m5K1REaJD+fsoVXno38Hgw7Xu7Z
STfDVgBzHHwJ09Aa2nPU0J2Fg3CLU4woyL3G+fI4wCYPO7P5WP+ZzMbntgLlyUWA
ozvna36RA3YxCB2BMmyBRXFuGO6aQ7DN38fbrJ42BnjfgP4MUzlKRjrk9J5TvTah
hE934ajyij43sQ96t65m6eapv6u+BZtEaa8Bch6JPZFw50BTgZx2ez9vTCeJiIHn
RrC3ljfatrpT1ZOjHL7PWrenxlcBA9o9mikc6heGeq9/PDUZHp5k+VE8NSAK/+jT
akaYItCh9zGpNIXYORDI2Gt6IhLQa7B8kky+Xcw9bQkHPOefnCQJBplcyWmeTW93
guXhq54JjY0TbGq+eHiMYIqJvHu4nXVSqSfM5ahHNDtS464wbUIQAcFHd9r9Vhsd
1B+k9QjQz70fQRHLy22S2Gmagx8CDKvKjzLXNQr/NXfym0xfsWfYy6226YUpJnAR
FCm7a9fZ/hyqjRoEp6vDXp4yYDbbzp1xj76mpRr+uHn2NBYXa7rhblwx7LHsiRa3
XJKUtL2MhGKo4O23DuZZvIGoGah0YRIDaQz6iSdk6Ww8/WzuExr9Yc8mGpqLjfjY
fsXHnYxbCzW6qI+Oi4T7C2OHmIfUGqQJrIFw16le0wTogLMGCdU8DabvcRXjWp4O
FjDeoQBLy2iX222Eppa1v6RBcLOQ2WlxIJJRJylzaCpWijWKv/f32ZAx068bozyn
CFaoDesRFs5BvkT2vLb1ZnSr+huvlHbFtxwCdiVcmTV2TzsIPCZ9WmGmWhV/l4cs
yoJ3YYkIXhOYhvftV063MooB85t2l6QCIM7isYLUrZvm+HL0+BRZg/nXIYtcQaCG
B/OQX6xy0FX6AB/FfaQOaYq6IMueceY597ClA7yDYX1j55t4UWU9iPc8qNfYpovA
hYm1chKJMYH4IAXp658rSIL5I+ZHKXAwHcguKI/n/Lb6aRRQB+3t4CTwWPtM9TEt
51jlC5+aJPtvzYlWd8EhDeU2D6LIDbS30hgcyEfiCYBhtdG9S1dLcGgwbQE0WbRM
CXLrUckMN5gOO9oNZYvaVFpNhlV375nUl+pDR4fBD9LdN1RG6u402h2miSMvhIqy
Xy4czz1BOHhbkF4gpThya32pNGH0uflEgPwfqsjqR3Suib4s3wiuXhcz05FZ6oHb
s5Pa7uhsoj87lx/JS49bA1haTN9uRzamFtONdVwOgha2FleNYTC+9TfcUTUAmf9I
fuzZjvUmiA2PKHMo/N1aVr+FYyiligqFgi9FYDfSeBpk5VHNY8Sb/76abl8WUO5D
ZkP1TGM+plsQaKRes6iExFzQNT6DRetDtDx8UUkZUkz9D9NR5+sgbpIBch51B00E
JVNUBWpBIZvGRtLdabgjPiR1ihqPXctYugh8sdFo6aXdIMBCn9gbODuGvlg7j/I/
gu6AllAD0fSTKLGDzkVeNPNIjem0tHxVFHZmavG+BcDX1R8P9tdRhosqZuFKA+Qk
f2UvTyAlA61FBbNlpUMVwQWx+f+hIBqU+tWu023dfeGxi9m2oshJkmoviYlMlo1l
LyozMQcf991JhtL1EdISTG2KggfByLayB52FgpFTMGMYmVLr6I61AVgiI2nXLZow
zR+MhbO3mFI5x145P4rxSfU8Fy8aggLplN6ffo0aNPURNBogpOAFmDmNqL73eksj
z+CbU+3ngJIeejB2+Y7b6upG+moHpLxfnRE8/kd9cXCX9aYIWlQX1KDLlCfHw+7S
3kkmYXKJ081+ry9pg2+RKNnnoSor0rNO2KkllwoyUyUJgEjr4BRAT2rmarKnrXrd
JYlkg4AJoo+nQn52Dl7sSf9mviuOqNrFbbhNIyoWPtgmQ8GJwIIad4L7/u/nazWB
22nKBv+FnW4F2NF3/+vjwg80i7cnC13GdSNzguu+vyo0IJnYzG9fEZ0bAVFGECBn
ZAADmXYuohEzIRbYXkHp07A6vrkqBoArbzzZ3gIOkHSfGIOX7qTOPZy/zCRV5ydQ
TAPg4DkXgOt4cn8Q72fQaAkCm7RtCewg5PPx4FTPszh/r0OHo3Ah8wyIr5Ci9As6
Hr7kcd7nOVsVH3NUK8agYcNy2AwCjTPHXZdQAf7MF/3vw7Y/RcF2xwaUp5S1L5hk
aWebbXvSYABMjXanWjdqZO4ZFxFc1gfcI014IZgKh7sm+yw8wZFBYI+YVxMuUFIW
hTuze15J5u32ZmvwOs4sYGh3TVgXOfVuk4xj00c9dbZh6XUVXfYaxrjmPuBO4/wE
gB9UAucrpzkScSizyD5K3EzB0aUknIEg4CsoB+PZohJdq+TfZw0IhJu8VNdtBp9c
S+vLmJ8X87iwTdawLsyBVFADxug3577rOt2VcIFABjbszVZ7fe38Xk5t68+7iK6B
yL+mTqkc/s+zFnprh39uUCM4gC+pwhUxQJ687H0XVChHpbRr/Yr3kJNU4U9cSPGw
LH6PcKfG0tMaAqRTyD5pEr1K27kI85YoBQ13lBvguTVeK8yYEn7/YsMcQQox798q
ydVvVb4MLGF03DoVJOBfRIvG+Uj8x6Q8IUEklCGX9Y+x7t2bDly7E7AWp2+7oSHH
msryeTqVG5vLJ1J64jMzA48xWNzNcQhCJ3Vzucd/d2YSntdnItjMxdYowmJjeMvL
IRXiZ5lmGySFLIMKL6d7HQbcLgVRi5hTEbG7A8CnMHBm+iDt5cItTQ+10fYBR5Fn
sxT6JsaNcqESRkUf290LfEQajTAKF8sSxBmVgmlt3P1Tcldu6pdR/wgwWC24Vlne
W2+xI9a4BRYbjMORL7fg437hNzDROfMYEBTJPuVXLaqTiYuUTggqrcADrrZ7GWTs
NGj+hjZ5lI29AVeSWfV80EWMIwo3d3O1UpsqWgTRhipiWg9thqbAFkBothTUXlJ9
uGYEFvZwEI/cYxyZBYWzMgzE2nAUCbQO3jzaMb9jmAHyIbquq0/+4uVLIcOASokA
2+Yn1wM6v550p6NBEUzG4hyHPCvvNIHXGJAsxRsAKnlaSkbucvH8ld9x5Ir/iP66
c2FCZ0y93XdMR4x5m0jpBJhUzbrqfVuVSiKyir7oX6RqoooyofygCFQb6ba63VUV
fSUqhUllnY+zrlkBYAEOy0TSktVDuK/PTXPzBu8u7t/Ed7o6SsOIIluX5lgtPDAu
8O55pm6HzQYJdNDVgorcxmILJg/1HLgeesSyhOk/E3CKOBud++CR0qsBv3hjUxy/
nualt4x6QVTWPDXq/EgHSbM6oUwCV6JlP60S3/fbGSREFbJeQiGVOBymPIObTzEt
gwMdv9K0ID/R89aY9tcZyaSRrF7sp6o3QunlIJoyFbDSVSJYuXGSleYWUZUbMTEK
Etvoz1y0XwLEZXT3DDzoU9pPRHNL7sY1eH/Zd+FFeKt1k2xLoKAKOiHIrBOGdljf
XO144QRYgn7YsHL/xZwBigues2D2SIYEF+KicXl1lq7sbDT7vX/pc8PQT1FAM+Sw
Qefm835lKIfln5yKsQk6a9BZTftfeOx5OubAYlVd4dkkoTg13l1+b6QaRBybDM+/
JltMBlVUJ/FZYZKXFS++VmZNFixnOEWk4Cl0QJ7rW24zB59zfddOleoQ2Q8GK3Aq
JipzH8wUVNXAr2IkHnXUq8DLw5HrfU7hyGmR8QFfBHbFmq30xmS8tWY9xRtsvVPx
/cD0qyZVNMY6z7VjWv2dnaemaOb1XireEqQUJCK+5cVpwZrRDSCES2K1rL09zMzD
qB6jKO/THvBCWnNTGq7swj3SfxCtJByjsVwHglE8XYI17zCTw0yZ/GKqgIh+s1Rb
kySyVC3qlPDtFqS/ofKBvQyfU/0keqXY0ofSrVPRcHQKdd7fsmiVW9vx6S2ATkGF
ygJArxaPHhGfVNeIpV0ZSmmUuovziFivujWuH20x6xVwXzbfixhmlIFAuw+sdaek
En0FWnpBNtR14Ovfa88ZbAtjO6mpYJ9lt6F/f4xvwwDS7jyqDAsUNPGhVk7YaZUI
lxOLZsl9guVxzJDAloD3CteXgniyjqaAIVXHS2PA8lLphCbOsEt9qitOfEBcJuSL
5f0UDtKQFOjpfpycbf7u9eOxgEUYIeGS/FfFar6garLr44/qdiwjcokHeQaUEBdO
ZeNGHlRYVqjcFVi+EFCGOZBMqU5aZnQHF4eEVu4YUD4EbeVhpagFVCpemv76HPbe
FC4sY3tFMwl/CUnXMVL40ZPfdxLl+K+Fu+s4KO07OcrgYcfPwcHpUKQBBVM3ANSY
U2G83AZBU5UNLsutBCCgLqfzvSBNH4xC7QZPRxaUHNt+nymgEttUDkEgJL4kqbXV
3j0CAABT9TKrQ2SmafhTxXCEzqy18kODn9+/6cIvlaYch2jHkEqHplYHN6AgIIIh
+j6rs1De3TZF8J29H1viAQrmH9jW6azpV3taON281D3l14oFo0hcH24CyfIKeuMT
LNuCHwkN6uikuj5yJogjgq1SGyskKujZUW233A058tT99KTlkw9pNCBmAqM91ahv
1oog5CaRjEpIwsnxFygzHLcMKVWl6U0qUe95P3BdtTZ8vYyII6O9ZW806i9X9GIC
sCxSZwS9nNI9DJ7SzvnKSe/AE4CBnJEdvosqVxqi/Q+8riHk7fEwWHP3/HpppOkR
8WkU5Ak1oE8wJ4H6FwyaesPgBWtQr2DxshOjpLF51msk78mGQKk5q4ErMiawPhks
SHpkdK0e17y1YODydOPJdKF8ww3SSWoqJ3vo/tI/tpfw5nmGzhNSOvOF255WXLGI
mELoxBTymbAOaj/0BrvIribGmo3aV615BLVtHs8uhtRcVqEPTphaer/2bWdcKCJC
145rlFGZr66H/TlWJIeBXyY+GLupGo+eVAw4FHpOd+vbcoLo8Lz/E3pO6c6uq7GE
lfspGyLkbs0rtFaLw+OZuKlp13BwPloZELJcTAqHcMRNe+rGpUJoLlhFU6cgin+O
ZYBr6lmyfQiMNCXIAsbfMQHV8UVvaBTZIn+fyll7oAp4Uspbb35sp0dm4ZCOxmr6
wiAWvCwJEcTErWOVavQaaqbzzURaRW1aItUK4ag0WLrbOYG30iPuXIr4tLDO5p8z
4thX81LtRdZL8MobjdLfX23qBzKPHCCLskkADgbdzOnw6IW1DEHmiOta3/GfKFNk
K0hev67vcBcAXEwCFl6a/lseWpztcHW+W9f2PO7cdG/dmGoeqsUk5C+IELvyfoHf
ITqbPcYPvZVE6PFGTBxIwOu7KqDXZ7hYBvHisHFoyg6lhrYvS6LJTC1H283Wnj8E
+B+9s8QtUE1Y6cTIzdSwJB1bXATCJdc7M+1y2bIOwmirj1sEOx6nE1Mk2kzu51qs
u8f05/d6g8ZHJS2o/gwctTsSBAw8w4Iv58y1zCtkfPgS5ip+w+xp6orylkkTDTG3
/JM+LCw88nLuIoGrH7utXzLCMwEggV4vF7bcFWjZp8/YtZ7Z+K8ACQmvgb0QxDWO
Tqti1ioVsFaVm9KiKv0y2cvhihlb1rTvlQrfUBebd1dKZatq0Bx8AdgR29Ji/EaG
V1te64oLzyHSip1TglG+P/GLX2lngEiXXqBv+G7K7gWiJJnig/+nZ0qDIOuzfVrY
+2xn6LhCQfYzmAx8K5rmxHeoZ+hPoJ1kRDlMASdSV1eLmqpSlpqcgWibQsbDbI/Z
KcIvJPdRnc7NDTTEz8bWW0eJY2y3m4HywZVoG7fkH2j89gc1flon75t3QwfuDtow
YTx4m7kvQ87RNb/b9wT5I9eKR2Weh2sV2NNhCZ45hbySy2wvJ867gL6rwR1+CUHs
QbIUi83uBszl4EZMd2xXlJ9AmpsDsT152zqARvrefL6eG+rAugs6G0xJ+ga8VdRF
NqJt0Amv1aEyRdY3BxSlvyyofwDPbp4VNjimkye2Ayvh9Z7N77Wv7a+fSycp1aiW
W7MLu16eGlxaJg85HNpJErxTzxUY4Mse5ZDZjcCrG6dhW5oKhE9yKWolxjDqnvdE
ubeUwN7z8zGlBjrMttZcurUXP3wcrYUMKKvmSurSf7dFHHpyG3mzr9P5nQrxcCiw
7Uiyc5HIjnCZY1YJLIFMd8NDqsgqNwdhxt5g+V5LLewq+dFqwmAZ/7giG8+7/Eho
cDheKIYTMty/RWw61TAJ6gN9slXQAoWxCFOnHoXG8N6G+AejjJlvmr5vRSkSPwTK
wJhZjIwdPX05S/bm96vZEUzRw2lcV9INtYwezTHs+/SyCPyS7CF2uOQbofGF/YW3
uCt10w0FrTV0IkkrbjtBxe6vJFruPTpBc55B6/phKT/3NSmwniaqy8A8RKmAUMAJ
O1VeV/qP/WS08pRMLi1lQ+7nfbPB8wE26GORw9mHmio7ZcnScFttwJii2w4k2xIz
j0thkKZJWISP97ep3sic8rOrZPavSasCXYmtI0242IIsF2jZ1E5KqUfN1ug3EmIk
WBRlHqBSHND/MccyqgMuO6+B7qMG8szC1WtfQmD5Te0fPkdwO2Cr+88nqSiAf7pL
FktQRQawPpOG1GWIzGKn9BpGFbeOUsiITJeIXqCbdummy+tLvKZOIFZjhpZe5gw/
TURNphrNp9L3hBvtKMw3tQHKEQGR/tLeF0+9d8Go7F9r/xidi/3Z1zVyIJnOz+Be
s+/E+2M9wHQ53XzAbJiML3SHD0eKwCTaMQfj2Ik3/xJBWC1iZVrrikCWGxoEMCGs
paGegW+Dtl+iDFTI13wSfBXWcDee+tcsVdR4fvYCJgAjcCDJPPKxJ4ekBgsiCENz
hrLdpMw8pEo/w7NeGDZ+piaqeMDgX30evVEnikYUDCBFkRZEaeZR1YkIKr0eQiCC
/WGaksU/suEXxWhMkoLGNBYcL7sb1sIJB8OtXNPdNjb3LBx01MHeKv2MXa+6vEtK
r0BvP6gJhwPYfnQ/Pagnqslz+DtAGfxoPY4hyizKUtibB5g3MqJl1X3R2FotEhK/
QAYKIgdnvL5p7pghW9T2GDsLdOBpoHiVFHAagFt+BfSx1Lc9jv6t31eekyJiAfDg
uH5lhoySQGtcfcCJkQjbMrSunANwT2cyfgOW3Vk5Na1Gm5UfrBn8x5mwxnlrTEGW
w1yDhEOwYzlF3Z/Vc72plQLt/6H/QS8xW+W9MC08v2DhEdDchetBaZG0+jE9id4/
J1FrGRmg7Uoxu5lTC1J0ROQN/mxtKN3YUWhjBZNjZqy2NuwiFqjO063CHiOqbs+S
6mvviQVFt7BhRlQvDdWdm953/3zRAiiz0SX5ceL2o2oExK6A9kfV/lSvTONNOvGH
LAMUt6gzGwcT+sVBjyjP7Lwkv1mRKjMXVBqD5EBWKX/YGstddm4Wjt5XbqeRYD5x
Rmb/o36P3rfsMlUIzRZI1q27vzkmtQ1uY2KYlqnC/VsQpGxoEmg5m8eqWsQqper1
5G5XMs3YPjbW1MN6jh/MCVZQs8NMGVtOz5tRoVZAAudivxqZ/YADgS0sTlbEum5M
8OZnynC7kCrIEH/OvBTN6uAwQCVZ/kGQG4Kjgdx7GVRba9fRMBXCcFGgPbHPFpkU
rn/hoQNXQJxljmf90v4leEs8hPkBINQ7chu3pYuJ+twbhsE6xAhkEf1JJfIN0n31
U/vd1byYNZLOLKe2G1jcWl13vaTISYjDFbQKHRyLOMfUCXQIKItBOGf4eD8zMUj7
1b3hl9WatFPs4JJBCv0sBanMnMhRuMcVn8LdhRueqJ+cMpZKr8z32fAGKcSDYH7g
3vHJ9pZztIQ7+fljyTzb5mI9X/NWcIcFk87iSAB2YIF3HWdT+YSqcV+3B+mroLyI
Jx+n53hHXEmTblwxyMzQ7+uzO78YcIhgm+P7gAxdPhOZBmSzHkI4kqBbeIYWAStU
H0bbfKHy+rnfyprB9YJL7n8nnNBaRN7wF4qBWprQugvfflhwqlGrFHwH35Tqi03x
H3tKghW7+r7IRPBUBF/OYAcIWebuvrsu6uN2be8heRx6zvQ3o+FV/vn7tsboEceQ
fgh7MEtp1J2bL+Mf3s3CE2s7m7ED7hC0wRoi/UUuMpgHRYPo3IV72hq/Gwm4LTyc
SabespbI1Qk7lRlwcrJRFMmgAF2NY38j5o35EVXHsF8mD2X059rGfWq1b9Mh2sXg
uX6RzPwjhJ9AO8FMJJ6wuHAbC4PVhFrnda4S9MfLdnGKJJ2XKHMLCMpN5EerItlW
0iOOWAevn7jvpKICWDKKu9eqGo51ZFupM+KWKB9xomWSRCcnxNh9hjjNRqTCDQgh
itZabUQbGSM2lj0pbJXnvr7yAufaZU7/xUlB+F7yXRL+nDxo6ZDQHyRXNX0htlw2
Sq0df4wlwHaLbnG6nRhFV3fcHp7hdzAgshNGgPCUqB25VwhtiPoLu3EU6jo9sLHr
7a+u8z/7bSh4gutnBMaRmG1vMLmBDqI/cI6p28MWogWe73U++enu1rM3sIHg6u6O
dtSxhbImGn2eT+hAcP4GU4MFWmA+ZBZSr6OSCcWUrYOF4YwqTHtmWzyJM1eGT0JX
73cTvaKo2hHl+ETfFo2bYtLtIUrDfxvwNlzt1fHc5Hj6KkaBd2rTVwTvIm+TESfT
Br6H+P75biNcLV3ACIihc2Pz+YQ38CMUMo1B/f9Bba+ZY5581B2x5m4AfdpnveAE
gjQUbnyg8lXD+9c0SjnlB4003FxmGYDOwVqHWQM1DPLAHVt0pB+Hl2UNdnAozwfw
orJ98o5Je38LICgQWVVPNNjqrMzfERuuTj9M/e+Y/1CPJKahkFeDBkY8FJ0UiWVY
kA+K2I6C47VhAPiRf8jIIr8aW6l5rnGUCkhFZtP5z/vj96zN5xhrQvOn7jQCgHqZ
mV2tHuQdhWP6ORJgPXupHf5bHMuBFhFK0JtfBDWqSUkrwq2cVVpqgGCWWgnITZpA
02QUabs/Wtko0kePrgQSQ2Y0aPF3qfjrwLRz7rYFQZM7uprslg9eZA2lnypxAWE+
VzK232pVRj1cZaDDw9a4TlDOA40IWl9DxrRi/ps+r6BX0nh6IFK5YHK8QO4nHgbU
7HwjJ+ht/dl6Vh9ziZzp6Y1S6/ycvZi9D9PRE6hFsktgFjM2a+fA/Gxvg+nDwex1
Kd8ciZUlyZX9RRUYYu/NtT7STTO+/1+W8TFs+XimpFpNyXBfCUuDPp2njdJVdVmN
8YdXNGJXWN0IP0o2kkHFIXMwQMRIFwg6h6P3PhBgnnZfhkccXF/PZiYp8qxq2l+o
PJEnOOEchUJ+31SVb6YHzhnw2YTdWjP39ekqTwqdrtSaXMH7aurb3KZoI9yjlYIX
e9ATA1ghSS357yZZk66IN5Kr85LB+BljGB8NZ9fpuNe7jQtW1Ig8sqVODK29q5bL
hI+bE0DSf5M2H3B560d0FwAKnGB1yDQRqzlbfIfBMbQCIUgCaFz+dY8MgxXr4nHS
OONwNfRIzMv/a5HkrX9bJYtvdHbPj6Jjvy0jlQxz1rMPOAgktWoFjBdyDJpJX3NH
25Zm1KqxSTiIdO0ZsGzhzrgC7OV2MHfDIlnI5L+1vl/JPxmQRYn1hRDYD6kfEalH
7JtKAMmmIucaR9wpzwpf1VYHPWmCshh0rkujATbAT1RY5+yvGhIgks3fUa26b1UT
x8qSFyQrmZ0ZpMNhi6w211b6qadd7RBOpmt2VWASB6I57GDE7rR9ndBJpCoZ7kG5
wCLkvUTcSjVMnd+/foeZ3BsabWZXu7tVgNHIFc4vp4gUYxDM5+N1trwbTfKwhkca
6Gso3TvSFxj6gb5FfAhf9u7qKd755Xf+m5ETQGokPDCgAXQCH7Y7Y/+jZm9pU3Tg
Sd5E1vvK847j7pJCUYABwehhR/vz3H+zQ9RRKoiDdC46ocxWCGBWpxxS9fLZWy9b
XeYNfpiCqs92iwrQrKhoPCLZxoLiqPKPwT+aewMxM3GRRj0rPvyeXE29onoWvKTa
tHXYThtG9YXpfsd4yGnHGiIHftB1pDyx1NJ67l7ORAC91moJ4rUVT9R0M+a1q4JZ
4X0mE2t3IHp+aTGLFvFUj3DmAodY15zwk2BYX/QNgpCUGyz4SgRXu/w7oLqmR37T
vk82+RUzMsQUQ+lESI+ovuSbDZci3ewPxVJJrZtj7VtHhkahg4WcCiuuHSu9folS
xlxJMOoTWVo3HCQ+FtXZT9axJZ91g9mO9ftFsXcvA2tA0cazwldRjRKeQbyPBiJN
/HZaTMB6bH9yebo+U2TPycWl6DXp/Tkg0bShLVQotWabISoK99VKV4yiwG0lVajY
ErtXNciKB3vW4nAQw0xDwBYqyvpKXUcgIOgAGKXdlxjmsVU7L9Ls2IiTWbvX+OcX
MymEF7DCb2r7aGMpg1kSAqH6s4eOtuvB7UtVB6gtktzDBtqersElbDAhwGE4H9zz
1DoPA/IfmRmS/EAYjOFMZ2RhbZ1vNqiSt0WqqDwsEewNnlBPJbLJOGl9TWoBShTE
PNmoahCPAkrZ4x56L6dqaTGDZ+b5CyxSmyK8pm59HmVk8cgiHSOfxywWdjDyPQGd
CWWhUnRgW+fAvkZ948s89ubWIKPzSOebKt+O8T3RSkX3VdCL5dWmSPZ6IQcuLJz8
18yzzrTlHhW++n2rPUtOuCvOv11TcmNpWK9DKIQb4/GFMU8X+H536kPLfzUguWMM
wr/lQHEevgoQnFK3As40k2xixCPsCQNdhRV1RP9cEHj0jPkEF7Re7r+xhTSwNcLa
BYqqNmW7eF2RMz1in8+FDBgStJwcza7x2SGA7p3XbGQ+ZT5NIilfu2N4KQTu0hwe
csfRaRQX6MymxOIu5axZq7MQKtFdvjqsuWpoHOAhvFsxYWr0UjDcHxZsrZWOZmJG
ymPD3+p/PtliQ3OyCdb2AzpmFxO/TIpbkoz2T9PQzqMj9YtrQLANTkAOOHFwxog4
4Mco+ESNs8oemLRYA/LE4g9inVDL2j7QnA8Eb8ETulUxYpsApU9uGqT2wGAWZQs6
P8LONKnynVKOSyza5+PMBq8mLuWr06TIiFZDXzYKaG2hQ6YV1k60BJhxbIPzD3pq
/ZqLg5tGGj0xeOgZFRQ3KpUUs/XZX9OOZl4Duhu463jHubka4Ii+20GUOlHS8IaE
XA+0ZxqHHP7MdtHTt2G26Fsuf39cWZ05LOqGrFur3PyLoH1E5nu/mYm8b0zq7X+w
nA1+OdJjwpwd/Xlredyssx919jKB2hlYroIbLq2V9DxIYgh9fTN/nO29MUo89NDr
qSZ+OJzfyDWKDVV6/nTD26hbwTAYHBc4/WozqK87oWsPo5KVKL6HD6jJ/porz9nq
7iCiUoNskHUt1Re2H4nN4vHzBt2NrafpPr4WSpKipN3F/yqyiAAZ/6/zIXkizyH/
vqdnTdYRG9a1rLUgpQsFvnzVCdPKeOSJLbUWCJMARIll6FmGMKsh7DC183ipXGhH
8I5dvH4YQKilAzUAbPag6JF354LNY3c6JWVaBDZuZC8WVlNiDIXI87lCjoC33JcD
/3a7DcVqkbkoAnKbXaZ0KLbUuqx7Fn76Wwy4eQAcz8g4IR814zlldmiXEJ5S9rIZ
G//Tjd1x7EXR4WxVZoj+l2i+v94HLJc2dLqmA8y1Xv76uynkCRyn6ytgOJnJc5Fg
XW9zYeT39niqfqIpQnYLgH3aHJhPWzB5nLKbxtZVHbvpzN/pbVUgi3DBAlHe/vVo
eYU1Fe37M6oQIYzaP7sG9/pa0RuHAPG3O3rlzJXOWTu2sBHs8QMRubfFCx8uOF/4
i3p9Ur/JLSiIrVL/OXzOXCqleVkulKJApf1xtBoav0V+0kNaSVBnp/c/N9WucZYM
7+y1e3wkYffDbEq//wcmCLOJsw2ErldaLDDxuEHCMA3Q/NWjJqQLQ1M+bJeGLQy6
tgKOwTdBYruJaGVlEZ7V9Yne/dSk8rlyNB/LDaHlxeMn0EbxeOk1/hcWsk7nuckl
I3K5Ur0iETih1o5nyUlNpKxUcO5vlC3X9ACRUdlYZ46DBgIpywGRCs8Yp2yUcO3H
tPgHtpwdrsZFfus+ZGHnuVolC0T6PRHzn1a4oGWW13PZeOsJb1sMi93EwZNR22da
bYIY/VVBWxPyOBMC7dIeYLBg6i4L8tmsz2iHXHUnoAV7JVqePOrn+ITvnTOiMahb
zl+1CYiIVSa4V8g2BKZ7N1hliuBhCA0nh9+7ZMrB/fLI4+MaQEcvtSQ2XKazIY4z
RFdtoIoJO4dCKCwZfwiZLXelGMlKAgCjCzSvHt6P9WxzUzNfudOTf3a4rbK1wkiS
8EWTPYuxNTpIpZtEwDthDLxGZxS/77tzjH2zpXcr9SBdpCsRnpPMadb5x/WJPdA5
fZZBHHeG/lFs2r5Ng5oH6nFt9JISZq6d9aYR8C7AdmNmqAowb/+AfFjreAMCSVMu
O6u2M4KGpU91RMFwAJlNi7Y4xUexvQATcKjJWTEnn9wSrgL8UNXdI3KEvMGYKpQT
ypAU9m42QUJCiIWhfhbabJlml0a07nQu1c9Dpj5doL6wHgKKZS39hB0JvoQRAB8b
7FLqDT7ewAXeZVoo7VLVTsPyD2v02oZET7vraRN4RoNAmsWw6mOxsO1CrVMUXHHl
v5FLrUrgorE4jPeaClAWUea/QpWjdZVFLbRkPo/lvKqtzzrDGC3n1DfcD9V/xbuf
H+9ETNJbb5sdndXI8yFE0eToGys4uVPfCPBhhNFySa0QOask281yF6pGDNo98vpU
ya545evf4aPcH0IiRYsRSE1yl/tnQ7455g8zno7BzCEjZ3LROr//urBIeHgRnr4P
eH+e4+BOjDecJovsp9aoiQOr1+9ZlQTr2BRv0Z1UOCAvHRBXgDncsDPTHzTHoX20
tQr2minATbGiW061El1oKqujIlMDEb3+AdiQ3jY7VUjxikTR+ufAygK5w2Qd9sL6
zgSIhKetMa6n381T447P6mzgfrlMGUZmdHz+USrWv5Bj3t8WbJr7Lq1d6uc/vhuV
uNg6MdAcFJWqgJFaGaeJJrli4veYppEni3Kmwq1iaXLT/Cj/IJ0hZDZbHEoChNcs
+ANX9ey0mcrkaqOIpOXeRUItwU1S5di51Bl3R9BRtLMkD52gdYoNl39n+fzD0Yq3
lL75pBzXv0ENIjnOZ85yhGRld9NN1hdrUKhs/6NT0HEoNDxeD6UjW7QLfjaKXQj0
nH/IeSFXHfVCVpLOhjEkjgzqjwfy/1J+sZeuc5hmIYAf4Yyz29AXkilPCtRi5cXR
tN2pWljnmyGhvMlf3cnlEjL2IRL27phC3miiFjJHuySXcfw0cGO8L2gZ3rg6LiiH
k2/ZyRQR087cYRCBnvTFAGWwAg3BcixMSLEbzpl2YboUUSpseFaeJg8qB4PIN+PJ
i/hzxyJTnzXkxekEpsWng/R+xJeC9hKGec7y999+pWOylmt14rW8kbRwbhfsC6f0
2Nu5HiXKGEDEgyUdhCJuSdyqUkPjv3Y3F3joUMWqjBgyauc/DmDm+g1Aa1P4Ig0M
tncUHl8maz6B42YjGj1Cx/jtt92kXePaFfKL9A64D+KOLrQhh2KEWfxXoIG3gfT9
dZlxDe166e4gyT/wsr/1w0phKPbjhjmIYY4fuUGyEIS9Nt7nTtKGRqdxBQHfvI4j
C0a3LNl+hSGy9aVEtarZ1wblr1RUYiSsxLVeDpFKxzAXDCntIN3rDIg9K8teMslA
ArCXT6GvKFsVG57cuj1dOUNxVacRQYH53MCntO1wn8T56bzOfLm1PuibB5plVo9m
0eicVnHnb3j9ryMhoFb3okMN5uCCd9A2a18EUFr7kQRPqzviLdkGwk7arYYykSO2
XRx/mb1v5keZCp/DItJqDgbrxsoRzeephuBkubRrdUUCZ15b/Ga3+98GAxCYyLnM
zGT21ZJIzNfbao3jsiAf8Uw11BmeGO5kINhpqLSTokPv1EKf+MTKD1Fq7XrG1jYm
SzmL6xK+ObmfAbFKnh4ZL10wgMlUvI7QSc6xSyU6DadgxjmSS3uHTuCskcyiu27V
hrUWPBZjnqAxzHfImhBCvLPndDo6ev4YCLi+LhtutinBuTh/lEN26SkPP6HvIrTX
s4ZIVGgAMvuDw3wZNRmCXrJPI5qs+6omIC6tnavYpXKGMQS45WQm6RjwhWNie3II
ZFa+PNUNGoR7oFL6tjz4ATzY6qshPXIkPBkgoXPx1Najzegx3TH1bzpckNi0pqui
1aVjlEXQZ49XkBfjBGF6+0vEEvSa5fZKLKTV3CSBxv50L3vGcz180hm/kavxmqVh
SXfbIk4plR4lo8FGpR0kelAp6mlxqAjag2Fd+IERsgkst0ZlwG/V0XRvU/g17xdG
n/cJgQEwywqQtAj3EvPIc87b52zDsq3wGzTEo/jwqNNWRy681JXESysK+LR4fFQD
QFTNxIN/lgtWFiCpjTWNKbMqpfUNZZSDKiN5M5IHWocd45mWKlGJfs3wZM/fNv6C
Tv1hGa5lQEgi/1DzP+N2HuM0uvukIazc1jOst1hskLB/Kvdo7Hvoq474uBxy4/jW
9GWljn4jaWXK3D4T70jX1+x+Am0UKe3BP5UZuhcagQ52TO4B5occg7+FSR0gitXh
wCFISZT5kd5GSFYQz8Td2JhPrDf3kKmNHnaitiPmVB0X+hVAyqsnGTaqfA/8mkBS
nodRtbOxTF61r5RffRJ06Kqj0CS4eLP3UghxGrZojEuWvr7J9yKQK6b1meQuzx1Z
zlI5BjQy2wD4G3oTa+X7DIIlos4xtC4G7TfieC+jI9Bg+2Nj5MoHd04OQik36e5m
YP82UWMir3wPIZspBjmAHSoSiLuyLWpx1wJ58FXrm0q5jft88fx9BiydwvAhztLJ
w5FPxbHQpTevLi879nCfEoeAc/4OXi7XZnRaA/Gs0to8g+X1/IV6VyPOD3ew0gbY
RxFPcAp4LCXntgwZUVfO6830nlO1xQUfqNekCRBT1YiqCox/0tYOvH/WwmLuPWrZ
Xm1XVWKGJtoifYa8TNkbxiZX24zIveYcvdZP2jGzTZ/0aJRbv7C2b0GqDDBi+DSi
SAV00EXDMVbhggOjYE/v3GlA6gWQEZb+pMZiVSpsmsyqAfRt5kXeeu+X0RxcsaTD
8iNeYwxvxp997bDqJ1pBn8BAGN4pTTMwn32nV5YaULzBGskWNDCBSz64d5aGbieg
HoP8I/Gm38wYM8EV6Yma29ZdoW0R9A+W03n1kjctFviwSTlwdvmVQVTmYLcKwshu
XvM+5MTFPb4rnF96Pb8Y57LmtR3kKUc0EcwhLD6iHcearpnZtw3wGRRaL6/Wz13g
zXgIIIHsQErQc6AAlhqci0S9uAJYiGtYM3RczMqf55N7T/ItU6eB1WW/1Igwr3S7
Ftf7iZSO+H1CD02a/Wgho8txTk1COLp4paX39XvPhot32y+mpbwmN8k7hrwklGv0
xtb52DSEO8d0RDZ88JvCjFdk5GywzLgFd6Dgwx0ndjuwjfTWFTEjxCHseSBE1J60
TjTg6ik/OeQGVm8oCoo0XCh4krSMedQp1TtyETNPjfr6PHD1XpI+tKrn66f3ya8U
20JyPqOUUl+4Scq0xRL0goi11D49lFpJBpybzdhmv9rZKOCla7CpZwG1llkwY/ui
NchAULM8UaM0QL/9U5U/ly+BwrWvrXm9biLxgcapGQw3NkHCRtyw3BCZeSVcppYM
nWkaeFX5M+zxvGiODxKaatMjiouIQqV7zXSTKyBHwvkYOGBtw4DeULMh9/YjkEKf
6Pi5EBAR/ATujfpIr2hR5Qb8O19tSEnvZh6zzSlp75t/ciSgCua7SUAAu3vkYpJB
xknpWK/2a5NRrprpmQO9+QehFlgvs+D1WJSdzgR5rDhVFkbPQjgPU6m54pSsAPKt
9jM+Q3ifKSASNhWYb7XjHrTBOOVyxnoS0SccAyamgS0OzmpLr3P/DTf8YlZwjgdf
sSYW2Vj8ZXDzLmhRtP0oDzGSm0ZZAyI/SfpxTg1RiiTeu7YmQ9f+iadjkqLjuoJH
OMih6gJkMUbjExDnFb83Fz/ejg7oXF+oLjLWpwZx+WGgHd5M/GqLTI1RJxXI3wj/
Y60yIsfAM7DFkyLpVHnTGt8dG856Z8QS50CjhmmsTrNX8FTeLh6VWuf/sQFuDbG0
yv0SF8soSVfgIrQeU7PvCp9QbENrBngvzWGudy3qI0JpW/lICZeVmry5yk1eQCCP
EkIl0QeNWWeZ+DxwKu2v8/os3X86eQKaQppbUTaFiFdh2tZUTRKrXyid/rXf0yi1
Qhnu5TmUlRz+TVTJeEE2X0JMJHP3JQLIMtGmQPLTZ0rUw6LDG721C38x4vu4l0fB
QhHhg66EIQGDGTIKnaEGyp+EdbFHg/3ee5tjRH7Vbryb+ILHhOnwmBNbIle8F10A
glAHV5yxnieymrmA4QSmCR8/RxqbtB/evO0sG2avrK2wTVRXF3oFPWnMwowp+NRg
0Vwaeoak6HJ4+KRoTpesu62RvfBpbJBj4TgJatRG4W5/Tye8RS5/xrRJHCZnPT7k
i+ECyp79X40iBnNavcFTCtTRUupmir1KTbIltlG2VtZxCO8o3ttkGA7X7kBCYGPP
IJ1kgyVweDa/poUGTi9rQMZAzpj4HDDvyK9LYMyRxtFmWq3psQ4VXpaWjCN1VYoj
qUhfsCdgxdoJF7N8Eeup/a9YSmmCUaq3xwChwZE61g1BrC+m7sYrd6pWjdkopTo1
7t8yLSL7f7s/kYgA/mSqlUFYqm6E5nDaclgNxZXcCeoGOS8/Of0L0T2KqN2HraOd
5roQB9zJNErN2wRUbOP5jszXUyhoN0C0H5LAUR1sDD3u8OO9okWcl4EAu5Eos+G1
CugCpz6II/CW1dJP1AT5wJx5S5AzXnj95r3/NfAqHfQzbgfGKAeJcUPGUGBNkYqn
mt+ljgG7Vf7KBKvrjsjzSv/kKk6jhX82AMS1OfOsdI5Dh+UYXIl4zJPDnKL6Iha/
0dKkH8PSrK0Q6RhCODJJO2SmX3I44AM3gVyc5Ms0KbP/7jVNmEWtCMWqMvHLy1A1
FKmnb31WAMF6lweT9XacDTbKLoxPlr1nfSOhB1IyfyPhxnZYHZmrNvPr1CxIziYB
ctnA6ugoCOoYV1Sd26sUqj0kFh2gXfyPhhERodCuIp2iEE2zxblcpUBK2hEtfQcM
bi+Y7a5Efi3ZZOfXMH0kzH2/bUb3fmZnWLt83EPBBkruuzPQz/6XCvk+w0p7sAZF
TqvhKaVCMVKF5hMpo8Di6SpDJQihEEWxXhXV6OVEVrtqbd25QQrgrvsJjERl+qP7
sexnk5p2E/HM015ZQThhPxzKVkp3M+rHK2E+ZhpOBj6xW0D0u9Ar37WFky3EOWyQ
9r5mPCAL90xz66IIR49ETVKJ6iZsZyZPcyDsX6TrSt6ksRYyvccUEXBG/XVh5fvI
m904jn24xk87xKBI3t3OLW/Nqz3MMx1QntLQem2eel8wH4kDbY/AoMvylKjZTGYo
9UGTzDib4ocygxCCA/5XoxtnameLkzG2SBhXp7pmMcjJqGl70e7nqeQ0xhmNlEWI
d8XFA7PbIXNfG2siGQu21hb5pyvmxrrw9fj0t6dMgbOF9xTRWEiHgFK/2j4Htb7b
tppW3daHRGnSpgbfo1dRpy5XJAb6utJDjb7BBo7kVCqt19+F+Io7XlHUxHr6DS/Y
jBZayY891ESrbqptHJJWsWGnV+cXgA/u4G4oq7scld3BqJRprPBDnrkzfJzYMpxu
cHg49qV2/dNXnNs3pExy1F1CnewYT4MNvyOJe0KIM6zrmMQq+oP6SOPBXTOOqGO9
5Sb+2H1jTGszBAwb3eE9ZRrED1NLcZeYp5/8NZblpip054vbw6cEnaaaoqShywpF
uz/KP3mCm/JjYpRW44TR3ztp0oG33xlHXBo/z/DnRT1TfVnklaQnjx+1eIhWf/TI
m0ZWQ4x0Q/LBs0i9U2DifrpN4IjaxeEPVu+Qcpcys+iCCLbuFRSmIejuFUUZ8p/L
S+MxgTRM+tOTwjp6TvoxhaCteKY9Q5eZ3kuZNcmwffeVM52uPInBUERcfG3hdlbN
0cQ6vSlcsn84uTyw0UPug5mMy2EugjivNMblm6qyvI/Lf9DhbrQK9C6AfI/Lq0LA
JgzOOoK+stE3nh7pY9gDv1lQHQ3qhrdsB9M30NUeZ5Q4+mT+gV6Yg4Mb/41bxd0J
gcjTX96VSWTRnX99wB2mBV1FTerqPO9oMpZAjKJ6vpBbmCFdj9/JjFrq47lcwo87
EaONk77qMQXRFhFitES9l7KQWJrgFtSCbTdpf5VopzYkPfK8BtvzRVBfcmCMYybX
Z4vZyZCXivFIbhUkmBA2ACNi8msFQD6LXFfmyK8NDeuv8ee0vg06H+fuhhBzAEBy
YaO0AaNOph9i1qiMM4sBJzzdBQDvI2FBtZ5WCU6mGKaq9iwXi67z/vtnPauX0lv3
cAePIqPQxRljGjZCbgsN7YV3p3Uo7xZNbkM7VR4srB9Rccl/V63lwHuc7Qp2yp8I
NMupeYOUGrluJ3ort1NfK0TyFtm7H6mIge8djoe/dmWbRawS+ogqKTgqowsp3s0O
mBvIVlCaQPl55PRAfxD9mnDLY7C/GZfH62NkTqifju6F433afbbllnoyJvEF/TjK
xvTveJsXWBqjbV701ifwOWDNTxWubuztNPBaxAOx/vuHFXt5fRT7+gOHoTvygmmH
BzWlmD3lDGyaLD8coROqL2hVJitC0O1/4p0FdeBPY9TixIvyLmRdxQGEwTVv28Cc
dxiPtthBbVD9XpaAkUxiQq3hVHJ39VlTwGe3hINqdSMQax0YmqH1nXmN+7sSyLUI
CdZo7cLxqEzzQABSa/RoFCAm4+YJArBogmkTXGSnU/dEAjAjkTRcdgpwwd8/HAar
OLk2BleinuRR0sZrHFaXohYjG9XsQstjwsLw00+1nCanPn8nLWIXBC0GMw+6/vJV
rsRd+nRazuWi3eupQwij2qqARYs70mV2wQVeR8PB9Hv0uR0n0aPnlAJpryNOQ6ph
CH1UUJs36SRVCDEQHBaZrurjT2XfSRvRs2XZDorFAYky17xPwBB8WgPxD/hkXKD1
hKMzF6zrfs5z9oBP7RFd23DQzRtQiwRAOOWCwXH1vWZZbCqts5CyDdXRw4Bl2NNw
C4TLJV5M6YJvG3lw3GDaMKMVHnOVf9u0KGrJOmnUVLktie+HD9dVx6p/Ddx+0AlN
z1ChtiJG9quzx/2+oV7XerBFkNN4dVEX78vh27fyJkDAkVJgw5C09ZWe37NdTWPP
Y5MJG1we67gsHjPa4CxZkJ5uCdSSE2NwNX7jlRPvJxLPQoG8XFKJlY1B3q5grHbL
swhn2hGFcnMEysV0tyELfAp+4mDNrbrjH5gzABiOFsflcfUksQKpwZI6Boo+pEki
HCMwc7sb5sA4s8hgpCcsyznOjKwkNUW1EkJ8gDIdmUVvY6MRBewvrfZGC5ilmuP7
15XvVVfdrIQ2DcRPhsZHaD9hiyyXX8ZV4eKHyRIwPooTbNdNiV3k/uiLNQIam/7/
kltyLnPnkzuAtK1Y7kyYtYPbBZBjqViPdEKh0/J6C7jFo9y0VANc+XSTdF8qa+/r
GoWbJiEJvrLHissrVWjZZa91rFcmxpfkKOUaQ6j1GoEeKG7a0cnn6RZdwTakLKW8
+DFmd/3wNOFzjBd0LUVl2lJmZAs1QhQqWGWK/No9hf8ItvCRAICtAzuWpG328YVh
5OUb9laBaxqnAqBCXZwHr4U3C4DOzjJ/NPDXzP6tvNt/eHrd6o1oIE0ZxXbh03S8
PDBu/JNSKWeFlsxs9Da/7zpXWjVha2nTvyrVtAy6ZH/dgI1YXCiLkSflIB9OwXL0
4WqEiPUY9U4g9O3eIn1q/UqCQI3X0AeZhYD0OAbNj9fHKv9002lTXsyiRdWLGi28
pfAmR+u8l02gv1lWXwJrb3WSDAsSaDYXUErX+QSRIL5uXFfGTPiTA0+yRJU+C+0s
qmNABcQ73ntGZYC+LtrK+7ZLQOUruX7CanOluRRMC/Mw6M5GD+s3dGlQBNoy5V9t
sS5MxLlNDqr2ABkreVfIRjvhUaUqHq3fOedKWiv8gyM9SgsO7uBDAIynBFw8hQLE
hvGWiHw604hhRN82c8muom1PqNRHz5z6zownQ8uIZCEsilPaB6WiJYZKrdWGjRIj
vjxCoBok88p5iJUJN1ZKgJUVQiuyFag/RqG/yYnGmXjNXi5v6RGdj83kWEKhHpVN
GMmTwC/OFMttatpJvfvJNM2ziCA/3O6MV1xIhi8I2IQbbBEFVZO1lSM7QsryC8/r
7RXLxY39C6yx227o9zoonlitEo+Ry1231loNgTexQyVmLYWlbPQXmLNJmbUrOGyM
UF2tMgLDcjlz1bmgbSoeLsWkGbgEnCOZ3HETUG5Ehn1u294KTXazRSwRbB1Ueiiy
tpkpYg023s4PXgv+WUWJMPNBeCt+T16ZMLceEnI3thKF9uOt/aQT5SgxyGNDgU8s
wpncf3XV3qwg5MddQwwdLyKZ5va1ElZ0fITvDVthzDrt/LKCK+4d1v5UnRvQFeHf
NwZ2OcH94uU+VJBioqJtwVP2teNm4eWOZSM1LAwlmmcQLjDvvXwCuQMReO4WbV82
tVNuFO5rYRVuZj8x2kDjo891qE0a8qmge+yspsjm6l/AyypcUoU7Y5+Ces16HsNf
zNXopPWimmZYbtNIKwYfMTylKEFB/l7rto3+RI/JCGSd908mVPTO/pqcpx4iv5Tc
UNsGjQ6aXGXLZLV0amHqc7f44DuZIzdyt0+a0pr+/mLbOalSxHePQV4sr8vPpvcG
/ADcNQhhqyf7yvuGA7dOR0so5aZakWLj4xioMScRjIRO7sqQJSGZ4x8Z9FE1CFVC
xWgajt7/Of2uNQwRQcyhuXEA3krTXnJg+1VTE7NkhWnCEpTBXbL8KsTb6YflsFUM
fIFyvgXyQTEUaK4sa5FwHKZBrCnJcTUQeX5wbAIV2pNhQRMk0iCtiyL4fHDxAPLs
7ukxmVx+Sa5XjctfpwNnk8YQRfIlrht037rAOftB2cYMkwcgDjCjZVo9j3fc0xM+
qJb+ijcTIIP12ZFLfFD3u6Q9WWX5bR4sl2pwE3JDAv5rZqjUgJlSwuVfsxrYYJ0e
Lbf4cTnSCi4VKAG2zNo0KGGfh1yzTjfqXkV18e7htacRRmqCNKctFSWTaAPmTZBi
uKpWln41EzGlhB6xPvTqMq7z1m8tXHSqBzMCToVg7Bb3e7GbVDpbTepvPJ5PXkCL
mgQmBHTKI/XTUAt7EbNyjxXSL/drS/FXR+aXny6h/wK/lAKgvyEwbpquWbVC+wdc
Qu6Z/LNWiuIyNZwvPkgRpOGCOQEXWD9SDMX3Uk++uJyLKyqzLpDEGb5gaBVi8ejl
kPx9u5jItOTH5Vr8ENSjZh/yxBwcjjG8tYFcW9iPTmXZzArLOJb0qUFZTVJvBhDk
WfN2JgtwXsDQOr3mUeno21zRuCGWqiEAGQla8PtqVsA0rcEJbFDNau3N5vvLI4lg
47A2220wBApEVdu5hdTvGHCktmnS2LZL8JJSFbvKH649a5RJMiXedlXUduhHvSHm
+XpRFqXffvYpEs665RX3DxkSEcAB60cOqeIIs40diK+r0MC23swi/Vnjxa6dLX8c
Vzmkh6NtFRy+Q3vD3alq7VUOU90rs5JrVqxHi0DtbDWnd34bcr98g2Y0Q34csyzv
tQYxiKaExXZHffR/2CdlKq5CWgL7kz2VCtwOPV18ckz0uknGx+YY+OIlgM3HXbM0
7wdZyMScfyPdtj5sL0RNoXPYqtG1YztQPGRyfonn7goQvnGZWD8edOUDPcKJwJRZ
1H90hYyonht+EL2w9JsuYLsCp8jgyWmd8bVc4BqegrQu1DzgKnNaP8tSR90Q/V33
bBVsZh4Y6pYDNjwpEuKyGbRi9RwwLh0l7AuXYzgH5zaLBvRknx8zX3GR5rfoqdLa
9QkJM+kl9hAbifa1y7btD65fuItwile1n6XCeigoo42RAxbEk5iWybLTNft8TgKq
6Uid8M+N3fcuTiTf1/yupy4AOl/oy0zipmgH+3YE38W0KcORWOdt8yYDt1OX0QXD
4G7uL+bgg0w8Ihm2Pqi3tjKUWn9AtUF0vCfSzLABb4NOPLf6ttBVvYp0ydkKuS0H
EOTQ0+TvuZ4fZohwVYKAE697wdq1Ek/pCvOM1w3v5yGZsv1VVJpHMXfdaFzXWBs8
0yjnckMcnk4sM4I/Hk8SMEvve4xeQ/4/pmMpm3+Q5+0AXl4QIiPW65Vy+6PCCwMk
o+MqCrHK1tH7zJgeNMzUsFeXfOHZkBzX76/8PImm8uGvMz4g+HRSKQylfmkxtSFi
wD5xitqC8E/jt2ACZWOdHoOSqIcecYCwrtcbnjXTkEOb8nWoglwPM2Pm7c6OZS8W
SnQ1YOICy9TQqZaHHFhJkRLBbpTjIFikHRn0yF60SGkbIByLAuPr4yKQ56tABUY4
I9Jekqs3iXh0TcmA9BvH5pfXonsiVEtzlC7VRDWljQPjg2DKF3hlXLv0XOJPLk2Q
Fe3ozUp/9sbaAQRhYK4R2r1k0H2UIrf6IE/mVVcXtpNoXiHmAlMwmFcT0jKG2Jss
W88xPxtfenhAZTpAOCa5crEnoDKJ/AsaGf/UvcYaF4ifnqbftERur1m+JqBq/ClX
bh2L0C8u2JTvcIBm9DD8C15jU9gmmyQcqSjGdBc0Jb8g3CXjFnU2+ZYiYfAY7HQM
w1/9K0qlV/hoNaabeWYQ44o3nVgm0VrjQcZIElcz7B9lbie6sgMvaGu/ViVvctSH
mf5yLJblrPs9OGxi/BguifVKoqzCnJVcLT83vs1E+ZLgMF8r+kOoGpyCUYDIHWZp
EQGMjceraMuSnNwo5/QCfsJc8HcxWwxZLYNGJqkG+PU+mFG7pAnnbq0moCGjj4Zn
AeNHqCB52kckOzHvs1EoN4+YBsWInIexuOErCcYj4Iup/GZxHriz4FaJ8ZcA9UvZ
Bgd+n8bODSTg/E7UyZyxLVMzr6+8muJE1no6kl3yv84SniWZERnscKRPnrDnEjeo
xmwpK1Nt5tBJggT5jfZspiB1tEtthzuVhJ8vDLvr/NA4sbOr6FIKGzxp4x2P1Yyl
a6NO1L08DCatHaVIuj/lFDtkFOaenDzrGtz1Hx+RaAmeUt1PVJ5RVQid72JVhva7
ey1TQ7by0312ihjoz6j8qEtg6HT7alSl44vqxR3dVjc95iSMYG82hdfLBr4ZwjTs
5tqqPV7YY+QBo84JKFGPGOfsC38Q4K7CHeKgxtUwkwE7Nh9e6Cw281xk2QduEhCQ
eIAF909NicTG7sQZkjNjATmOxrwmNhvWHpYHIp18/DDDOGlaVCsKgurV8pVkTruO
OnuaQS9Y/BdA3xMYrWcX1R/ePTgVFstwCrwW9KtaUOwbBc8LFpLzsGZs3ksoaUme
i0U9Zxnu4bd81YZ87AwUHjgwBj1og34buvoQDFecOSahvPsyHgGO0Bl+0FTHiV/Z
4EBIWjOkxjBGkUfAeapNcJh4o70H9Oyr4cz8jHLvoQVRMUsySfbxTJXSkY9phuEL
GVCFsjbZUA943yZr9v9ir9SBZCt5v6IhE6gmRj7v87LyZ5wlQzgajaOBJt3uubou
VVBw+g1r9jH72bGJ/UbNfxtpdZBBZM5Nhp357c2lSokvGwxWzpUBIKafJhiI46Lj
0mXVmFRB267Odq2uDwBfeybD600VAoKmNuVfAyI4cVb5ufhaq80Zbmfdzyejlkp4
+Qu+WUL9StWEbBoeyA3wNPixNh9McDBEa4it5khy+0/ILzBThk1+pP/0L7W1Ak5U
RcIwECgAkRnWX01rOtVU9UEM2Vhh0nnuctyQ//YfWfdrPyhPULzYJKfd5wNHvFbf
x6P/Uut3ZrSJnidu714+QRnJhVRuBVkRxRVkHCpf3k+kvGWDU+z2LjmNZRvwifQe
PJPWQapszxi0dRmtmV3mlB7eVo/3TlwnYkH52BVWyeG/xddl34//tk1LW1ZLYd4I
QfKYfj/RBaecL0KIm29L9NxYC1Vj78l2dA75AihK3h48/3PQmeRuPwSeiW79QSJd
Tcw4rjxAZT6BhwWQPiWUIko+0fK9RhbOugnaR1+fxLGl1zP1DkVcVOVrfwIPLw3d
/OtpX+Kz4JqlBezrYSrMGdfvq0RR8mF/VC8arp36+Js4KfO0BEcr2ESmqU/rVA3D
IXn8MmTEsuY5QiqYl4cglXOU3hrn5bqKC/vJ6SQustvUizY3LxGZLMmFn7QJunlY
8YoigTGrPas+1EmTe93Mv4W1OLoIfqBo245riZmne8TlkQfu5BjpjquOaYpBbF8o
ny7xkSlcNpmJFJaYWDqJnfeeYlAIpxo6PNjpbxMvN/OBFPm7aA/8UEFDFmaf3qhz
gvC/ObMdcbiafO5KH1GblDFw9Qq9Od0aQ/2vPYUKRTjDsUv7sbXDbsN81kGAyLZW
oGHcv1Utoqe8tbKJysq23+zqqfudiEb9MuMDCe+Mdmg7JXeRWinZ//Ujj9CdCbII
wsjT9boOIpuTdW3PnG2m1x+3koRwTJuM9+GytL/jFOsyO98Q6dT8+kQVUwvHnmZJ
uvcE9V4DNH9MZsqSlsCMcbz3HqM+mNfwMNSoGSSSP2u/KVGAsztZnYCW1zNTX6Ao
YvYC4ri6TKCO6SoFhxryohDMGBo3gS+uSzHrWzcNr1w1TtvwPLbxyQfnygaIhftJ
Ur7TJ8kY7IZ0GbCx3DR3BIYYlMuuS4daG6bQz8RYkyT5Akdn4rkDnFrzMs2hA/gf
V0ZrqSMjHDtGgdLB+FlcP5qbvuaaO8BLYE5ejzsiasTKz7kkNPLp/sHNYTComwB8
F7pj3tBXXqfvaCvDhGJuJ2V3IsjsANYDJ/8xdjHt6NYVHiWEk/8sTN0Jy8+WxzaJ
+AiCQrcF+LHjF/WkjY34WGBxIxdQ9wUVz1SaXH59f7dBNuUQeVxG6orsfMD14Kkn
Mhl9Jc+/1wXtU1JGwOi2zc5X0oj18PzRhfMD6285jgSNdIShE911qvjvnvEyBtCM
ZTjFruhXarbvZgEEjMylKtJASBZM+Os4O4S59TrGivdnkS8xI/B4WYIn0wEjFE8F
rsFctJYL4MsYbs+0xc9He5RywcVz4YFTMUs0R0felCzL2iQDJn1bHHnXNtwmVALm
AjvWmW50Wi+6sdJHvIPgFxAgRAqkvl55Ro9BQwwabsqBK+xc7gYTj7iX/Kms8yWa
GZP9k5X1jJii0f2jHT78FMSwoxKeDr6FuTfhxJa/RfUC8YxaaXfX6ZgRQqRpiZwG
3tRmxYAaBONynW4abBXyDOUGwFcyyYI750DYYMJlqgd7c00aOOLq1qYuGBY1Qsnj
/ioVr+3UGHyXJkr8lmqptUPE1FeK+IeJAMs+iTBmnSOCJFh3rD02vrqfTrfOBo1i
fUeft/uDSA51jvq3QCf4qMc/uIr3nBkSdUVjxUONxwjJZHI+QUiTrcMh07pOFtUl
tYiPODmjzsHWAqcRy/6qkIpnh3kM52rWHhspjSjt8iTISDSsvBWr3LciF27KlydV
aOHa45YhOLmsiPb1HDJDK432b96sMI8m84b1B1V0XxPYjeicOiwWU1secD9avy1L
wQY95l3L1OUDInlKpJ0oH/3pBg6HPp6v/HF6eaYfO+KsO8rHDyQLdAgNt1PXjWAE
eSiVxYDcC65YlFFzkcpdRm7vUYcnzILu+0tBMHWjX/0gpNJPyeNVH7tPmx6p+Yxl
NYwmHTl/1rjgb+w3mbCrn3lJBNbJWbUHbw8rGkNtEHZ4eb/J3FAeTVtIzyQ+/SkN
DrHet8C+hOK8F1o9eRJ0gn+1ixGerX/GkTOwdGFTtibJOaG3YOPpdClvpq7Q5BSC
3HJtabOOfMomqdjXSAskDB/RJN020m0ImKf4EV0BYLH1q74ojaY2BbDNzlR6NysD
Wmveq4diVFAOa6ttDVEymKSkNcUQKTcF+bDlcZTzqHi8fPUb/qtvBDCPWriSkku4
HAUub5jcszLBP8x2kRKIUMDM3kIOypmClpSHeg8dj5WxkmYcrNfj168jzsxvZxlj
xYJcYtE27p0bZjs8TD9BzjBRZgaoKfG2m5Jp//Gi4Vv/rKOFkZmxCQtkb88MGJ1Y
5EPtG+YaVn4NDJMsMgFE49zal5B90ypl+iQT7NBH6B+9MyPP2tZjn8nXwpAERKZH
2I8UMxMLMSYbOJeq6El8pRm/r6WzKcW+MQrgW+GFZHd0SC4sxSGg8RmBr7VuHuJM
1zEVwTHqMDPDTrWx2NlxEYCIcB9BBTXtwOPlCgEWo55zsUkfszjauRswMKv4vnCG
BDxiwK0QEQ8zIhr4xf/rF1XxwjlCiUTs1zLe4gcAU+OQdEDrkl/Vww5tQ2SDMSNh
Oc3O3LxRpkLbYvkVtZyCNk8hTTuqAtFL0R1DCgeq0TmHZCxacMzJ7xCKcO6fH61U
6hrnOJ28/AlX1eevxFjqFK6AvZRAV5A75JT4YS08mv5lRwfm+w0gr5uOj1PdiglM
Xa9zdwCnluIASB+orqiVPdmW2EQFZim2DKkBCL6Lk5tY5/HHsu5uH15RwHifi615
zVL/Asye1uF2zKBwL2OabjfqAgHT4BksEm3Bynhyfn7ko90R3EXy35nKfM45H5Wh
zLTr+4y2+Qwx0sl2Zn9UD/kXLUeUXwM0keedokqqutH9d7J5a0dQOz9+eB4uhXqO
JSx/Fpft2Msr0sgIgleubT5geySu4Rh3cV7xvMfZC1Z7pZCmgSKcy/7cr1XPIESi
pToSwHYsRH9sVzES1fU2ns4zSZStVTg0yuwGfgTDM6PuY/ECuGcthCBu2iKjQtaY
82ayoRluWh3kXadeZdrnX/WOs9D1OsCeoRNZSSlB9tuf4sqt5RWq3a4ZWxfRJG9r
Q6CekWcrO0ZJvqZih3DgJQNm9adst0fULsaeWGLghiUgGd6Jb4ZZwERQWpcEOoS6
LON9dGTkaUJ8vMsCDvdlaV90DFa0Wyw3z8RB9dZULQ18OJc8IqY5rxZEKnXvFMBq
Tzq7lBq0nibaYxDqKIWIDb57InGLCrpotRqnrd7af+2Xj8yyYsI5uURACDPcYP69
pfQX3909WYznpIdlX2OKorITYTOMmUqdthe181ClCpvyQOjsX8GFe3DKeqyY7xp/
R2z96EvqSwkgK0COorYNtfZvnG3PkVikHD7z5bxDML2poo4mw+Q3sxVXGO8Mw1O1
en1Ln6wPs8xgUC9qXSQYmx9vYa1TaNwsTxQ+Wm2+1lJDah8ODf+mv4CeNKf7PEgI
XLxh+aDN57laH6EIqFOM7wO30S1CTokZM8luYB0LBXy9dFaa19BhL+WRVCJRzkQe
C8hn/Sus3fBFdxL5bdkAoCcOKBDyKGYhlev81TK56jjq+d03b+avcjakN2rvmJ7A
GCT8vw5xn1sGkttko+cTYtjbviPLyp28nAA3/2c69fIJK/7RJVUw5RsIiZO8VMgp
vMr8x00ry6wLKc8R2mL4xiRlD+PrSPtdKL4E7cmUsm4JwMw9CxCsPddaPJIEGSej
gd93dpYM40HkQn7GC+AF/Cxl7oDtNovakD5nPERncs7u+B0D2uu3aLj0vMxPxmZ1
zw3ekFHf4tt5YG7euSh9NK//FUBlx8fZD3ekEkZYua+yPpMR2r9QTFLJFMrcCco8
MFnNssHFlt6eVoz59UwUc5w9wLein8APme4x/i/KTa4QvuSCWt8yXYDGfoGFQzGQ
gjrYFPPqg76QBp2Y7M+lP92EhJK8pdREucgQtDvKRJZ/yPU1/g9NO5nExbRIkY3K
Exfg5vw/+TtKVioCOOwppx1mzUIWS/eIwigoM09mqtRwoZvHXlSu2rckg5XDLL/I
QZ4j2ulE9kdP3BlcRxFlSf0xIkkxUdCHFtPPKPiGiv/dCrSOagwv1HvbwpIzyJYd
jKM4b2e58dsv4wTIXdaXVlnxnbRRkz17nbeGJOX1GJKzxFzm7p2Rh14ckEcg3Qnu
qDC15rkYemSBuLtS9/mVoWMyhDco6TEF3qtBWwJYumU5WRTJiaeFPH2KtWl+8cYV
jybJBJdirBMpX7J3kRXqreaZbHKY8o2OFxvq5JBciFYY80TfWGX6uCrpKNYDM7au
wwWLUfsPr6eTZVJ+vGd6k6PeTqEc/ye5x+vmAIz2e8gpc0dYXbCJPQE6YSwHVzBd
OLgr1/ZGP3h7K5sC+mTBTRPyKHuFTegjmYIMdxCw7Ql7z5dFWKBoE6XsWQJsAEua
ujbOuLp/wxGpgypdhJEKVWotzLmDDjq0DuArVe5XqavhqMB6b4aUMofqXJxpzveZ
W8drLaor6RRY3CQD2HoWMkt9gelUHfnPnzK+yOLy5282MuTYBry8g91zx7P9vJXp
U/YpmBh74ZYtGEvc0kZgQJBRhPw8U6ljMu47Eqk5pHvxuukUnDytGXJnySNr9rJQ
GGTv/Ke/oG7sLyipFPQKyDiO7JQbi+9HPyRdLgo/1l3twBVGH4ows0p2LUtYVQus
znx8E4VcV7eOAcrjLr8ubSlOUMwBY+XknbWM6jS7p1vN9m0P86jI4WXrqX9pWsMg
b9y5QvsxMQuT7q3/KcFjM1N35mXO8jQDCJfgMu8JPBhXEYhxw2bN8jfxBiWpqCpG
np/POVhPhyIjY6FJLJVSmU6e8aR4mroU0soJffM+bjSscfJl5dq2KZACLqT4+JeL
xNlvMuRFZzaAffkx0GCo1vjy+MzGDHlyhW0Q0yQSwCF8Qr/AH6oe9OxL7p3eqjJ6
1BRRhYQjBxguXLBTJKheFdawOcUZZ2IZxdAyjmGI/X7Kq1PEgzTnluSAPj75BFmR
nt5ZKmpaEAcyTY2sKbEh8OenP7jEoGkuQCWYjwbfETR71lAEstchIV0kshnwNjy/
Hs0MSd5Avii1Xv+4+hEcpk9+ZNVFF7CI4ihm8ZZyPQi/3mQ8GX0uEHU+Z+d83a0G
jeqIUhTh0pdNmUyqkEAPwRFg4IraTSJVCIjEsc/oIorlxkR1kcn5vNYoJWpuIzor
gZBn4CO8UiY7dnQz0hvvh2pBhZqlnyzYiyIgSIoeSyX7yHMm79Qnf1AaT4o9O3WI
pcTDdzYSfGcj4jr8HXFj3QTgT05vxoq5xJLU+cvC9X0+NY7EfoCeMCLUMS8u51DK
OCYQ/BTkMuWtmftB9nAuet0GwoMQ6Ab6nZEfMiNeUvy/qhmOdyX54iTXB3tld1Zp
rk3wB63W6YOHHx1t/cyJs23KKJjBu8tMOqahNwLv6Nlz7E5pO0bmyOdEoLkLc8Rz
dU9B/wZ5VTuVwgGpxMhC3Acr3p8+4zk3u12Cfq48O9yRt5czbbJKV+Sp9k2LpfR6
WDx/aCV/niQv+UIOThacUoBfBgUoS3+YSfhlyuY+Itu3hQrFkruHgIsT4VGdaAmc
9usWtSk3KzwSF1YswHicIf6DwdUVG5LS4dUBgrJJeAqV3wQQ1gAtaYYgMS3BmvC7
qk8GxIg0l0t/Gg0b/sk3pXLRJi/2Zn8tjvVXUnGb7eTAJrPeKHcBIAs0tUBlQba7
q67jDNbMF0owzZB3qFtwc77rZEfRrCmtJd2mldyNyW6Ap3U8acTknbOEkOHlZ2Yk
INuMEH0/Eqnhp75FlejW/u801h43VpjTgNEuo0zDy1dl4SmX8eqjP22APjH2lUta
9jXX7jnOshLo6bAauy1n8J01/sgD2/Iynq64wwK4upEf1QXW3/DzMI0oZAsoFjSe
h04W78Ysb9AdxApSuGokWki+k8mYFPwLEffjv/4DDn6jOzefxajifA4XatjUb/yc
UUH8dneQT1KGE8+2Vs49U482S61Q8gjSHMXw+T8v+AeLd3c9mJV2Tj4smRADavcT
+jMXUy3SSqjdj2Mv7e6O4P2V1xavqWUNkMBZFZiT9S8kFS8EWQwC0Ut3ny68Eico
o1ZPz7SyKjnH24PrlWaClZUjBn6O1EJmoROPo4jk9+n/YEcVpo8PJwlcpgKRQvUN
xKVIQq3uoW+7Jlk4BTaE16kvDgk68XCAFV7KQjnqXQtKCqbTDPf0U3DXObj8rNXN
dpPSCwTintcqOYZO0yDMl/vgpaxzx4uyKld512lOV/skY9zKHwwxmTKcyZNi+eCG
s5MlCag7VQXLBXY7/OC43ujqVUoowPaDGRb+VK1xiKzmh2NCvBhwK2yiVrXQ/VOT
ng78wPzIyNicJicaZ3nYWgHOoKFFEXsFJewW3dPgtZlnyEvTP07tT6yLuiFeXfLc
Tg7jltXhRomu6O08aMS1CyeGyfb7NkJate4dwt7/8iwDuyE1x9Tbh+KxiLfFB2jI
fetcNf2k0n8+GgCnJyIBYbBLX4pB60Xn5PaFPDYfBQ7L3xdq9CHvCD0ZFLP4UUlv
coi8FmynsIVZQ4847wLzKQM2IawZesPtK9uFq4cZqvMPdQb6IsHNg9CrNYdTI8bf
LGUX8lL0GeeZg4rTgL5y65bc/6yyecVUNDqtTbYFnhZZmfeqJChzlJFgTj3wiiDh
Ep2lLOtsKSaFZUmFkjBP6ztLtLViAf+XKRkNFeXpx1nJAx6Owi0zL30GECXL7NgA
WZW7YlpGx4uTrS7inbXDV1P3MVKhmAOyBDU9tLCZZIBRC7DHgz7zpeBhC5raT9AR
lEfR3hInUh2zISXgXFdRVNMxfpOMOA4EM2wANPMZURcUxcZloy3RsiAwWQ5xwCqK
W3ucowT/LzVbcR9A+9eVOhC7mgAsBqsnnQzHmWD+xGKXwSd0xqHozM3ECQtbDLWn
BvjM+pnBynAz3/KVPwNG3sQ4y2VPaQTe2xhpGj9PfT84Dj7lbQVxV0hJlUDLJNXj
WToUwponMudUMTCGAVjRrOONXVrGpyuKDva3205sAL7oZnoH1g9yK60O4XdUsy2l
6PVkpia8QJEa2DltgDtCKsKn0cxmFgDpNbeJsJcC0vKZis8PbQk8UawCfVLwzy6B
fqTGi6luKc3Uw7bzhs6mF4HemJI8mulFIRtEYS9HaxhwCqKwieQdTH6ow7+xzv2J
HTv4FJvE/204rBKRcWt6Nc++MQgzgEwMgpePxauziKmA7tACV2pBrKHjf3pXPTe4
lD/XhPpf7kvLdQIPQnGWwM8zwIENT4TDIe+C2IRROtqleeFfUTIZ6pGYWGB0sMKi
itHLQAXF0jaUdL/s9UG4+vq5+N/AhTkCwj0jYLy8yc/fAtIUh9MDLT6IuIZPn9J+
DkXOedpRd4BVv+A3AmS8jKK0rLrC18gL1cNT/uWrU6AIMbndJZDUFxQ3QlRCO23G
Fo6dt3udTEKkbEYllLDDSR4+/hLZxgXLUKdzo5jEKxZShHXh6yIfdAL77K/NCDUh
SUabjNw4T0w10n0ofW/H8YCPFmkHTHtn9oJSXkwwwHQeBaWLS9KSiDOK7HpqKbFL
ILbJXOJQe2C2obgm9Nc+92a5igmJloioUsc7mbDR9Icu1fryV9UFyFvUrCBcD7Sm
7beZoyQTOBnOCxikTcWEzXrogq9eCH6V6NEqHpHrhhcR893g7ScDHRErAlU3Jz+Z
hI7SV6C4pVNmUMOhotbFRKB6anxd3Y4ogvt/7VvoG/7Vh/6G63xwGToji5HkHreJ
F9Fdo1o4zponbhH+F0PnhtII+Pgbld4n/sNE/o1PruQjiPB51Uour2Xb8wDooduJ
D0Zrkxht/LuKPmvofrAmfZfzpwqZk51zKvA3233R9H9U22qolXSWUlRJ2yy4+bU3
IfK6uaZAjy5zHu3B/pXwCL3Yl+YzmdAqynDUgz6+k0rwTSD1e5hB1n7H/rSfEuAp
F3iXyIbGhJu2ZIog94uJYJqm9umucGThCHwN8gOxkk/HMlKL1wxoPN2IpH3sW4Xo
SqBVKyuHs9NA1A3FSalce1erloqIKYaXXL92OBAMKv3hs+o81tJQJXS5Fb+nLHeq
32Yppkon5Dghta1P/PuoaRXekDEkGa+iDh3TEsuugYcKDc3YKHSkLExfuYS9r+hx
9MCx/g9MBLZUbFN/w17bojYskZ5/Yv6SFfZR7U+AA76QUgR5iC05e88PFsblWOuF
Di+RAK7nr+5lQCaPbiNEctlzloloByE98lgDMoV7jc8T8vxd4vXJHbNndDiQMiU+
YcdwmrQ9aTnRayUyQF6a+GZGPKtslC75DiqCSArG2GRMLnI47i7Rj3vK12R2T2VP
3UBIkm7H8iugvq9vic7du/bmRBduFaOj2ZZvNODiL9E2DFRC8Hcf64E7EsULFTdD
HPPZ/o1XqkzI94a+dCTuX9eGeZLVkK0FwYuqJUF3IF+VLX0n14t2HNUJJs0skfkV
GoP26suA5Hj3chZZZ5x9RmtbEowuKcXU7/b4jswnNon4LTvNK68cW9rYstodSUsM
BVRH0hrEXpoWEjHo5KrT7zEf671w9B2x1Aw2z91FDMpVtfpqrMewuvZ+Yr3UE8xp
BV/uwhYXghw6rY9NIWe168C6cTxsqh0f39BIBIjbBx+5oDn9wwx7ton8c3XGsjip
IqZC0wcVjehzwPsKMaeN7BPLZOZCH+3sASX5rFIYS/qgzsMU3F7ym6JB7j5F2yQv
mGQd0KcIxI9Pc3LFhLV4d51o9sobha7yewpnu0bgcLMGTM8TCx0HsH/tWQs7eTvJ
vglBcsOb+lZeTOKTGHr7o1sYvSs9bRIJXYv8blBUWiNln+BLcEVlJzQwxG1YiTjg
RFjKF84as6z0eTAMJlPilmz46S5150awVL8GLWgHFbYjp7gai25R1Q8zHRM5J3kb
1AR+vsNtnebsa6MjoJM2eGk9ietJ1eWIB1DZoPW92g/NrmoR0XDQaShJvBKeRuRv
Vr5755CT0NsN2mvA8fM4uDzCHVuWpRDRCQ/mYwW9vL2cBI5fe9H1YpAO1J+snALt
e8WPwcIfYXCjbYjbxNCBW1jL22sXAr/daJ6IrvNGea291tw578AXt48zfC6uE9bq
NJAgW+2nqcnOn1lcyu/KrMOGjZllf4o1FKOYekIkrd/Cxwwakp5FkmPPWrFFOiCX
59jGO/JB5qQIRJglWsaTYmdbXuDtYOwj3BQJy2nJ5jpKv1QlSYFr9DfnI8qjtTxv
RbWJ2Bf0sRh13D1HJeL7SV6MvzG6LRFng2Vcg+8wZyqPCZzI99/vRadSQpDKcDWF
VnFN0TU5gd39WCAOwlLSsYgeBeTLwn6UxR3OHjExn9vfldfhuGdUkTWVgiJCXK+2
rbf9PYJTrhOyAKCAW5miMONdkeEldPRNrtxWmkm2L1LcVDCJhLvYZW2WvNSB+0SF
QLckZOIs4hStTD9iKDLevOP0w5427T7ldMPoGn+zsECV4337GobmqHbztbijhBEk
clVrJ1A0P6ASsTezsQwUrUu+crhl2nW6IgUnF1nm11lGLuWy+yGCSfQ86EfbHCpQ
iQCFctyYeU9i8OEOYsaMsecwOVMW8u9YxMwIncf2pKTcXB241nyR5+/CcT2HR+RZ
V13Qtrzey7utQKIs99ta7LJ85JFP70P3Hu9xF2FKYaHKqUSTcvX6NtOKEG06eMPp
Wy91+V3QPg/WfhoX5FleEY4hC7szE1vA9+FI6aWKqXu90DRrIc54WlTN9L6bFeA/
10SRlUvtt2oFnyIIu8dNX9ZeEWvTm/HrheJIrOGL6sSGkkppArER4CHST7oCSsJG
vdgRA8A7bboXwlIWu7ivOWgqYQbDcT7jRJwkgUZ15SeTmQAgNZ89Tg4PObH3st11
ZYo617CJBna38UWTZLKEytSwiTDZq7Gt8ffW0TF84FSC0ki65Sao09xKHIzpDJEB
FxnfG/EYdczTG9+rl3LjU2Qe6f/zBNPRBq9mKe9uSF/5Mcibq56pX7XwOkYeQgRZ
6lcoPMuzCGYNWqeLW88lPhZktOCZ1xj6SaWq3fsQC1aZQJlpp7D7G8k5pZ6MfDTQ
6E62E76COWnIpYFVgJ1yQI98R+pje0grmNJ1tzguySrLs5FUykUb4QWETfVDudLf
AeE76lZFA+11tjd0Bcf7bY3rLBZkut8eXdcW/WCmOmPDzrTqB68MBl/gdqkwY+xL
lfMUjBzGT6UQPrtQ89iukLbdUsIjMQx2ErVtO8LekKI05nULvSo6c8Pda5uBcoKC
C5XQX3wNVKdAfnzCB2/wDlblSZjeuxyzfG/zw15+pXcHgaHVJIw7RBjWlAWCcFUP
iXjdpJxAsdGgD1RHfnc2r/vnViXkXSR/2EqcOLxegYW+xOumgl1vrTRKE77jcI8X
EgBRFKz9bbPPwt1PZelD1tOQKZJqumoDk+Xa0G7ja6yqHYgYToBk/NdFHihkybzV
sSza8F1gqWe/sZ/IAO2xpMiprEglXWktmmC+oQ3SwYB7AowC0QFTiTPY+uTRTvOe
GgUUKiz+3LABFoT5Maewo5qnGdu3rhSHglhT3NFJCKBOu8g4KYVs5hqvN3cTxPeV
jzU1fSQ3SANeewFT3JWYWXIYIoy9nEHotYHxKZXTAjETOTYTL4jqydMjGZPA8imb
3D3veAqKNbc/YLiKQJVemsIv8g8EcSwar75Ri1oAQAylZ2u4Tw14ZomKGcjnXPSf
gS4BvLQ1hBYS+WNSFYSbppbwKbRwlNGJba7Zhk7T/bMfNqTZkTB8SJ1qOnbU9xUq
7DaxLSEbK9j63qwoiEg6ZX1C7kI5uRSiUa49oWFnYRd726Vdh/Rk3cXVKk8npB53
bKhDyQwV63tWFmdeEXYAkI2cUbZB7Yat7mXuMwkFLzhET7IGEzYvw9MGe15bo8kv
MMCR/zv7gf79CesCPESNw1xYqdjs2pJBqROZl4aSbJ8OL+M+wgjmBFdFHZEgfpqw
rY2Ym7Cxffazu7paTI1EDpIAexPpGbgf32+7FuYRR7FAxp4VYgslJJZWy6IRpjJw
OKcMmlTPQ81kFnFVw8NZY+lFp9puSDRfpmsHcGogeV6o6Vqxgdrc/AYSFLlrR/m/
d4UK5riq3jMu4GJEhQWEjynj4gWbzzZPM+e71d8gWX6PC4j24kbfIEhyH42/yFUS
zCTM6qK2n7RB+lQWF0y+SrynoFjhJ2aiPrA+jk/2E2uFA3XQZi1HkT6u5m8jc6uX
B47KTVtbrQwQW6j7HYtEU39y55xDawCJ0gWKCYFVTXw9DNvmrCVRy+LbmDq8n0VI
KJvc3yPGHkBVh56PU9MqRrbiiWM45bx01NzCUYi/gGrlUOFXQR/Kj0cuopGkDfHk
SFRjLzwCHDOLjHc2AgnyDOz6BZjRWEMlrLTjeIPy57FZEsDOug/pZ1v/9tjlD9rW
KCLQ2sV9cs8W2mRKk0klgFMzEhuRkliRDt6/N9bkJbWjuQk91Pz1EjJwcgs93n4W
Bjx9fBMN7ajWMUapJb6zbpUOmZifxQXPaJ0KnJG6PaT2Eim+4vQ652vzCbd0MkX4
uqyVzrHx6C85CRKmHy60X1hp1obBtcUxa7xm1k7Azm/neZKjkdLJnw/Wy4CGy9GQ
FUd0g8a9OmaNYAMuUUsDUnoD42NefymtN1HXIM+uWvsKIELosNfmuezBC4UmMr56
o/feKRCWa3+I7oiGuptQRAHGajZKylVEAhXNt2aFH2pr7B3+RYURvgVR1zO3YL0i
ODg1lJKblDgCDYNCFazL79+LXa4qA7ru5KxNgUb16CBBNkPM+1QaZfSQo4HUfraK
lLvcy2Wov1nYG27yKwJUOCrw5vAEXcPjjO/VZ7cMaErMtFKs+n2VQRJrYQ/LtmzI
LROG+focJs/7PcnzqPeX/luGZWm/8xjo4HTG3GAjHdIspY9+2bLWspox1iS3VZWW
YQ13Is01pf0KIDmlWIUart4YLQueS/quWBEM/fsBZBNDGNYN0h76vt3Ig42yBXv7
078pRRuRDNyKhyl4yIWi6IGu3wSSomjIlo7qfs/xZuNqItxSXx6U6G12wNa9FeVe
5wIdx5JtnrW4Whm9jiGZwu7kdpmXOB2c/Cwvq/M8RpTPMPQoBxELa/6CfEUOmddC
9BkUTQ2v9D1IwAOGeWdW0dKtMnsUo1MPbVGOei9ENqmC+Rmq+Z+CG4EYgivivckW
/KtnPm0zvuoCmKGHao4uOQli5k+nORJu7C/YSr7fDq/XrBD63CBAAAc23zZYiXh2
y9WDJTFmmFARF2GWsY2HV7EZrlQTn4uojmoueQbQpOPmMd5ukb91bDAd1pM1iQIn
dsrBtdcUP7A+7NJ5myYOQMT3+wEENrWS1uGVzX++xYxOJj97j9/mN8fE6xoLpao/
9ItdrkfTrYWizsnkygtHFz7zZnPShixMkSTd3SALr2WDK45Bfakes+ZeiQL02CK+
scd2FDsbG40RTvctUJ802YApg55M6uxO9yfds0CS6UiI2YL4kQyEOFyhJT1ky3SG
FxHZTAM17lEZYq0D4TaqVyal1nyIIcLWTMT3nPjLbfpC9XESJsv99NKD197LmR93
JBJhDHiVBUmPZJC5GsIafgXBglxVY004zxr57ysE6dFHomaOF8D69b9X6fodhGob
xBrWHkaTmx9sWJyShGBXbXyN0LVnzImFSaRfxeQWlZ88JPy84DTt7bsPpPasel8c
SFB6lpvw4F1Xq8PgNNVAwecGheKFPMm1YziX+FhFkd/LJgt15XHeNDAtLywqdvj5
skXAg0x301Nmv724HmTHdHtzcOYZZ1XKIVJTjQ2avF5Y+NQFWVYBCrn1JKYpt031
5dLrlN7BUh9pXfpvCG/PeVRBf59dnWUoXFbKbr4QhxpLjx0TjMaM6QJY1+nQOAJp
ctzfG1YPk3ywsj3c14IHodbPxw41XmkM+a37c38QpdnnwhUabcPHDGNPK7eVoQ1H
tuYwgP1Z0YhFh0+63VeIpQ==
`pragma protect end_protected
