// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:09 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KOF4VwQ7bwEtzkOU2FZNwrEHRAitY45SKhwVLASNIiM3wJc40gXmMaC+F5A/fsf+
2Bp4qOVkxKy+KQXyOHoOc7HSudU9Y4epnifucfasJGTThZ4ezxkdih1YuhMSMCvO
UiGxuzWXSN9G/rK54+GiCJMHi5DOwqARecbAJZlIBuo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3792)
Ny/uLJsnWbUjiMpyPN4DtxAyXrbjikXxM7TbOgIjySqO/8wEECZljmtqbjhZfR67
79Ossi6ynCFyK05UhU3o+JshUrrnhLs5NGH0xGkB89w6xUm8MObXl8nM5IBbNwL0
Vk/mwAjOhBl+al3NfyfzPtwNR9103zopABzxKHcy23D9sC0Jhiuch9O93B2PtTrd
tjPpxf9hGspCT1pHB7gB2gtnTioOGB0uzBcSWi+TQ2y699eAWMnndUxjhHXXsVYE
V48aEzN3DBBeaQgLLpDtzFMZ2VH8MJOGCrrAu6zpIspLAZNRS2KKeSsylru5FIRr
u9/0yCgxjFJwDI3LN25rz2PKJcjJtS1tKCv/zBhEZ5oJv3/m+B46tH3tG6PD4L8e
35BuSxEtEpNirxbVjfQzevi320f6QtJdMPfr/jHUGcHs6aX8t5IbjgUGUYoIkxNx
gyqx7Kuj1pqBMxfsS1zL27t5t03krNWFzHjQ4BJFIoHS1NLBCVC2W4rjBoBWtlIZ
czBZF6PjaTP6lgchQIXFlhAMAAJjB8mDNXzi5FEEG7jvF9loY2JkPksljVSLzDkn
8IBvK3X8+cjRCOkTXgQzjTBIclSIU+QkLeQnB7cDnCFaHGiB8cOnz/IufOK3AI6m
o3zug1J12YACKRoTa54bWt1TKSpoNKQvc1chu7/gRZYe+y2CuOhdw0Stoy0RK7me
t1WUO4v6L+iG8TpoyRJ7eQ4Sw+3PYTvXTjjO0EJmtnauQNDOKbYsWkWJ0LKEHaXI
x0Qj/zaIOxwnzIGqMz/qRWd4sEu3xJMtD1bW4SvwLWxsq2xkXI0HszEJsZe7WNkf
j8E6fGMFo4QFyYjYgwrP3RuKagcBDXE8z4BWYV3CPWsqn5wdmaEkz4JTud07/0ow
HaGI17ehQpurxGdAVsb0bW/4VmHcVs2So0eGcZBaZdXqfCH1lPvDmGSjXeUUTZ8L
ceAvx2cVgvvNpd5bA008+sllrhXmE0S2l1nnXJCzv3VuCz46jJwlOqCY+DMXYrh9
Eesi1NsUuxL/bNJMTw4Bv2Dc1Pf0hv5avZBHvpK9bSGv9Ic7Fygao0MfSHYZl9wr
XR4Edq27tNEcWa8QG4s+amtB0SUUmz/1IbWnZZdN0okLg10tPeGGgN1bARA9r5o/
m8qDTmaqASSwVU4hPCR9lDTNVq+no60ibuotRe70wHiCeFJFzysveQqrqj6UseXK
jgNioOMkgeYrfWLwglH42pQOickArBIaUHR57lgUmpwnfX9VLEAMvJXNXU89H1sY
Yh7+sMPI8P7B/WSNzWtai3kZW8nWUgkY9bpnzP/djKB76/VaR/YHJ92SrU4ChxP9
+oOsuycv4uF7WrvIYf4e4l0fjPwbgWMOmpO+fTwV4d1h1ervUO4Ijb5Qvl/2gTn4
k9+1PnBbF/BvQE98JkBsTNjerQmmkG413wAjv43Bb22Zu9vt8oXj5D4NIDViZtbx
6yc/fAgR0kqw/4a441xeTdtm7MvmWu+Vgzx/wqy9+P7TqNblt6U8hk0nywK9Thit
y8zx94qavdKGu0cTvhiaDaKmLjRYyfhdxZFhnuVSTO5wxCS1CwvmVe9QudWvf5DE
wC1Hg7QbL9ZQjVbnz0SHbL4IpqoQvNofZmOn+z1BG4KLyRWhizED2/HWPAwn9AzA
D0FvuYWqbNQPBvLncaEMrPQuHdMxq7OQu5LT2RyO7p1R3MihOlFL+BMUbaRvFKSz
Y+BG6OtVUYUt5av9usFtxllRTH7rn8h3uU6KWlU0NMUYHfsw0COIhwOd9aqplLA/
iQhXwzIp3e+LUA9hARQJUhdQQfQSBgPfaIZznAWtaWSmKyQSJjiuG/iAv0dDXJnN
zj34WZvLPG6uAbUmYFgxhig3+vnnUPU8foUiZxymQJ2yvH73AP5UVNUgxsn6ltZU
fzMido3OeKD8uzOKeEgyRe5UbASdeJ/nn0oMweuoRBOmODQF0Hza3n/4QuUBONU0
Nzi3NLUeccIUYSXP5uXK9Uff7ro/5iNv2GF5JX6HgEoc3MfmMxQo5oruhwk0SjE0
umNxxZ2QV32B7jRyEqGNgEjE3xanxbwDxJ3Qb19L5oQpTpvLPoMRz1VulIfib8q+
SxnXyulgH2GZHSNnZDRJH25DAS/gK5WMM4WDQmuK+RW4ZHn2neiEvSILmslH/Zb5
lXCMcXlhWtDQvdUUUuTv5nu+PB8Ix7hRXO/CE+3Y6Ws/FH8BglIybPITktIIf8/e
+M/rHvSECFrIFoN/cPwZD75RulBg1MbJv7IFGHWf/J+VRDmjVe7NCTQKgjsN4w8K
ke5/PTkuYnp0KRnTCpOAXHNYz/k4nIbUdYXh9o3Adft8inlDxRrFA9UvxkLWKGPB
p6y3+Jz+8UHp+ME4Z8cnXmrikNnWVRRc64dMMHYM2CiUXYh5o18LdkDpnEQU7gN1
wE7h/2bWYL1k+TCXXpA75bc8S5DIfHasjzkfpOrDW/LDMVtzEvWIBftanWvNyXPF
i293IiF7udF7MAgO4w9M46SjOe7bIjdMllVljNCclnjGv7VABEwCLLxDTbZfzRdH
s+NBu/gDU0V6+3EPmGIgf0HjoKfYIuC7R4jFIZpw8m31CNVP4esON1FxuDjnw6pr
JLZRuVgDYbT055XOm2xdU/VLd68/vmpewoSPOM02h+ofXU5bdqFSOLmfBVhz9GeY
A0XOPrtnyW7r2JqSk0nqw+NjnYG/lpqWf/piVS5Q8BXEcLlQj0SBZtCM+aYr6H1L
Vlff62UXGV5k2ejnqG9eA1YZKOYOaxymmsuiujl671RH/MlasQruKiBICjT5ixgC
TJgng5CX2idWIsSJpgZRKPMA55oTdUKZ9ogMen20l8lFbwReb2+xn+dKN2tX24th
F5YFJk6vBHFZwy/00klMENXUlPaSHAE69jGAdhv49JLU6ZBlarmEaktqX4F4YyjV
Kq9cJWCAJHw1BfaLjDColXaUJGxlH8w7g7K0o7Ap6DQhlNwhunTFnbtmDxhDn/Yf
RNrLPI7vl2bdNvj8e7i4IM2B+k0pUn55rmDqclXKhg2MBxPe5+2rfjrwi06S35dQ
iv1JmpADZyofy+KHHujR/MUO0nVw4yjL4JML5b6iysi3iI5iqLXDr+uDtpaYxOYl
C4Za5T5CCHssBbskYieHnKh5QiR6Tr60aTion8bXJnQ6QV1rjTRk5Z7ke8wlb9q0
BsQi3FHeOpxx+mxCWUDjTkkQJGwEHVgWMnttUCf8t3LTxH8ag6YLyAoZ8iNMruHS
l4qGsVOl+T3/90hIAY8UisT6jb0xKM3trzmtI9u20o10dWlRTQNZSztu13nBzZIR
t3OVxbVh6sCgTqycaJjwThZnorZirkGy8mg1j3mg/MpY6eMhPBtIkL+YaDb2xQ2x
tPEd78bJHQQaKl8zu+PCiG/EdPY8ucgVlMDMsJb2F4LnODVzNb5mpVqx/jkBdNXB
2XUBm2hthI54jt3JIxATq5R9iCZBnAo4p7LvwA6KE5wVn8K/+NKgvYIRdp/SvB2a
4noyRMwnzDb3YbDFnj6JFd+XMv8/OMVwYxThv4UFm1T/6B5zD+2yY7BmMHOdln5H
sYS+4e9fW4g2oimpVnQ/3ihkhMbXHI3vKuoCwiB8vZ6cVWezuWM0JD1CgjkdLkse
oNag/Xo+ybjD6gBRhwMYAJZvCwleHx0SMqQE1G6vyiIooOOtJAidfKvGVcs2GdKa
x5MYtG1m70xqUzQaSBSozEld3rQG+PS59L6zuItzxEBdSYo/26JdawfHuUKHU8z9
iXr6Un0cZIirF0TFq54yf8/VRTOXtUq4vOjJNYUyRSW+9/qExGDDp7rhQ2KZnOfD
V5meCxOgHG+mJL0XFGDw3ff0gzxZci8LNGdRZxQ80caeNr7kwKts/hiUGjIyfTZn
HXpl5cLaMwmG0cGNYbsBcl2dNnJ+JP+EBPIkokPSlrtnE2hqnfVi1mUpIVVFDazQ
Ch78ol9tVnnIOqdQ9ybu7ewVvZPr8pF9qOiWG/0CmxCH23tE3qmj8xwEXsxFFfJ0
lW/rc5GI/fVuCqPhbwe8ll6GeLeecvfzNq/1urDSEarLrDV/1mYLspEYV7lC5crM
bAKpbeSeTRa3aSJ78KF6DnIoYnbkc38HCSvmmgCoOj5LTVJX5hC51WGMSET7IUph
K1NVk7aoSx9HFvZXnS0iR3BWuzFw4gyHiPF0UqVyDnh7N+nBB1EEPAwLo2D2tMqn
Z3j+eTzveyKVI45U7Sv6SJRB+uaUqCX9aqj4jeYsSURwJKvsCS2rnVdeKCISCysq
fKBEC4luSH67qCtxNpwsoNs6uyLq48xqfk4ZYTdhjQdCDae2Fq0sgZFev1IinW+F
M0oCs4cQEhkuVFhY+8JS7Zz70uLHNHQGl+rR2O5JBGHAv6/6kqDL75eDNyl9wPeP
pj+1sm3A5Cxci0Ga0vJ1IDR2oj/9xDAY8bAjjdAZ4qhmyanWAr2BSDdXFT6PX4Ug
52Qr2At8Nuodcz+GQTsMP8QSt2eIWqRbwKtQXBt/xpdvMjfnZCfAiRVfMcLAsUL8
tZ2Bsy5eJREQ8Wj/2PjtEl+GdrFv/UB3IqXbrnKsMGjPE7Hq0aEtM/kvQvvBLrNn
MEgQmxYwgc1qBxqlI25VpLrHun1L4RvU8ydbfmXpkRlnL2lnGkuK17xA7nVA0g+k
BV9RraQlkxy61R4/QLsN6LeJy/pdY+zqGDwpfe5XWYs5p7bdNaItyo9j54ij156L
Hikzub/QUR3zA4ht94A/3AO56PV3Y4JZXBNNgzEgk9nqWuzuqje/hK/5ROHb+5Rc
v7XeFcfSYt/I2ObRj0MbA3OcSRLJt+4t3kI2sp+EFXGQBY2gk3Fh+Tgxk0Y31Al7
WDmcPA2hb6pcsL4fYGLuZ5lbDz08VHaSdjVSWxV9alYmiUCdjvVojIXxX/8e6tY3
K0nzenC5Q9jwc3O9DgmgUM6/KB/TAjMWoaf4fTHLbVckxKdX2qsvifgHj/rDZ2CG
IXNvp7fi/xRTv/xN4awUSpY3FnzCMhLwtUXfl0I2R/JS3pkwi1EhDyzZy2LZ2MN/
`pragma protect end_protected
