// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:12 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ltVFu6nHrYgcMaWUN1WmAe6lZDuiZ3HNdvtY8ZHhA1Oh8vXxnGUxULQwKNVMTkBG
F5Pl87a2OyO+/xm08SYCYzM+OPSUJoQM2iUOV7GPArmoxNZ3Ct174QZ9CZbpZ9Z7
Ovpx09Tq5URObPc8RbNj9juYR7Qh2BrE11esrQp+alY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3040)
ywq/9USBqIj3QnNKNs0PdPeFYPJO4yyq7y6OwuaK07qLkENGqUiu8RyiriEWp3BV
0u3vUht3BEnngsuYnI8VPSyYQ97slAyD2ebTCc6NN1FP/VxBW523sbmCR3QMv72y
1T/jh1zIWj+COd+XVWjj6szzz1QelP7pawGF3RZF1yJNbJG5Vmy8gKk9BfvIMp6y
yLcS7MQ9Aiw7tWL6GoJQqyrLSF9y54v6ZWzs5YFGDPoGQthN93v3MP2sZdOglgah
lZUpC+cuzba9FfA8Gg9oi71AxGKGdIOnuQ5O5AUmzP47IrmVMKduDLJoOBv4UiwJ
I2XTKCWhGih07kqbh0ZEqpPnJ9mW2mk+9FF2/IfoxlrzNQ+qGN0Mb7d8Kkil6imB
B2A92Z/gf5HmhHopUcxQB7sWqq66vdhHl/DTZYIPHDGman6Zw36QCNlvdv+GBl7d
kXR58W1A4e2VDYQ/mJkI2W72HRXG+FOOzrRtgzxFrmWXboknjxs9/262IdfFlqMF
xofHJZuO63VDXggK3zDrGjgbmxGSuW2TEdA0s1cdVGejhboBf6tLJPllRm+cCNU5
jcnCnIVc3aa72HOQLkRZlqzE2UFloNFn093o/f6na1lvKf38agfbZsWxovEYXu7h
XEy7uoNmIKZPxE6NdFM86uIkeUAHm0yy4sBddvpI3NXk5wE2rNDcTxUx9FEKXS3i
GqW+0rcnbQUu6Ua8THOiECETRfDX+Tu9YtfOUhqzb+akuS27QGf/9B/4UCi4sodY
HRNSV8CzgdSIkIulzWlPSNYz0NwOjSfE9200WUJ6IN2cJRiEoT0zD+Gd+JpkT+9q
t/PQ0WVSw56dxHa0s4jnpWQ89CTE/F13ARPeXCRg29EH0TncctN9UE6gMCV/AbC4
zoyT2rnoTzHEMUXNwovjk/fzcEUZ8cdDzCCJvXs5doXFO5ga0fGyihi+sD/6Rf8p
5P39h9Y9NnVA+xjBqmjM9ZDOcwdX5dOLNv1Qo34BmpKDGC4L+Di98NoQw0bKz9QS
DOl4Zhxez00nshBH2scDokC+oMT6k2z/saKcg31uy2E2Z4bKF7dWTKe3KT/MscF1
KE5a0DJw7U5Oz/Lpl3Pe5ouxXUEWt3O+e4Gb2RPl9gOGL4RGaJVM7dYSDnHqoMoD
7Knbh9av3Ll/1lvy/g81gz6N7EAgV7+Kcmjd7WzHuX3+o1xImPGF8Lys2e8/rxa6
6/OgzRi/MHNvniRHr09x+ekd3GcwsSEFZLNc5wVoJSx8nltK2vV4vUcfWRXcidmI
v6MonY2Te7Llmxhcc0FN6RmnQUx42hrGUKDpG+g5rETQjQpJVCnVmlPJ9V3ASbZX
zNRE7azxe5PSc/UY8PrhPvyevqial0hga6O8vzlagI3fDrGZMj8TEEqpobbk48s4
pNkOCHfzZeVQHEC3H3gH7U9wyYLNSSNwRm1N/VMYvIhHPPOX8YT/Oxxhq5NhoGL8
AaHZeUmcIhIEMsxP91Qg4HyjUhSlCIKFduxLxVXR0cqbgQgAXeSxDi8FTvy3a0aJ
mJsYV/17rD07B6zSB9Q84UFS1N7oSWYvoEiJ++EJAZM8HjOwfRuCITwBwBl/XQLf
zLOjfMf6Ldz86d/7rnnJIRGOZzvaXoLvhINfRqkcWNR+UpXt7dJL4+IKCm9twFe2
OzVJD4YKCi0i5elAtwwmb89R9UHitlELYSYLCAJMtnHEItW7rwFaG4146lU3TU67
9EykhZhul5MeqPNwyugQZ44n/LOSuQErQai0fHHl9/gqPZFkeGwuZUQz8MjhIMTK
SoiP9duJlNSCQIuyZ7q1nn7+53rWLOdt97iI3oRbc7ixn6pW2RZGMjYtkZMBMwDg
wEui8Ee9WLwJNperGZU7qmp1zU0sIZ1Je+0sKhbdsSnQoM9d3gydZG3H5M6PzT9h
7gqTzuzcLGoKm2zfJsMv05Dvb0B6nUPPBXs+jqdKKS9xBcaWuImBijlaEFSJdQd/
aqeQSjLGpbFq1+jMfzphN7jnIOPukS1YR7UBC+1yUfv0ErBu/Gp8JmE473Q1SIJ0
3MucBR+9cb0CTtiE/dgtxJJL/Sbq+g4o06p3mE4B0YtbO0gn6sP6/d3nBfzss+uL
ac/EjOeayp5ymbM6e/2g67wNXRsw7oDZH923X7zXZJStvqI9welXeFYbbgrAjeWE
P/OYjpKgYeBkGhG6NWB0VHZW0X6C2ep2E+ABCP8cpB4A3VpltRL6GhhbCmKxJ8xM
L1MnqtYBCdRhy2VEl1E5hCc1fQ3kAPqRmwRKWdXxw0GeBxNvL0fzsQSQ5+PNUC89
vRmA/yNWVdErWl6sPEIVEAFNvjFItsoqPtt436H4K7Jak34bSW/RE8Nb+W9BIjiA
j/rCiQzZWBIclvMaR5FK1PUpfNQcPi8ch5XfgfjqbNeA+J8YGyXru1CerKvPpsGp
F27PJc1zCLpF4L0PnQAJl7tatMJR/GsSngRvQd/9MFydVNu1xWN+e2w+J9BxRsHz
/E5CnqqLIlUZGBOo0q+hmTUEJ4abNdfaGmum2tuSaKiExRja8IqE+6I5hBvwFsMd
Gs1jwnrgvGjmS1F4shUv9KOx7b5Qa9aF7A50BGMBBQy9/NHeo47+0t97cV53Lyzo
aD+7hr9zEvIsL+f/EwPBjBiPcKfA4PvQrraNj5fK9TIftZR8/uz7Qgah1JVtgK2e
SvlYR8q0GPPBcZIyB1QjqLDgn2QQfpZGMFoeSRL1fI2s/MHefpNX0qaNAMwQGqR9
yrZCKPm1wqfpuSSW1AZaaG00VwFeJoSaP6f5UTx90PCh7/VU2+rumEd2RWAqqD8R
SzIhcj+M4vcRF/ungJwxNmCPwKWFsubqyZPe00aN9f1rohREeHdzPNxqnwtUCVrC
FL6/LbF+Ww9VIX78UPXGgypPNnCHz4d1NXzwLV/cqHtsE4FvFLo/hEtbDYgB1ibe
/j/BnENnZH6rearrLJpHnIp9qBiTIwLN303LmasAY2BcRzD6kS95GumPLHHtQ7kr
6IVNR+JqCvULPXv6UPiEdfo/2DjSXq3C/f7KoPLLVPCv8jqUuQAEYs4yUbJ6S8Bj
2MXPtUs6pOXgd817F/NiF1lpDc7RdUJyODEUIPHr3xlSq+kq/V2O8KNb8+Jlpk1d
MjfYwcsr4ZmFWSb+hmkyHcSauz23Fan9PQKIaRj1VCl6gYelO0tdQrg+Nad7vpmc
tvK/6S9FpNRUiCKYxZuZsFogBnXwyFPHHSDWJDp4zQxKgd0kiRJ4XugPpLel2Y48
+eCqvtQYoqCtIIkeN0sbYNb4TG7Wfa5Y428CFgIb1p6/BYC0vEvLtlj/DmUGlg2w
sM0AcP8G687+J+pG4TpWVtOW9ctU/jmuls48H1mhcf7zLpUmJH+V+gKZ/JfUr/9R
w8X//eJ9VYzU/NC0PUxAtV7HEhbr3WJdn3vY6NfsIZFF5jtFmsDyqX9/m350tgpE
G/oQWpnqTKefcNLGQsncW/kCkGDzdJc8snf2HJ0inJ/CNm1XhGnwjhSa9MffFSL5
lS40+rVllhKZxYYswo/sFgdgiRVEUxjGxZr18dx4Wb06V5NYKYv94WcIKumd2gcl
va9D90hGzXsmSvW7igvgbsOpMTGVyytD+hqng2Fzs76ewi1xy9tLK3tyE5T8voHE
F8LH2RXop+bZQDaouCffNdZ2Wcgtq0pmOfLVi9t/izerXvTgDh0dC6JEcL3nxsiC
Qsw/sVTLY7CseAVbyvAc3LTKhGn4e67iy4pswG4JVsF6mrRbQ6IdGeBRLOgIMPcX
DszU1aIeROuywbocrQSddlYtf00GtBKvgH3BJLU0gGUpQ/EQTPpnhn4n5GbtR4B8
MM3ifcxSwKIE93J+wExggLhXzPyyrlDbUO8asI34tz8Af0xRdn0VHPW/lqbTay7g
iqF647dx97Mddw12qPzEv9IsLL0fgYw0hDBbxn3hlplKWPSCHO+m4DUpL9jfyY54
+arhHtKlD7V5a6CScf663CFkZa8DochLxb2hfHIBsiI+38xh9iO65e0xgaLVyUmH
6WnffKEQrqFl86pXp+QGSQ==
`pragma protect end_protected
