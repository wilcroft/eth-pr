// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:13 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
B1puM6BrjxqFruLTmiuf0FYMhR5MPWEbn7bZwzrjdyCqDu8FpCbWZq3hPavbfYEX
bqQXhOgE2dTTOg2z6A9ZpRB23fhRPpK53qiTBe4vfAiBfJCzk8ci+sdAdx3Rhn9P
giAHYxcH8+hcVjtsqgGTY/ZpEeGQLoUszZn0RR1jROY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25872)
3POQFHWKuem1OS1uP3dlWyepAJ8x/UCgw5lgADzAa4eDvc1Lh+uiyGdIv3RF0yAK
3ac6zK5JNdgLFJx93zEE45pGudSEBSTT2x8AfVEDhyXjhZ7DLsBswKo/p7uPQSWs
Y84z7TulEDPWAW2wQouI3IzBtvgq1+j4+E31VNtUedVrWLBEEPHuIFbEQQ61RPXM
/1zRqqPAKNEePNAcq9ao6svJVenqGbC0cddK2Rb2EG3puAt7qC6s35KMFvyxRfW2
WoZ4P+a/m5J6IPrQcKQijcGhgB2HGOtT7FjpRjN/bWmbsEW/136Le+//TBOtt4oE
CDsBCiwzTrP3Ek9alwGkb5asloUby7NzEe5vstmJA7u2hwDbxa6gQl+5hpArRv/5
W6run26pegBmJNzT/XcJqCLwyjs53FCime9ayNukGU2bmQeJMJxK7o0vS+sw4PN9
DHNueZKcGxwClyrN0SaoLp8jlJfjqrsKUef5REAb0vbPsdbPY/RnQfesnyYGMbhf
ZoDr4+paVqUWUdXj9m8LEKQel3xEVWqbiBv2jGsXl7W5A7lW+zypE3jQkWzD3dkz
YwRLTLAqZhvc0CfzA3iELBiFtC+xjryBIhtUiI50lA2j7GwJ3b97gwr5Hd0DeDZ3
03VN/j8SS9GosJlpHes/o0lwE2s28Swcswn7ALK215y2jq3EHDBlI2kRF48Sg6rr
B0kNqtbc/JjqmwtRcuGc56gM3XxWBguMFzYAALaq7QBd9jQYBMOX/wyEOy5A/bf7
o6DDzLjo196QSttjAINJePHwY/7PTVHNeiBjhMuprD75mjqWpUIgiN+g/0yUQplX
451YyhH05TcICeo9azluIqN8jnVSdKez2RQE8A5Zote22DnOIckGWDJQERFPrnVx
AdtPLHonIKVBUoQakSWJ9c+N3ODtpCk+akDAKZ9HvGmW7JozR0KE0C715f90C3Mk
rkK6pp69Z1wuf0gluQyynO/GvSwEHq1AQG/9Hh6MEm2K6PBPfcXBSBwpsf9bcMpf
1xopPbJw8/T9My58pJC1J8OgzkBwe57JcXTbDA5sl6VuyB/Vn90SzdB8kdOFoZwe
HY7VHhpXaKVfNTv2Z1mSxc/tlrgdY0gk/9pmA9kTgZru6RZ3fWvwl/znfWjdhlJB
7NFNo4GKGGGESpcYeEbWxFVzl6TjkK1Ng+oULRhOtquQF6sxQ42YjLcGyhIyuKTR
QFa+nEAJ0jizBzHcYs5xqgsYwUS/os5ev6EkCN5y+WfI2FEMqohB6KuOZUHslAJk
HJPJccwidfra9dPXPHX7vJWKBtrFs9Eub5TNy2/WUt1Vm/hw21ZR39I21+QEJ/z8
2dLKSwKD4jHsEyvs6wmZk5EiKuDx4xazIEcD/wq8eGd3Rexx5mQ7oW5QAcTvyd3r
bgvH+DwNSx7SPQXrEYfYafwVqCIkPFq6oDe3lic3kPZuOFmE0lpwYOZDFYWH+5Tn
L6zkAI0mJnmaYUUKADhPPFw6P4ne9tDfy09YffUC3ZODhycGYdj6F7OjxE5yl4To
y6oWKyNf6FNlYga/7Em3f6CMDu+fIZWw5FqMy1BGQIkpsa3t1a6WbMIXQGIvR9IP
R9rljkGn7mxAp+3R77sQLRGX3dDcIOSXOrQocNfpB07SENkxz0/5Xr+BLBW+rtkh
WjwD5VjWo4D+k/baPG0tMzVC6Z5ARizU4YjjBjskLyI9fSxgf4b052j4DS+H8Zh2
pCrjNJlNx4iqajZ0zUdURglIWIbrhLI6Bd3I9+vkcQdRTsjTR8Sv6lJk5QmGDg1p
OaXiMmPJoK6aQVeQDa9Mnsad1Dj+F3mz7NlvxL1ABOn4cBKv7fhpYt923ZB3aPby
4wrTLEf0bxmStZa/Vf/r76UiM+xQ7rTJOtRBmEqfux65dP62ELwoSpzaoWKWk5Jb
5ZagyjZ5lS+2Q9gwjWkyToBT2AW2s+dR25THBEaNlFcQWYPCVsm9TlM/XwVVdyoU
9vCPGlMXXpeEaCBKcU6X0a61bwHAIxOvGXFptEtoTscIdNh8tI0BN6ZuYqew2m8w
9HeFYmHdxB0jNXMCk252CDF8MVarzhg41Ef1PQ1WoJ8/6jnFsptqMXnuOdsQa/bA
MKKKZ2h9DfPD9dbrmQRfxJoJ5T5OtrlqqaMeRJTrOrKmtXUbagqA05Fp2UaDH5i+
1HH9wXtMal5Jwkh8Kx7O8ZZJS2U7w4OO5zQtD5oO9tBRlWwXwi7ZCiLEL2zgitnV
txTPAcM7/XG5Aomu0X5bg+clDuIprjdshRfd4+BzbaX5HkHFQ9wN0cnAbrxlx5oM
YuuWb/CH6pPUKqnWdBY33zOxxs3EZbdtdG4OtABk+PqSf4BkWY1zz52xKU9uXF8g
26+IPUPEMVHbDqaJ97Ac4c2sdTP+XzuCxecVK9JoAuwWE5hD/WwzioY70ohyggZq
VKD3R80E5D0HYLRk9fIf2cwhy16e3JTdokLKm1OeNtCOHICRODvP+Wy6BBIQ6UHN
cvhofJyi/u2vvByeMNAQokF3JEhFy2ZzMzgRnBVaFCM5yO7RdDgSzLOoVX3CPl1y
nlXGL1VzrpBDOXcftd2RmFQ8w5TNCC28+Cqdn/1W8CXhLA7bTHBtCdab0n7awORr
Ln6V7RD3oKdMCCRO+y9u+ixywIW9Y49GwzI2Nh0CDTTooIJAnWa52ZMhUoLvlPfV
ZWuApuU5Uj7sMWYe4R1S/ZTv4fFbuB76X5bc+HqjP3dcl5x/RgWcMrG1qXkjQZv4
CLTZ5dlSFuG8KRnrjiw+lotM7hBk6lF+1bQeKwRemLjjLySx/UvEPg15wC3up6y8
78cBBeHe6hVULTrUFBrUOgnb0a6jJkwhpI+JAtJTdXxlBjjkFyRS/P1m8cyHd6/+
cCHj4g8yNoTHpCbZlpTY4327l+tiz1WdKsgNMbHmu+NwmCNGtbS8TCbjYC0yyvsU
If9hbDNXPsE2MhIdJsKkAAJJmV1vLeS+tGPuuCze+eF36AC7BtjPea6kLSQvnAcw
GwPPEON1lpFPEpxxWQVsrJJEaS/qkALlidw7j+tFYlXd1BTmJpCvg9LTqCpkRsWk
7SuW9J1h2fV8wZvwudour7Juyj8FNkvhLeZcwlJF6uleqeoBTDTrnIh5vztxacbf
ZxoP71mAJP7RAzDG9yUg8u95TMZjxsQIvZiNN+lK+m7fu7lUqb+PtOyAqAFeylPB
iGhLyS7itD4oLWRtdJtSAC0ATbonpWg+jANhkS4yjvjYfntyWA3vC6AsC7rlXLHD
19rW0ALALysQifSm2nl+bA3mimmC0qt36yf4lpQUtyxB7WNqArnjeFbEmA8Yxz4J
qqoIFxuzmZAKmLj5XrQ/HW6SzwIiXxB0PJd5gimWThrBjRkcP5mZnYQfUEg9dcZz
yNybQ/VHOhO45OfgD5Y/XqIB2wAUYR3o7bZlUtTRHfaqgO1kXqhK7lkfB5/xis25
cMjmZKDrAzagKTKRdx1ykdezS8aH7EcuJ5rlTRsKU1/yETi2KMVeseIOwjDUsrl4
1zFxnFLhDtefbyEBYlo/0YLlZ2SefkhVsxf+/Nwner9nO1/Ti/EBfCr8Cm+3MyfF
wurAy2Y8K+vQCytbifidiuGA/bMlyue/wMy02bOAvaADQSgUZDJx0RS/FWAChSGC
Sl1lVeMLvM+Nly/pbhlDklnJSsYkyV38I/WUA21PKN7jGqfzsvGrbwWJqxJsaHiE
t2uXkCnHcc+jL5Pn3qdg//7eFWl0juVAPPlq61CaFjXaYG5plMZ6o76E5EH9TUlg
dQFRE6vw14CSRLaHycvRzPOAp7r7Gae4rSZ0KhcHBs6B5qqFANukJ6Vnmr1S3RB8
874BYgwqaW3kqAzkLP1LMa4AJPgRc+bnow0dCwR1QoBGOcbodvgRkphxQ2HWxsLk
EoKx5w0WhsD4Qd7h1Kd0PuzD1XlnuZkmY8LLti22uZxvjV19bOR05WASeXWeqz5W
w8RAE7bN4jd8jPYlFOAOZHo4nGNxC30bZaD9whTBINCYCeqhnFI2Xs3ACXWEjGTh
2OGRT5MYs4HTQyTDEUxZbnLklNP/gxEWcYIgAAwcYb6zOkJ+7sGSKAN5akNGR4eU
Ux118GSM3efZeEg0nXrIe2E5ORf54qvODAA8Vg3y7fqOCASHcoSpAC7aA6311Q7Y
W86WldMY8wYOSQ7T1gBlc8jtDeV7EYHS8qPrkR2Mlo3ENm/sbBTq+PIzEdvjmPeW
z0gwy/pwQ3Qi3E35KgTwvHsSHO8y7165pcgkfTQT98B/NbVtcGxKR2V1k6TD7z8D
mHigIX76W0pypOI5ltyZLONg4nUNzQ6kqWMOuDR505PScDKjeX6+f/Q+RAj8Oh5r
4OzlEULwTnSoqPE7AH3OexWTSmNYJ3i1DUAteqX/oN4uaKR07mpbZAO2VAJ2IvlX
pF7S+e0Vj2sksu9biJFW9ttZLJePcOGu37S7ojMtXEjL2+ygH034ddu+Ex7uIKJy
PdOY/bupWNy5vLA+aBuzuf+SI7krMUbarmPasxSeqXcInhjWOn/Fs5GJtFEqb+uW
lYuC72GQYiOzycYP8m9BVLqHueRY2FY/tggccJeSTcM9jJdCvB+/kFtpg67Av6Sq
pQtjNgSKlugKhRMGrI3Yp439XsoAU+11r/xr0Rp+yGfy39zi+/C8XgXO5iMjVUky
ba/yhEPeOR30Twe6gt3Ch22Nl/WEAaqT7WhP9/1+KYtEcaHRIdHh32ne5JIX/2Bg
KcYNmGHpBCPtRPVEJDLifgQ5iF9iSGb5j0eaFNLL92mxyemC6ylOEMEjyifM0H83
0rx9efn/vGzWJurf0LXPhgrSCfdCRGgVtWMkwiaUm/ktDWt+X0+6KLyt50rb0MMg
tkeGXdzUkQi7JOMjo+qfimCsojjiYHenNvN684VeLWiVpyS8SZh7ZbdsUgki0911
I6pw0kKM3SCYSEwwMdZFkSfNMz+++WrEYZrLsPKR1cWAuyABv1FjNxnsAMQYnRDS
esxzh5Umb+KuDr186nfEeNIZfYPfxfoAvwG5Bapqxcc+q5wIZUe0EtKEMa2V5/Ma
5jO2G1sMXtKXwGIfAbrwEsh+arxCu3UxrliU7esc3fOUx9BIfwpSNF/iXcV0xyyc
meQ2Y06RAzNATnX/I/VWBTpjiXqh5Gfauk879GeZNHPWbFypMCjJT/qAF8S6jo45
/69ab8VPrOm17463MAM7E+yBgM7bCRtknkiPCyu3cvICWEBKolTF+teZ1eQ1Gkjt
I3FrhgUG/vOw3qtqevv3gzxJFMg/lDGodQsNc+oslkzVjPcWttR+33yWeq0QLoYb
DJEMrJEM2X6Rb7qwBGSH/SAnctKml08RDVxgbaQq2iN1r9wp24akNz0OInPLFPXp
HuWUqqTE+9Pkml5T9RDDPRozoISwwgzwEDEQ8mi9/9zY9RsYUu4fKlc5wJcHj8s5
zdl8fiHUHs8IuSN7KMdSlSSuVBik/JVDarz2OJ7e/U0b4U6GVpBApHDKyEtgXWmn
z9E2/9UVCqU5SIo3ramK7GaDouJcMCuxJyjdLJUHsNMUICITibdkOwLp8m8PZ/iq
77LOfIQoJI6IrSxKX/31yIwGWGAqNoJg8v8H/s4QKndOdhsp3/kpK1brtZAhqnxR
gduCZp9NJqrH5iaG2DiKjzPcZKM1rV9r/vEJdlSJCJqbmAuuwYvnuK3rVUA2oqZv
SfobGPRWujiVsZMO1PJn4FYn4yCOeMp6Ch2IwTqvxe3CAz/8skmfZx9CB9ftVqaG
YHycYiRfyZ2dVmnJcvy6enxmwrkqGxUrkDQRDk/9QLhIbGffbm+rDkZEi6Q3gqMf
eyPSl3cp8i/0NR7JlpWqJ0rmpTngBDGLenfzhI6mcwjF3c/LeILaxUJVrirS3RKV
mrojlLUwViQPLBIY0eeEM7Kw8J7TrMR3t0WbofnAo+UnkdFFju1bkAhh1Hqyb/17
zT47KDqCLLc7C7P/A+pJSmiDtYW8Mfg1AeZNvNJNYZtlus3A4g17kgDx+b7sh8LQ
IB/enxw2o3toGQarhhZ1O3hHpLGGKTQlxlfp9ZYiDVq4i1YZNm9grfvNLeSDh3G4
fhfjK84uzXtpcZJRFX0wWVF0rKn2o7Q3PAA/XkuxEGWZq1PW7n83AhvOBjkYMWo/
sovpJ8idxus03b4ojQxA8biJhfXo5/1VLAIU3MeWz3NmNmp5+s2e1xBrfqbFWtaH
UW73oPQO3U0dECoGlwzPIpwvyYI/RMHsbvideNpQpgR4ybFKAdcMsUtZhl8Mdknp
+SNwIclUmi6BK0kygGBI9NkGxIikbf1o7KQ2EnsEi6QDRZx+G7PwxAs51h3oVmMN
RPnLDuMC72kzzzWO4z6mTpeNJHjvgHHOf6h7a6hH51vAuIUOGt+9ho40VMH8Brcz
l1HgrlgSbVy4QhvFa4F2KSRmAvYinworxaMPXoKgiBR0jsToxuZpClgvamyx7RAI
LWlcw9DT8nuh/dpCg3oA0VwETFcliyo09nQ8drD+yoMLrjT6fpuKPxNxWsHe4iJI
dGQ1Xf5E2Ndvl/gxBJzP/7HlH2+UMFQxa2hHzKT+ngYFrFy4HQDimW16QTs9QI81
OQfn0pm6fmySra57HBDmh4Rr0SGWhUbb1iHs+6HHQf6lBPJT+o0QSb4d+E8YT8oD
F+dWD/q2ZHtqeqB6BJ7yAmIJZsIQFVcZ3SU+19u66GpreeOg7+V6uoN2fUGgabMe
ftPoFrytxlBhuyWDgzTP8dzgmrnDW9o9ZmXQq7Ak9ISZ6/DBWmuAEFkfQHbz5lL6
0qV78316dyAG9KuKUxuD9ChVgu+BiAhUrJLlhYGR2nvRaZkhJwNyXNtYpN5lN7S+
fwV1Jb07vzeromE7PpZUXuqCJETNWdpRfCja451qbun1o2jdWExnZRA0lWK96m6O
Ewj4RB2KmlgBe89fRB3i6imi0tAVwtBNPscLXcqEhNFsRcitGUpYn/CxNPINnTxi
MjSdV15YAvBwwtSo7ZwCGT1TIGE51yUAYniYKqxOihL7qvZZv4wFvE1JSAV0HJ/f
x+nHPU7OxpK5FJJGHrC5bTAzWcJnOCsiqAjnWxdiNIUTIPTL7tYXwZ04UeM3JLX9
g8XvS6AjvTCovkexxkJQxMN210erlcRp4bcqackmaix2j4MhqiNy0iwVvGGXKSyq
YQ10vGCvYkq+0DxTDMUWRbLslWCYy6VycP0q5prEi+WLR6FVr/yk5N7UD/tspDb2
UI5WerLHKQmdhvBp/tgybxvfvKxFP6+IIiR61QqEhvguWezWYJF/MPNTiuXdz12z
akPP8pQzqCJSQMlkMkxXIWmhWATcB/8Ml10ONqcCJC4jmwxgl8P2kSBm887Z3PIR
JYfUf73nCr0xo8ewQNty6ZhdGD1PTlaZrOefuEu3G5hvs1bwMnbUd1gXzywUi5vT
x2beRVCYlvlBNnQsGldddzCGGmZJBPpLgHCbydl+0VMOEGhek0l7h6H8upa7jeo0
5jjl7HaXCfdSAXWlrEt2lTMkZFysPwKANcd3CRZUQgswXYwfq52JS9RCUt+SBm3i
73cq7ITwf8Z83VzCUTVlyDinpOavYHzlSiAr0UF08JpVmKqr7OS1tNc+u63P+lm9
GyY/JuEWq8omuqHeBJRsbEwy2gK6il+99vkmvUSANHmVbhgtKGlyZFJ3wbfoZU1m
PzPXy/fGDMqC/Og6IiLfhMN8S5LP9p854AfCiPo/Z2RHF7/pGoROAYhtuB+p7Mw8
KEwnXvdb7pEKWW4F6svr1q61rAmBt5Vba1DFtjPSQA6PUwXbV38vJ1bE7B3Ybc+0
yRMKa859cx/FuNKneNrEKw7kE/kXmJllVkC5CTjvDj9IG1sJJP/8Xbv0BgATsYd2
HBRCsz0yAdc56SD1PcOg8sJxmcXc//j3l7NFZr+relD/SKCLPbVXtmEBUleX843p
OwfG2a8TiR0V/gJyqSiLptW7BZmnxvEbvcnmEQJGKziOPoJoDEO8nHHZ0za9Ylce
21c7lXBQ4qcxoUgbO6vkY/ySrZFB3vvFxMtMQ+QxpzMvSC43CbzxReBPNHV1pbGs
0wXjnMocf6qBkZO8ZZKYkUZrhlq4PuyYxwSn0RcSnA2bhLabYXA9G9ZT7JJRK1Ox
XbxVuVI8EEFa8SZxHFbiKWh7jxgkVwWS2pJ4ghAUEYneTB8tnUZAkwiB2Ptb0sC2
oIMROYkKjiNrd/g0AZnQ1PlXVtC+024fhobK4BW8kvgdyeZAsjzkwU4cifn9Y5qh
ZxB2w4VzBqwo+yK7BXWDZN/Q/4mjo6lQmu+IaVqHmUQPJcv49UpOuWkUZX84unAO
Nrhi2c2BYBaVFTimOHDjtqkEAyTZoEMdPnuQSZOkZMBN1AcZz7vb5Vd4/2WPfdgE
vbxXRKFK9XPpzA3jPVgJlYDblCmpJvwQT5UNIVhERKSkerhP4ypE+e8Xn4qipDgu
4FXeXz/dEgQU92quz3H8HaiKIVx0cvj5S1iWJZauaK8/z/lPtdprvNdvF5dZJHYS
1n8osXyFikCC6whunTf3StjS/quFnVjAWde2j2oR9WQeSugf6UkuGX6rG74ltoFd
jKgqILjsOxTnUPH+Wcwl/sNhXTUxg2No8IbYSS0sJ3oTXZ2/0ddq/nUQRwnlDEx+
h7imDQ3S1mhPSq/KGNqQaHGv8Gq0JKERrmXMUd3l7gHtc4nNg+Wcf2E/a0ZVslXG
WZtm7AX+wloz5nCUMSeWxFDLE/9S6qmMEKj3TXyLQWzSucBUO5UlO1o8kXbtaM7R
hnABXg5Z6HI4jwTvmL1lfm5m+ujQK1Fe7DkLb862jUy+MR/hrGO670yg0r0gy3fd
+DQdGNYsteOs4w9uLp7MDNbUEb6w+HiD0QzdG6djiHZk+GekjyXqrS+kAbWYTTsP
RVzzSXv7VSJSu4BIt3ulXmT0MR+n0T5XhjNRchUDASyzY6u4k/3+t5uDZB2/h30P
81uNvdYz/KuJ/m8u2VA6CUCtySSyM2ECIojpK5diQpLzqrM8+vquyqPEdo61apM4
o7cKAHa1kxeNU8+S3BhPoFeY8D1u/fwxEJmQXd3P9iDn7I2HCnXvCGj2SuK+glfQ
PbuMGnf8K1Sk8p2nGYSxCN1Z84bLqFHMJHUQrsyeVmKvW2ML96t3rFRRwluVtQhS
NZugYug7sUAeD7hfahCYSrZSGcOMa1ElAytWuziZabAgo5NhKUem5G/XxYNNhHhW
dAWkL6ZqG5ccNZ3OH+De58Io5OxBVxpGBZ941kJob+RUiygeOb7CWTWdckW1APN2
zu8wPD+Im0kSsRaIMfA+21wYyTfXkDGGLU1qQKc5GHXynx5dc7syB8TSA+gcC4I2
lOGZt8Oynb3aRjL9cLAPcKSEq0H2cd1fGRfwDsVQfaiORVoDvtlSoJkZsNvxoc2F
wwNnO3z8WYv/MMBE3O72xlDbF1guVe65vr3I5exuNjO1/p/anmir9I2PDIpAdlkW
mdqPVsuevmBOT6vWsxpCJ7yRrKUymBmlCZl8Itm1hMZFNElUog2fau4urEhMOyAw
WrHFI7v0eDGP3Z3QQ67juLP2kCRxLYR2cNyNTnPpKvbn85zGDdGCvxVP3G49f+tC
l2Ls+riEoBQWEckaWNwQuZEvl6JN7W68jV2ZwOGyxJc6HJf7qVzL5DZ+6MUJ/Eid
JX1Pnk/X/Fe1z9AyYFaWOA9kT7sfDHkijTwstXka8VRcGgOWcp3z4Zk2am6362pC
t9ig2ZNjfrnVt+TLoVXofFeAkH3g4jSDYP4es/uTOFX+ePAx8W+xMhWzZ5Z/DJTP
r8Nl4F/0Hb+QgETfo7GSmvYLP6QQmbr6mQWpsAGCjEK1hLfxX62pgBMVuQktZnvQ
SzNXqi4PCkf07gzjnbmDVCwU71UlQ1699OLN/SolE6QM9IXC9M2c1kSnU079Lds7
tGx66Ok67lOKGsgetL14/rJUT2m9dpDYivL/gqQG8p88rqSnhMDAFD4KEewfTFcz
dUkNyF9HgV8mA5Jpxu6Dz5G0LBlnj8G9pq1KFyHCkG2HiruaiPqM857LNCj4Wvjh
EFwAqqKR70NJa5cQxsJKdgdgJDeYhuyCpeg6EEh49Cew9PIbWnpsLSdhw17/LCoH
TfdP3yyPNNejCZbCLZZ0YoPLAIvLeJWCwJRkKE25XI0lusEwfSAsXjtVsxreowfV
cbxQZQ3sY/uyRD6NfCrlGaP7oOCSzCdx9TIyb6xehZtofgGGj2Ev05rBi0QicitP
XnFxrjvd9PKO23WGNaGamlmlrv7rNNo0d2mz2TkfjIPoP1auvQc+HCMcG0w9yneM
Jqd9gP0BkvKs4PDoC3bOJN4LDG5pX/GKgMUA5HDXaVQ5gVI69WFFKauA4ex9LneO
pUQuqvFTMAV9KfCtKJU0iqUlDyWpaUkL1vM5jvU+rzDmynh1qHoDNUqi3TuglupP
AZwyNN1g/fF6nqKqeT57jwzO8jhsms9MAxI4+thCfl75RK2XS/my1zV0B/ThbxQ9
rQ/RMDe4bNGLtoXUtdtWbZoJFQMTVmKuVZ88Sc3jeIuGoCslh6RCrBVpczzosGk3
dI9IQxwiZqFx7npU9IM9Htk/kQO31nUQZOhqG07tA+407zWn+tUHCALN/QK5/+6E
sAzWRf6UTypzmSwP1nZdh9tvGQusu7PqjBMbRT50xAgwNOr6G9+nYzOaOOiJvmnI
GSpRDE3wL+Kzw63tfruhFsuluwbT8dS902EvKlKFzLm1ron+M4NGqNs0jUqPGufC
cF6GLrgfjOvn7bx8TVJfcgHWtq2/WKdjgTYrVbLpLKL8Z44NAxOqDqcsJYuLpMQo
bvpHWxzjRYR2pVCClIDJFBbdlmyn+n3M17+UXfdl78kjODXraXw8CBDS6cUB+v6o
bmRR+i5NMBrSTTC/N6AjZrD2CIJ2g9POyW0jDtzw4MIHKRNGp5eusA7NkBNOAzc8
3S43AAg8CwBy+MXMa8fkJalCfOvWAPS7g7Gv6GlvTSdkl9fnDBcTKZ1RECSqm9f7
WxFUANj5U+nGKsF19IwcVqHSo7bY3VrtCWCcvJDA/Gy3y2gX96pdQJtFHsadu57M
oogp5uZNkkK+yBzNQMPOJxZ041UNAHOGTL+3vmhjRY/U4u7UeB+VULKgYwTEAiZ2
NJoClnVwLgAHYIqTeQGs8LotJ0wiWZ38qLlUi3N63jquaCVh1CQp93v//4c47A4l
snKXslRtYpTKYLS32SZ+5OesG+DKa2j0mgSqyHFXHkdlWOqrb/s8M9i8PtFtO8Ar
Ser2TItVZIl2f3gAWVeY86tqVQfTUQhLv2PpyzUeGf9wPsJteOilrY7pRqDG24Pg
APrF1By3bfy9b75aj2D67xJthVlDZq0xGkuoDP1rIy7s8tUozZDWXj2RsiVKmOfU
GaEDElK6yV3uioTTws/Tl5lO7VBEUjBAIXtlPMAH7ccsgdcGMwcfuL6R5aGTpCHQ
o94XNmoEOU7L/hiU/XIXJmKU77EDZt8FDDRox4jBD/Or9yk8QianIe1k3p25xio6
iGgsx9k8G7ai3kidSBy+84zjfiy7rqOKDJTiaWvf28K+tqwCSXYmj8W1V0vjzlrR
wwOPO9urVrzu3eX+0CBWeWoG6ZUjbqhiqJawI9eQQbgz6yzVKLBnUO4vZQzbXFsM
UC4L2A6Z43eA+0fSYhZYeRfIdJE9l6isuMZLWYgOXAMtOj0vfMXIHWv6tgDfmir2
lZJ+Vq5XqBfFH9p4ak7zMvnOCR761FnMgzU2UxAX16VvQnFowVDF2FbxQlcA312s
ZNQgm6IgFt7VGXDpYjvebrftfkNC9taWEykAixp/8eNQzgEtyN+wrypZPMkxPdJm
REktXoICk8LzujiQRMau2Bx/OxnAVoLyTZAiey+dIvrN0VRtkzDa2JaNCKXOo8rd
9zVfMYkj6B54vnQyxGGbHagEEiZT2/THeCJ9xE3MnddngVGEnJz+aPmI5P86MMDv
togF7+xQ5F8yOLJiC8K+yg9x+8skdm4uch1l9VTgRFyZlR5AyEW/ceU/cSXY8H3W
eyD7UCc0jM7QOTwRwLj8m+JfcZnN5aZsb/B+zEL3vlK7A4sCqbKOHbC9NfqLEiBr
Tmhbhi9G/eVKbXwYKzaVrJysXi6fF+R/uAjXAChdfVXgKOHl2+9/b1AbYkIECVJx
997XuKgFZblKV+tDBBks6JtpEP3oIRtjaj6uFaQAEPDuNx+7MfVoeTwwufy5nHqm
CLtk4RRgcOBgaaIxGxoKNPYEZGZ2QrLofBL7OhJgDVZFrdR1WTAm+OkNdCe6Nc66
lDdF49d14MSb5t/zw2JLfK1/uu0kgiJvpuK0gPARcs4LyEnvef/U9GLF3ri8w21N
hU+UpbAtPoPAZfW7POj3D/e9/IQmNHxTcUT5YeQVq3ENDlVFfazQQEuxDyGRJqdh
FIMwnWtfGdMOgue+r9dYzGzMw8OaQ9t4xyOqRrxqKXRizO3g+tDUwZFgrwvO/vLc
weYEYpmw1sOclkyNOINKPByd6mH2idhWnwlChLpISbkbmRCOwrbdrPPDwYiRmGWa
HsMnPmQhTXDPDq/4O+03/WOegcznLgq9LGLz0RZ3kb0rbNYdXpAag8tjFJDLdQb6
ZR4DrjGvC1uBu0HzvqSvdWIw4DrXdMwWB1/xJI4Z1BNk/wtqfcCJKtWN51yItwph
L/2Kb0FySJISk99NmQiHgo2z5XfrUkYzi2loO1VutZfRzLikoi3dvXa3xW8A6Jwd
lLw3aR63DUOr4KyJW/rfmYtBshfSJhdmC9G/HZN+tCuM+/SajmjlQljBm7ebW2SW
dMyJFVfJGqV9vxDFn/rUg+lsQIMP8R/zxegdeiK/ysXyokLFsNTh+BVfXxR5Iff/
t8qJ5pPVvx2pm7F/N6L0b5JbP2Ixi7oi9sA+btC401WIOcCkC8HQSplpABLbr/7H
LQLXtx/KgsMxraNG2j4Q4yv6y5MXMtWJM2dWKvv556H4k9sFwfPDQZ0f3X0ro3TJ
1vjzv9bFI8uRUnymHa7BoPPUh991ocLJwdFGITCMXMVsBAlmFKeYT+TtZMLnRNxE
49gMjcMMLj3fEJMazHIUDzKUpEjP7I21rk63gO2Nc3KWqxFtxGQhcRCHWvZNUGcJ
myBU87ILSPL4pol1RuWkoCEKjy1dyP2wZMrUl/Ii+fweVz4qM8rXua2ujrh0sKOB
vDUXJRKipkciam+0hbc5rtc6p6Jk1EnAFGNTmcAzImA2ZabTp4/1yCA4IsfAjXa7
2PhKj1NPjNFNDDaFkd6gM5AMcI8e5NT1tQdiBZ4ZK9mkvxK3pElV1ne3jIz7lhQq
l9+YvBKlB5HuO3HwP+5L7F7SRcANU4zPzNXsknpgyJUQP8IJ3fZRqHuB2i5Ox8sx
eEs5oTWbNvMOH9wlmBBPeDTfPto+B/Ilvdv9Q1d9ouJv6MOBoita2qvbvGDkeHvD
T7AtIgEU6AxWGq60d0T2k5C7trLaxda6pwK0xZSEnUuxGtuKnBcKTyllX3wxSS11
7J9efcK236htWQnroCo5F1QrYPTMD3kPDkZ8lxfgIw2c5zUokmoedaPCl3Q5sULw
cr8JP0GeleKa/VJSUyR7c2RBeJnRW22JGP5hR5ruYMnlht9jm5f/vk4B0hwJKCJ8
3HkCm2Q8cD8xfs7O+IwJOgqvbT6EqWiHTA2YdeU7KHa3p0S97zeQuIUMuD/yw6z4
k/UtXdCVpae0EfKBmJbbN62sRkYTq2d1T8CXViRlRqqR3DK5KLWWTZG0kS1BdBfd
jKVJw2eCK4Inp5c+vldJox2qju8aqTtlY19qaK+AU3/tXlS/fOEr8xnndG2r4I5F
gTXm5qNSbi9kk07OcllpEALt2NHM1hN3vvDH22YY0mcAvneAoe7m+6rklFYjcN1O
gQUNLDU0wQHkXglIzACO0tcxJtxqXzIA91kb1Ot8J1pZsxlrIJ0Rb8GyxBgKJwZz
0+4D6IcH2ai2kPus0Ytbxw5h/x79z3qBEgRMg/MDWoc728qcPSet2tt09h6v0mzY
sRc41blIhYgWeYzNHGJJs0XbcyoCKPLrLMbMlsilW5gSeQBXraSBKt+v8zK9E9VM
b0s/PlAUmhi5Az1KvuyiyKwatfR9s54qo+muzmgVNuSgQ8e9pUzBDzZ0tHHiB06P
fWhNJ45DRYW8hod1B0ErhqJqcG7WWeJzRUIW8/Sq4iepbAdYsKtr/AucvGGsoSXD
BvDglGyHEIFaaKDHfHR6lj5ngcRJ/R6G/wqexuT10TnCjBWH/cfvyJ2INPug1guh
0e+It4sIVPbQPMMuvodX2P3Cy+o58I1cuq7KKfiQGYHPWLCtB3TDwBVEkPapH/U7
hO7QSiU+I9IOket2i9Pf1xuFlx9OyKrxAdHFW/yX9iu9qWvnKrpulSMrBlzEeVPj
SniqmJSOwVeYn9ahzfHzl8YnVq7VjbHMe2lLeHR6DDRvacm0xnWmUAPaNOdUPtWQ
jBGn4WqjEerFZDC/jybjIUChPIrwCTGh0gI2Zm2S+HtyxCVj2k9RQyNtwcpabUdX
cNNQmBj8E8UXsgwMTAojLWWUnQJeoNI5GEK/ZvkXcSQXTIJDr5JjSzlLZEOJnroc
+nwIM+yiUIUnqg82yaQeKzdyNZQ7PQU8dKNeOxu1+24cNAEKx9qvF88MhDUn0dee
pK+1Lr9LoFj7jz0EyEHnXg/oT40iSMaeYr1VHHJjFrCuTpDBfvqtuWQyeQR9JcWP
R6a2j0BoKU38+ntxLaKWrH/Ar+7ieCzIpD9AQoHiuvYq0TLTJ1aMXnSR89eyuskP
Ry2/7yFPIpwdA4ceBa0+n8kQN4rIrcPpZf488cxd/srpMj0gnARvWyoOdY8iYE2A
JxtIxSyn5w0WVM/WZfKVJoXtaWH244OJ+jGkUxT/p80NKq8JmzmTCBw2zqIpYfP8
RI5lOVivpi6/nIY/T2pZk6D5o/FAcK60xq5L1D3r0OITx86SQZcVSlcG+a8iqRhD
jL93usTGgnR4Wgr1sqgqPVcRH8CQ8nei9jQ1A+D1mLCqDyAsFXhMGE0o/W3lvmzf
e1TR9QUVR+VOeruZuSuFEfjDhHCzHRhVkz1P68/5wJt/87wQ/7x0lCntrju1EyTs
uAgQ8Of2Ra6Pn4eVTVHNU1rDPhVBtjahtPTG9day30x1NuH5IJdf1c8v/re6sus6
Vqy5xgD2quA8yYTcVC8YfFo0fUx5SrHgdIQZ6ZMh0S20Avl4/M1oZA5kpelDW/PP
iUN/U2k/Jhb+s+18ACQY5QC9uPq5gclezJ0rFak7RTgg69eBi9zYp/oAJQtNsHn6
cAv5A4kB2WTAdWIjYIZ/LfqG8C1YQ96RWRMtQQe/MzZ4rgX4zqUFSMs1zlnmUTno
K47wfJ6M0ws2KhcnVtxWmL9ICQFPBWgawNk4BDfqF/1uPR4T9Mjvm411RomiDQrU
WmjoFNUAiwev/0SxIWnm8S5cz1MKtDMgh5zpXyVDLwS61554egOhA4hvonE4Xq6g
zEmaKLRCPx8SMamXWcYqUr7UrLwUkRLh/LjIpm3rslPT/xGxduEmdIKRsnjdAO4F
RS0kjnp++cc7JurT/lSIehzqACR3wSPLzmkbe+6R927MkRMBJSs+mVDyx5b7+GFq
TuyLasfNoleDHFl+UyCaB0+4FQSVCA5Js1ij98lvzF6IIJqHaLFtuZ5gekfaOr3B
tbVsBfXh2G4KMhq2OXkgIpyN9SpXmqugIaGpDGDxC+53rjP1KqOs5Ovhpy69Kr1u
AYWkim74re8Gk308RthTMwUPmrc0rUUcwD4XGOnEEp+bSKPNtXggtF/rYxhMvu7B
+Bp45lVWhA9SHNChFMe4qY0eAFLr7VskpgUawBNrpk2yzpeJChwgGlUIwkxUDVBw
CeQOqywGNlKtB9G7/dUhu2vbQKjb7FAVV5lI5JOkHoOtlWz9IGKZlPeam7etMA1/
Ds/h/gplqQc+V+ceB/XtgIv3RBusY1Ml3EYwKELdyDGZKZOrWpVfMyrpTRnpc7Jf
4NtSzxNk+nLppZSxCCdhUGImc0yfUF61rFiJoXzUGE75iQHPE12r9FyBKliwls3N
/Snriggrfyc6LWxqqvjpzWasfd5cd1r9YFJ1VQEsa3PCT8umfgL3+NBmm3w7FrwI
S6JOXh3ZFDUIGMPyYirKKqtycubVdLVH57TEGhuO1Jp0JeGYqzL7uDFfZp//Zfu6
Tuo/mFcoDcG9mmBV+dsp59B/J/ZD1ztIBTAaon8Id4WWUm9083N/YKiZjlhVO+U3
4MoxaOMqRC+5Fro87/Zf9pLXyUTE3ImXkGUGM368hK8jJietZg119xz5aJB4HBTL
+Gvy7yXwg28c3ezfkO9VgRnW8kpCggHgIPFATh3PG9pLUVotaoBc5v85fQdfULCe
FGZ5VawrTd4HyA8Ll4BomKfCrGXzVu2DL1Mr1/UF0BEYdRqzvqxpSCjiKBTYNx5e
L1LYPfRZ/vYt0g5BWqkAxHC1yeit3FIX9T6kjgjsdvwTNwv+SpZtxrqgucEMMGWp
gjgXkqXQUPDcy6uzzvw+Nnf4EzKk7PpLMHIt/P2BPrmnj7EkrH18nLDFkLWSomL3
oEWblsrmbqVCjoay+peNJNGdPZVtO2crYdLmgLlHsGRjjTc+pzmV+fn1n2y3iiko
ZCcs+ks1glVRufg7iwo6a9geKyfsXpGFeosMhR/iYKLiHGDOuRnhBQmmHIA5Iz9T
e/NbZ3FtoDEtc+FMEeTMRAfJ9mxPrDb834pSMtpqXeWm7ep8U5/rSLoevz1NcQAK
f6wwing6p/9gtDOhkyMkhOi+qleEXTP+ew7CeuAZ3w/IOOq9knljmc3XmcIKKTeJ
R6Na7VosF3HVKAXsUufj1Br2Ltn/omo1OCVzISJ2WtHBfI0WVPbV6cUbQdMKKJ0Q
qOkmIcu2L5WzhxY83UAnKIeAkU3WWxKZqcyil276zm2Q6BB9MciBusce19k7/nu6
A/eW46jAqG5YjuXx4Efs40dmr+RGDMp3Dqj52DFIqMWEkYzfSZSWgfeZIU1PVJzg
p3GxHXturR+jqPdoWUR49A0e86yUkcTAILoAw0xazjHRcEFMR44YrBTsVXhPbNgT
5823A4gpsryzzP8NRhJBy7nTXmQepDy8Ncvhv1vQv3mcpAi4olesjGevpaUwj/HW
sgo859NzVGA0AXLjov2aQO+yhYbs38c75eT2D05/cs65QScViemHK/Dt9AIroyxs
MHfVwpWmXq3xfehrvMw3X7CR6keQotZj0Dk++zoAWuCBbZUhnB37FyLdF+96pYrg
oyAcw/pt7UdjcUmDqLk+lFR4X/DTVQdQSvGjFLLDWAD+l+Mrgk5q7lPlMvZ3S5+9
oZCHhsGPgS3tIoy7+OChRwOPlNNHnQJc5yUiACoo6Iz6YqWsmMjYflkLWysfP4eP
DehU9fU4uNpl7rYR0MTaj0IoYblwMjyjgZmU313Je+j3ATtAcX88IxaZL2PvN0SP
mHboroSSkAhKwsSEmrV3+kc8gwSj6Ozh6jiUb0q1f5K9OjUXngULS2/sIDaFaG5h
ipDjdEzyMWmNn5h8M3wuOAhIvLUzhzHRZGkb94+pOFGeXE9pS2zHp9njFIVlivvK
Teu2AIiJWuoIhnpZXqhB6CjIlSe5kDCBt0guIaePl4SU2t00FFIR8cxWVd71XgwQ
Cso3mUraUvowGbnKXm3G7teY8ekxORnaPjqEQLXYqfw25GYg+pWNVni+2LRqKL/W
Oq10nUlYg0HyfMAL01sNTkC9lBbbi0VYOCgZzj/XfYv6AgYKCBn2Iz7L9/90nzmO
I6fIIqvZbFcVCLvzh3ZhPq2IasBOZMEa0lsQ4Bv78RUz2nqPuQzZZgEVp+G029re
E5cP/TiYNujPQVvc0i53oi2qXCgGNnpw1FQe4fE6e2+VR2JK/gG46NQwBjshlzSY
2z8pGIqyDTxEz2V3wNEsRKwYWe/lco532fxUAZ140STAIvhuePH0d6eFwVXtO70N
j1VrDxpI3yzOEzzDLCVmeFg0sBnwoRhrYbanka8Fk0kzAndRrJqPyklx8QLA/NND
NPcOAYErfLyqLyZDKpjPItA2E5euczYyj6gkg2lB10JTSFPuhS/SP04k71IcQNnM
cXWksDxWrgdu+J/u23lYB6A+3QsoLEt8ZwpnlfIPGS07WUBHx6hpxTImMfh9nAL/
kC9gsC4BIeh7Rr7dj/dSkZFMTBwK1pMPj/xeu3Kf9c1mCFNlznoFV396I35Cg3ZJ
unO8N286CVyigBUs34jBoP8jwscLo6Ma0IbPhACbqj8NSQwDPrL5pNBvkAZUndpu
1wjrVaAsJqKTDmSQyZigtR46lAy7F0c4stq++DYvWvDOuykkEAKUJsYVARNA/mr7
fOd/yUUPQtWA5dvh6/ziUzZZTykJd1/fCrB7G8nrPGQfDYEnc9nYZEHXhObwDO4n
fp5JFr2oFN50SYbBglKeOXAUBT72u6SMCwFyHEJHR2ih8pymx7LbkL+qMLPXD3O7
z+ZXR1jgUSv9vATjfPKX/gEDavvXtb+uhIc6gqIBzSV77iUvk1I0ZXDAu01dBwj4
6pOAM1HBypiVTtDZDads9Y6puofsjq7oU49TtGquodLwDjq2XZpkr9UItor0+Pj1
QcUeyk8tfW5T309IgdEGSs8DLZ2bhPdCNd92E4zoJyZBE6IjeMYIY5/C9rIp9DyG
ld4ML322IR+uIPyDswsjlOAMANknhXo1Fj3nd4+za4s5nVWsLCxwmH628IhElMLA
QA5anHN9qEiKWi7OIk7ng41YvJfuze9Q3iBhfulAjkuRO9mAyMn0VWYQk32a0nl8
a3Xu9zBVTOjxQ3UqggX+OFggyr0a2uiV/s86DYBoOJOgP7ptBHeTxmOntj98uXwz
cx62NdEZAXxjgne1KKlLZ3YeUJ1PxZtEr09RtmwniFF5DWtV+rFRX1oePJVDJtZW
v4qBNwLmw6/8PzAExVPRp2Mb7p4B3YolwkWKEcND9gfY7o4t0YCzkC4JfmJhsAHx
JW+LglsEXg/l21lPaiwNSjBAzrqbydwRprpfRpjXDezbiXa6VReOPCtJD9pCgvvN
ZtSnrs730/auHFz61y59sncQbibu5eDOWdeCp5M63HTViBwWMK2+Xig/iBfGTw5s
dkbF0uDGvwzN6A5Brx2dUGAnbGAwDicjtrkDS1kem2HdvfGsYtKf91nIDabV4bER
+pnfhU6z7E4jeaHVAzCIW47L2I8ScefOEt3jjsEOjDl2/FwhWU+ER+Aphid/QfFG
ILVlBn8Suh4oLtHiIgLONdJV2JzjODYFqW8SYMNyhfyBcZffwcvUnOeBqkZeR17L
03VnjUKDLdRxBjClbp3A8ohbUEp1VjKkbOkWTwxsJVx7P90ULCqslMMzQawFz8c/
yCv9C4mmievggpkmxebITHaPErgiCWMVuKQAZ7fv0SSvtbmGkkm/PqsYZYvRMdYJ
MUt/pWa0dSFb/NI3O5GsmdwzXITmcndYcIqqYIqmO8u76eO8B7t94vF5cAZRkavJ
CzCiiYQrEPMeIrMSXhFxtkPZbv3S3XgqeXm9BbecnsqeqFtaRxiTo4LxvlKDbcZL
CALxNjkZzV0fXkx4UgZbdxgIfJdO3w6/ZrHnxuvFutesF2Nc3imUnKVVLtPryw1q
IP/2Xg9ezVkIVkHyeKR10P7rLaHOz+SN0kCp3nEjInncCCMHD1/I+D8MLjGkM+QJ
sQuLgBz/JGd7UJJ2Om0jJ92HBxP7Ra63lbZ849I+CUFXOzu/jeV23Fan3/0Fdi75
hVm3rSDJZvYQzCvAq+N6T0vyMDHUg50TUXKzVW3rtviu1VlCVbXLIdYkZH9gqH/t
GNqqpoUxvtcUlySL+p97xPFkxBqs3vVUQDK+0KDeFVNEvVqCN0aeXE1KfHLGrSHy
vDQHtb3Ttq9k2u4xO7o/uhMcKTXo5mLM+JKH5+gSKDJT04HA5SnJcjZW30xFqISU
y6DJV0HUJegWO2Pz9JtYKY2H2xeBBVWElMZZgxUVawerWvIBZ7XGvIGPQoSxgeKI
xQgeFFjXSn8l/fIyHhC8XlRRh8kBSdt8XuHjCMJQGnm1iNQWC9doGR97bQycAeIv
gGm09qvax3YUGOVBb0FAOY00J7BciB4s1uEuofqX4dloxIumbFRzjRPHvCd70LTT
Gql16Bxd87gglXPVgNLpifOrsiXjo+LX5cGWSu0FNjF2T1Ti8bjWn8mWAVPlYEDX
ExdobZwvTuJfGEIGqzMOoWMDOSi1RX0N79Q1ELE8bgAsBsxeIpeU/2jIP525+3vB
6more9eiIFHzvJb1mulEy9tTZxw1hBxQvmNPuzE2J+F7EDOtdSNXI+IYv6foECMh
q0lfQFWC5tMeSxozxSx9gvMI02fimdZ0i6Cn4J2mMOLNynRol0Jms5iSxzn+lqgf
P5LzhdSNbEbrJQT9bJ1/UcbVaKk4w871ua+Ygx4ZLid1LV+qJXUTgKp2WZQZmgnF
mlVkfMqr7DcxTPcbeQcRZGi5i/UIJxhh+2D9F0E1cNWxlM2ZiasxZWgGa7qSXpF6
CnDwRRJQHIgE1fGKGOW3JUmfLJ9shMQ9FhvRCz/mvBY6kgHqG800OxnQ4Vk4oZxq
0l/sHZiUhv5WmV0GUrEm9PN6OmFPifhp/v35U14CuKcYskSVnlikW4Q5ddz/AexO
RpDBhAwJnn8iXbl7RQI9ii/7VZaTlVf1AiP+SlEG53WXp8IP35VvMaDIxpavcv9Y
BBT6SbWYqeDNVRFUKWoQh9SEHWWqlYwg8ga95F66iwNyJhlG7iCs5gFyvp2z1L3t
WCspZAr0E59tGPtshWQC5UNz918vdz2/2TqZeBlL2CUSBedEdF1nSAaXMidg8kAs
nn572Jn0kd5pX15QjKY0vk5xSGTQj46pi9WHkGq7+eGFiG7oUK/2DryKlmfS+zaG
YbspVpNZgRyblOBXTHG3mzckv9bO/PO+65FxlYImQlZrqGGtyyX2f69nVsXr3U+3
5NBRrHOyOOEyFcHzfjUnlYWkjvXETqVPWNBRLDDh24xyi0rl8Vq0dFUE1iE3ZgDM
n+k4al55GCK6/mPK0LIxCwlSTsEZOlT5i25Vaa3B0B1HWVJ6+t35tuXVeYj6o92S
4rQRM5E7Q8Kq9NfLY0GV/oetQhA5BSss7MDbhUUpSi1vs4WqjKM8fBu5ZaRASTEz
k5AWVW+BwKaYq18CmAm3hCsuwk33EgIxnNT6YvUnxs7mCfn/tPEMHnC3b91UdwTT
TM5G+42E/6FZt4qmJofNGAdQcHoJATQ92Xn6WRzSOanIJ/UnkmaKSJ8tE1+VHbdS
A8VUWKxKLLwabS+mu4bijC8GkUpZiUxwhzd1KPHxu+jgNFha0AJIiMZKz7zN5Fgh
pHLAPjIQpJ82XvQUA3eG8wygvIKCzBT0iHMSVQEiJNtRkLB9NUnPmktUavmfKCS4
vv4I/nnCPU7Mvr2RKSIYGD0U0tXpjzgBfs3Dbm+jao8LOVPg/UkAp0nkrx+sRNzL
DRfraFKYQNSOQ/Fp3KHxUOIUrdeJfCfdjgxmfSODEIyRhZoMeqfAgfMD2absi+P1
yQzjDQ7HvKIXQtGT9E7V4FlPLaShy3NMLfBnUib1ud8lyZBvwi3e5Q4N+2BS3coc
Lf4KSAI+KgY7cT2llqwmQQoZ2VRvBCw9trQpjIuqAnKbEYAHhuCd+y9o55gVnl5Y
WMxYAoX6NPBIGSeisKKn6HF/JdAy5SUA1Wqu1GpMkbNE8VGgfDo9pZ54EG6mM0dF
pOEZua/+f/lxnegK/LNm7PAFbXwutFs+Ip8HLBDwNR1+pz0YkrR9SzEsihwb26E/
w/N3rRCu+jePkHmXxpsg5IIJ+3xTPO6gd6U8EUahBz6uoCY5EY7wyciemEnKqTZR
ud7G5LbZXMFNEuHLAAzdu7uZnTFb5yQai1Viy+ojpHG9u7bpUVFZ+KGGPNpeKp30
PbGhP2OlZfpZUcf+1omB+370HBSy+H3+s7QqElSDb+rB3PMV35oDddSNd6DrVpsC
H1BUAOp9HS0LVIKf0WHjDnSFqWT62uujCQjv6TEV12D+K//nOATwsaFx4yhOJ5BI
SdAoy9PfMuvjxoy7k/bNKKYRT7GlxG0AI/gG6d4Uyjb2+OuN7oi0G5xi1G4jy2BY
Xg7zb+fz9leqC6EUch9StAR/xd0LISJlJ1qiEZdUlkO4len+HXSb8aFbpJwGfMri
JHmNv2iegIgKyGl54yBZBeFUm+RZeBFRvAP8IeComRuVN03DIlRAnKyFKV7WXfy/
+kcMohg/1aiPPOFlcMZqKTxo4Yr+oTWThIZxwRF+6oeYKkT8lMDH1gJwz7fubzn+
7E868aqarxvlz275niQc9JEeNIoAQ328MPwEmjqpgnfkStHpxiV7TFxSZDUs4RMg
LGbHG2IvH6m3SMv75lrcrSCWRIhP1UWs/131VrK0qtSkDniVSDOfH/aEGp8lXVwN
TScn8gRDsH0hXhI+WIJ+Jo4hGNSk9TNn8jnNvzxewDYB+pHPHib/34w4bTd3kkKF
0E8+RM9crHIWhvTU3F1vApWOZbiVfaS3SlEXpDw6lUyY6WpuWD9wytinF5OYh1LZ
kYGhwH9f6LN8P+XUEbHyXwCeMDMQBIjGl7JBSXtxnJnFNY7A4CeEgi+WP6YmoO53
K4Ew0OtbrNw4O886xJ1y7Q+G0bIsZL3TgCSjvTHU3eSWzbIW9/gdeuaAw6KhGDcM
2n83rXK5fscY2GSJdmN0SbI9Gb7+nz3QuajvQfk1OK9WYglwQ94He+rvh9sodLLQ
zlN13Az6KL+6gMl72sn2uuJ/sgbUnaxWtxYXGYBPxv/Sdmrp7iT1F96SrMJ1m1Zk
YpBPfY5t2xgHMOZtM0stBFk3M1NhFC5jGUqNEvjEeLLz8DYx0fe5Dxn1rSprRr7/
QKtJm4dvlAS4581KMNc0BusqGSPIIyc7qHzrWJQst+Eh8e9RuKw4tbOFIbp7a0vt
U4I3ys52D091KHniWzhmQGnGdbIhxF0m5hUOjj8eriYaPkWkpZ6ua98ibDl2YDda
UMO71npEZKoFwQWolQF+SNmVd01l54WpVeIPrhQVeF/ISiNkuAWCXMRPWER8Rajy
QrGM5ScuHvL7ln6T6ccSOp3TiWMphJvI751/TJl0WEL48v71P+MPAu25n9ifeLCA
fWMzsS7Xiybj92pN7X4xbXt70sbPdwgabqAWyfokSKwTeXwyGT630tmeC0xlHwSw
EO8CBkBotPQ5d6+Ehn6A/39LZJTLUl734prdRsOkQkDsHFLkc0jBruN2fdgRx07j
OIskrADtsVskAEmD9DZaw6MW0SWiVYaKUEglHuYPJDfn9vcU6brmwZLkVfdgMxTn
kbctRfllaux624Zd9kq9tFc6+lhqZDqIbOf94yugZ2+H4DLXXxX0HNa0Mpjq8TyE
aahtSfzzjvt4xW+SRvxuCoPF2kE8SxBOCafawJ0zXvPb+V6Tpry24IRQkb2KXLaN
frnIjwdXZZ4/zp4oc+W9OWsBfGZB0svfKngQsz+f8EKwOLZsAgmQzQV00d8CjMHG
tz7q0esc+8UWCbhQqPHUiNoB8xLt/tj2RJv6IrF0dXGbMPMv2fug9TxbQjQfuK9L
uzTg88aK6ub5aNWLTxgqucATK2iJzmI5LitixFV5VCTqmLfZgrA4yHWOqh45J/Kq
9LfIGgTiTFBVYy8YLKTwBbXS7CIz8TBdwO7rm1mg4nYuW+nmDlP0m0Rp8JyLxaPc
HotPy4i04muqTrpOEzipAW9wj5F7KcYqUKMTnR3c7NnEUilWzbM8hHqYu+ckBWWd
pzYhODMx+BSBl9ZEIwH1Mw9cGG+ds0wEzaS8PIfu1xFq0xrVV4PmFEyP1KRrNH9U
uyIwEYx/SMbKQGet3mxblR0Ww+6XXdINpI0x+mMRjvZtt7Rpj5gjHtMTlxbuCY12
x4EftUeYn2JR02RpqN18aHuZWaiOZfG50YHwTA/cdhe+ZsPyff1tDwhwMJ3g6rOc
H08PJ3YFIaUm2+nIJq7XQa0DzyrnewVc3X+o1S7vnLiin4NSIqPlOOO6GrVKsfzM
2XqogfxPWIGzv3wa0QHmvGbJMfZrXEGKQH7SaDLER0Znr8S489SNQZQS5WRZbzWv
iQ8ncTndORK5CPrkUcfdvK0XtbAy9LqV7DeKdnD+EeFmtYP1W0lU9WHFckOb2F+D
PC8DPRvsFOwZZ3YHSi1VXxsdEd31Q2cUm5Y6/97GYsUAwUg1lMREJ28cmeHwYCjq
IehDY5dznIDhDS5S5jF8syZbl/dM/DeOrLHfNOz0YclXIXMJCd5O8/LQDR3MUi+G
GVn7oKM1h+8HAPes4XnUldnbg+wmhhIH0eVEiXBqRyieWEW5xNSKiePJJXRphSmm
hh1UwOdkWMZF1vTgAyydM7AxW2MtbLdACAnGB55bRjoSmVN9Q4+bZJ+wg/uC/2da
ezilHPnLbn+rF70G+lYf/4VClzGOxEnmbnBwn7WF02CTEpz/ZZeA4EJlxiyzL1UQ
zCffBhNdLGU/AzyqYL2KTW2SfF32XhEaR+OD3ptUPqvc1NXDc7gLMQsTyYKpIG1x
t0o5upNNXUButsd9u9w49H/UFBH8DOTrKEpY7Wu7OUUABCOXdIZLo6CnaXOffH31
6AtjU4qfehcVk8De7IJMaKlPnINrqnYj69BOCuEHqW5oFbkymOcAx3LXn+w/zNCh
HcZLlddK6xOTVl9CAqGixZgNUoiQsSFhv+GUnLPCIfJeeHoqmIYOh3/j+VadCSff
5L78H8kzxICjkNPolbuewfbCcnVRvCINRvzWXFwpdN6jSMUs2WFSTIF8uEEUQfw+
6T51kGjWgXjx06AwrvY/lQYGooZliml8pHPZqbmczsxMjgzsYtHJnT0C9Nbk5iWK
EMi62Cf/MyqBTPRcE5X5XCsN4pE8tEpvmLq5MAAwYM6HemO3DXKkYMA2r1Nmg7zI
DHUdD74XNcJo4E5hwsci9567WYvsmppndTz2aDFOxsf1tu6anYVGwSsyW1WWCS2m
AVoA+dTX72cQgkeULXRQIeAO0Wr3D6kmcAX0CGn2r96PzEQ63K6QqdPJuNGhBPr9
HDVDnC5FZbFcrGGxiyvm5Os4DTk1uR9jFHVQ/ganTELG0jE9Kxs6A+iLwrifBBq6
KTMPGG46HkbPAoUEOJOUEVQxHDqHRB5W/Gpi3k1u5/EcsEsEaR/0o25IQ49Mvs9I
5J+V23LeRx9F3XibcKtbpv4WfRYuN6XXQ/CTBZyvCUweM7pAsYZh4V1+hULOzWCv
XUEF1okzcrAA5Fj3w9sqZQ1B+Jy47j8VgZTukRTlvYJnBSIswZH6/R0oysxvz/Ob
qIIl6fPFXIhO4HCFjQC/bqstlclnrpkuKYG3epODzvd4Tuj/NJUC31C4UfXnaTrX
0oEUzY4kTMh4+EK3SurpK4R7ohBxudPb+gnKLnfkCUvIM1S23WkQjnm6T7QeZCbu
8o34JJDRAVEPmXwQ2SnyfqPozJBGTrEPQhaLQbTGzaPu12cAEtvMBp40XkakQt9t
H4QqIWfB/9g3nhb3YGvnVBK5fFRz7FYJLDTmk0f7V/ZG5jF49Xm+Mp3/ra64DB31
s5bl10kSvBAZmQFNCqRMNU+1x/7bj04zlEYClob+0/9uzurRpiZ6Ysgk8xlvPxfH
/quJ+hgBCNTDiTBwuIUnSOxgaz+7Qx90cirWQfplBX0XX3l0YlnGI+RNgOdvTjHc
5eGpDkvxlY0Nl6TTvg8z4RzUQ4XRHjfBQ1JMqtSS6+EIK71re31t/1jRXXOBQz57
J8rFHDjQtkkOxhvQe682uMy0iqKwbjTYNfxc4NhdssDjcRv0hVEnM6OHUcwEz82s
ajJzQNYDnBiKKrckAsYfCH87Agp3CBjbok9EvzX5ehHplUfUt1Sv037NwZb/coEN
Qw/jnF16Cle+fLClKbRFLKUOMTpAzDUbTnnbRvoWg3/tFw+rK3UX2TFghm31oTfX
5rh6o64t7z+k321PV/9y4MN15JeLtK+ZEW8bcNM1E/Go0dmu0TjfxBUCU3VcPYVc
1oNF+lPJ+M+neZdJ+bEAjDIOX/fGNQbDVpOzIscv5cArXc0G751iSy7Ow17QuPJ5
QyVH7TzFZNFOI87/qWlziHBZZt8bbLoWzih8QsYuejPb3bTrKKXgVoEaFKBBF4oI
i/5BWMll8hszj8tPFasPdeOGvHfjGqegjBKDz/DW46WXkAQqP1kflPfTrg7SO3hX
zPfLR6mLNRCGJcUz2JSMbYvXPOfKgA2cReCZc9kgjMB13pMcr5Dlo22vTJbJV0U7
c65ws3QcC4oajaZtZ9feeZrQhsX8ID+PDaLfr3Tq6Xq039iiaclNhh+grytvk8r0
LYamX6tkIRBCdJBwi4RubXVQzUEi4W68ipKxa4aFnf6doIH40LPtYJ1C5K7GojHy
CvIFKitbqbrUYB3dehqCZPXDmZD1ihCRf62jOGtRMEgsGnqV0YrVPIp+CEXwY0q+
l6u+xac6ymYsfj71s27XS8qZtHObPj6GTO+Rb91xHr5btjfQCkAoTXRgCZ1xmNLw
pOSQGI6r1ACpWcVHbRtv+BrYqAMJIvv7yHuguv8Apy63yzNCF++ij8JvYQxlD1w1
xqDz/pHnym6pCw40A6MLLezTxth0iRO7WYvlfDKNY8v7klcGjqSbKw04LJBPId96
Do44I6tmqj3ohg5VgwVViEGeY4D6iHTU0Oq4WNmGQalu7oSH1FU73cf6UYFzeIJ3
HpGM6Af8mbvkTjsw/85tFHFX2FiKSLdJLSN74cSZfDbFm7Qzsw5jQUDIHlqY+N22
+eZ4sBCdvZlb4pGD9q/rO7hC69oKuQsi1xudawxwonTEIX3ywhkh0x+tPl70mycn
5VyoQd4UhJhvU9ceKQcH/slRubCQbzn8hjsgkdpNBmhdo2oITxXZjCXRN+v84mny
UDKNq+HFwJiZwXoRon+e58hC2hP+KLZAsGlUk6TS3RxMJ1LVG0IGiH5p8v7qEd7E
pky45rEn0OXgGyBL9nHqWqnkaZosH0j4NkmgiHEvrCGP8m5jRT110uoJEZQDOk0S
b/PqpgIy5CqAXo66RPbnJ09fxmjM/SfsrYtKfTQO95ZKnx1MrNQz2IzJg1EF9xzr
PnLf0MP6rHibmr0hISFlePcwEKSb68EsxuzjOjSESgZ/pAYEqb4YW1ov+6MnrnTo
LC+FwpGTiMV++eyqt9KhXQND68jy+EIKYMRgNOUh72hFrzaJg8yJx99uMkFOG6tQ
b8tazrRxjrGTdLNOoC+NAloyx9vp/ort5UnZqaWj0ODbWPrJ6B5NscaBgBeYHji5
2/0uAbxL7IutnODZdwBfgP+VTV+wE078m7RINIiUcIPOnKD+nrcTSk7LmA8RMWjz
GYA1DMdTU60/aGWl82JP0E7KLVTNHTlDV13GMUg0w/YQ5Cr8VxHMbORSzJBdsh7z
gs4J4fSLlJPPQmBbmTFlsWdCMqJHVCpe09+VJUFlKrb1OYvRT/xIumK0Q5IHEAlq
GVhSkYuSjzC9TirndBLNapt7qCTFW+Wwz4g4EXLx2/H+UHHSivBzGX319usD2mu+
pDZ0r/wZ89E1eL5daXrYrnhb9GP9mACnGdwmj3dgH1TCxA5J9Ow3SMRTnIVu6b/w
ZkgjaEsXbHbyw7uJO4XCJZDa3H840kFACATyo/ZJUEYLpa9xc6IDVwHYGP099Nvq
UbeQCQWMsc2d2Hp4iCT+RyXtsOnE0FXLOdMLWKnNHxVOUDj1xYZ5KREck2kghCsi
qcZp4pYmGPFRttxilgjOIuDJvL2pzFPRXzkpD+5PRzOas4dE/1T4chwbpxjHxZ2d
kO4n2tq5WhjUR/wS3knyUfdC6o3SBq7bBZ7YmpWDByBoRmPxZse0TCKXOiZxwdCk
WRmKMh9sOOoOZ9GeW0v3OPkSUX7wP6100zZBmhJu25OM6eXjPSpClygcvKEgtfDZ
O7OH5uDj3dxw6x3sq6l5srxAkXGOJD9+GLorZPcgz4W+S1MBJuhlojiwQvWYoRPS
+JXEM2K9KX45zkWoWQXFgOakG9JlP94YaNNdpvvlOX9J+LrAAiCmPd1k8PlTl4i0
7bbmac/srRwV5/YkvGwBDu/0sXrgP7wZiGCQ/A3jH002/egRBWZn3mgnYHQo/nEA
+IdhlFJ28Ek3WANO3jiiO0bgRtaxIFo9ttQm8OHu7gB7hxcPeqePAk4kYaq+bwZ7
IvwexJ1oSHRrTOw6sPO7YdvUqVGSFbjBYTjkhpQ2ktlSDdZ7IONr+DMv3zTO06WI
rErKxCTGLkFxjxaC6GCr4/R7vXimNrD6OiGgWJLGgYtHBQEk86UqhoRowYW7pgmZ
XL8Vr+CFp8DFYdV+qN46q5AHzROBPbMEcCdmmaL6qgRxc+Db1lzBGlTWXtBWG7d3
i4lOIBOduF84cHmfTRcZDKt1uGJh2w3gk4FVNw32RbRgj+bek2FR4qwQiKIhuMsA
cYspoB48EY/OVs0iEftzYyrflpGWgotGGr/OHQMurtWTnFKCn+cRujVLLHMjCsMI
f/C4eJLj0rDcwgXq0iSxWOkuJOXOxDbv7FIqEw7Ja7swrsaitxtO8TKFD6K9SfVh
3KjYkA/+OUpygiARLCyD3zG+Briy8K/HabY0OxKKdU7BLahrre34/f9dDsjLlbD1
daiHqrF141J4GoskJrqORAkImS4K8dGQUea58k2j9QHJYDKD2JiLmSQSOaAZg4Zf
aIu1d+w9PxpENgk+NbKl1Jtmofe5gENbrzrSLzID1zEFPevggA7Ja3/a/6dei4kc
7PPLs1GDQKLhSuwn3HaMkEuZtay7obViO7jaMT2jkpJRis4IV3aKsJhaBB7rE/Hw
RLpLGSdceNV1Btj7fMhg5FLhapGjCZcX0lUW33Dxlj22q9boLI9Kkqj0SXm9ZN6x
uoSgbBzardcOABNGK3OMNB+8KrPhAfatMDRRST7I9SUq6gKCOKKgJxEdXm/sdqE7
WMuRlbbvZY/3z/zTtojySL6Rm+SYPW6A+by/8CNA5R7OA0e6/mcZ6p7sk+MWqnWC
t/ec3x322J9x2DXEqf1QhmsaL1TpM/lYXBy6ogJH5xUNHqXZrWcD1wZZVNKbkQoC
GqXU5iFYROoDQVusuR/4TwhqJa+bCna49cPLM0wN8eXHYK/Nc4OvmO8fP/nvOY7z
J/rgKIpex7pLTX80vgRgXwVSi+EgNYI2qj3s6kicF4YvD0c9VgJujbuQN6KP1gxF
5rZm2eYcHjOp/LuDmngOV02Eex5CbBvjSC8W6jIaDzjsGUWqnUvUHqi2EG8U+B2s
GtgobvjvMWVHTZrwDFU/3PsRUoPiSlnkEHVIFT/SsoSPQUmptN9YWp0YzZLdMSfo
JlxMPysVW4Ci3yyrksu9kI6Iu0oXgHMN21hscASisCP7l8HDNq+/FG2RGV46WTJz
krtuwho+HANK9uuWZblKAKNTB67hBDVVCeOsOU89JDaeOyE05OXGfA3f20P0HPRg
CUUfkB+xybwNS8mC3HNb95JWjOijfpP6AsT5lu37GYs77p3FNjgKEDZwCfpCIGB4
Qlkg47GhMcGQVPtiZ7TXaPLWvFLm1TLVeuSnY8dK2nvbF0uzrOs9wwjSx43wq5Ea
FxcW91MY9uE3Q5bNEAT3rh7FBwSG/x/A51RBCGKSxAaDtnwHkFC8zo7q99EkB5fe
bTOybiH1YgKPo1HraEyORTxjpsvntYuNxBmXna9kCZxsOyGQA05RG3hMWzu5XRh6
EMzfn7esIbw4vACzRbyHlasa3iONu49MMmtAlzp1iEf1RCPqkP1n4GaDngjnBxJ0
BMvh83Dyc8OktfAlMycxGWJETEe2WrfGoNmUMVgppIafj7aMgWGcsmfzjoryWRwn
Z/edpGvqO4KoA27SM1W4iKoQHyOuIFl8dR3T6vzkOQArgEaZ7DRZFEQH2LpXPEue
R9llMrk2BKL+UTHIWmfkI17CMXUDU5h5oS+2oIIPUGHb0L8WMOC+fRX3jAZuzbnd
rLLLI2al90UQTEbvd2kVypeDDXTo7bj41jkqJyDu1SkobTeQnurxxyTgKiXQs8Ak
6zDS141YfLf32RcRoISKZFbE6OZ+pIiCrHp0e8ebVycuGKmmhftGDW2IKq1JIaxQ
+xo2Uy6drqGcC75mymk3eK0DcH3EOPnM5S1DjR+1IlFhkxVSKvrcp3KGBbQ485hp
HX3NyC5gMxZvP8OGi1KqFWQ3Z5D7WgnWo0t90Pvm7MRPK7H2J8KvQKGIsXAY6xDo
vggW3ifpEVEIPlCsiWMCadeNUo0+SwTlcmqs88KjWf0oZl2mXUMY0uVFdqBjSKAr
dfRBQkRuKwwcjaZgM8QiVv0tSH1nYYRqpW+cw7Q2dovGq9KlGUflQz5AiAA5JyoK
K+WDtft7KRoYhyRpEsiMM5qWVXF2gmPSj2LBzcLK6RphWNWOx3bXaAyhMm0c+BVt
lVbOGIkPQ/tUGX36KBvwC7I9EFQCXjAhru2BPujD9gJDm5IHQzLx1r4wwaRaHyLj
53D4t8dDVzn+s12cXS8nVMX6FiYBGCO/zQXbO2UXhFblLOXQ9fMZMufihWmgGWCl
WzU3jWTtl9n6txivWPMiDVMRbWCDEaE6WzQSeysdSxGzVpShaBz+MQG4au/t5BvZ
6gSRg4+Vzou5XvD0Gtf83KjFYWPzf0lgsHeimYo2dMVZSBVo7SJbfbQxgGFVMDhn
/hEfSz82w1BvjcF7vlXEuUe5oZKAD6g5/9+gtkRW6O1yNSQfIPG8LU4AGJ5i8EYh
3dp59znZSbXbo/vl/g5Azg33MdCBYM9iP++sJwUWaoNdSzGBvUxV4L8kriBZLS3S
BIXZalMUyNPVbbBcSys9bKv96IPrg9GaMArtAdw1t6yZfEGzbZsjCz/6VVofIQWw
QFqHFFdZW9Vi0OKId2Vylzj996oVR+WpB1X5DfxWNO+S+VtfHK0AI3Pj/etAUPYV
X4T3lc0MjutInUxfu/0AoS4G+pNL6Iwd+O1jLN7RDVdYryHGCNOXGjye0yCEHeCr
5OTle4FckLP1mFYsg3NehBU2pgATivrquUJw4EMnNavGoplb/cxy/rrnJGOfCkBe
VhUR1JzS/7wxuqJ4FKBHdrF8dsGnSzDaUYYVk1cuiJ58D4mxmqY5fPGLs6byzCit
1K89IPtmbeZgOLIJlqfcLoRFHj9QciEN1fQlOebzeupsED8zX7bBgKNzBfQ3juWZ
XkDvkEf0xUZm9DxSvc0iWrMS2l8A+Mpnnz9rv1jgfDEBCiZRgsvKKR9InEo2gB6F
LXl4pC37pAiLpzZhqL5GmLxb9rKwE6lYOYNRywbOCpaqAoX6I79FVn6xRcGw96qx
j26dHSwONq0vPKl+1EEcG+Zfrz8kAfdQsL18WElx46yQCMl5xh1W2s/lQ0eA+MG6
4ac9Korr5PKEIn4qlEhXfBmReIDAuzWW5S14s7f9ygGqHQn2yVj+SaNFADpHR1VV
wuCnuz1D3nEvwzgWMNX+ZaKRX5iN1BKYExuzqJLPP1lCNu65Wupcq3bKme5SGqqU
bdK/LGkkf9DtTO/bDU0LwrStzORafhdLKh0VfIfXR9XEYVVPCUfyThrFKMZN3Kkk
gjuNHTK1JM1SkFVPeeue59l1C/BIL2GNVk7GJDRQAx9MJz4/cvC1QTN0f4ulnrkP
sx5e3/LQtKp+BzioCl11VViYrJh/Xey3GcGZOLo7y1Fp9lSAfMyDC/QUNi70OiqV
qkl6fUOEX0TLSI4KGPAU05bbgFpSWCTX4WQ7+RO0Ho5v1nZ+HaxqMK8lMd6XpysY
tztGiEDirLBDW1VjcLpKvcOZ1neQm0V6Htn5etCNYpAv4ohyvVwoDvBjlD60Qbbs
A0RFzGKKD/E3Ekqv4uG7wE+UvYodZPwgB+T3snR5YTtKDvbWgyvBES6tQvwjuHTs
B8LW/BSmosaRtG+c79f0Bdra+ysxqP2uqVhF0Db+nCc3J/q7oPzB6d0+61mYkkov
m+ogNsJajrLmiCduwaOZ6nJYsZdboJ/nVABn1A2FXajkj4pJwjLfsBoUcClQojpa
5krGu7v+0pzW0aCUCor3UJ3VXrNL5uwDxDGObHka6VvcIFzTOpwI1yf1ev9yYTTp
QXqFNo0FVR7a4CQsvK4K58tRP957QD+qedEOk4laYsx4AC/OPSM5Sld7dsY9sTCz
yad7i6hKBeOhYCUwv4HeIxhyD+4zCiqK22+X0opdFTGi6oHbqDQ0jj/s7+ZDfzJh
7wfZHHL4O7DZz8TYQ8x9gtY40FUJMgntjHbydbnXbk2+kXKu/tULORHjTvgpLcvV
W8loiGS2GVYqFkzpnYDoaIarW08z6XjzJjCQg7SrptaiDqtRzWO3hEvztiUAGzZQ
Sywn4Q/t9s3/MoispIuVUPZ/elZP10v/fQYQGGBogqXT9VWGwy17SHUfQ/SjvVU0
wJCQXGlqTo1odIl8UQMY/Dfxxpc42Kxnu4mlR77i+35wv8eE3CYRpAD88ieKP9xG
k/ZpqMm4rCTKVj7vc0Di5cqEndzwluPAOB41Oz7vk4rZip4lM2q7s6Mo+p0OYqM4
elbG6Zm2HbY0TSN5EWmFgknVM3uPdqbDoRvQosLGOrqxaeFcKkOLj9zv/2vPVf4w
ptq72i/a5nHM5QStfY2ulejitn3X6NYXi3OuxDLBnEJsorwpKwlOZ0u4voemlJNa
4H/YvQi2lNKMBK12mxQpDACRm0tc/aCQSD/f/OccXaS8Z9VHKByjz1/4mix+8C4C
53Llq8kvzfgmdPdeBQtV7bTtjpjU7lhJFUafHmdThF7Xyc24TCWtviKZnrZ/apve
l9n1ZEVCK4oawZyRl2jcytPd7/X5gD2xtHgTyCOy7wGUr5oWc3RWhSnti3KunMfz
Duhx0DWA8AK1cnFbGHphQOQoXSrAURqR+32HbLb4umAYh4lxL7Zgjv7XnJy+sdr9
13D4KqQsKFz9CeN1PnoyJOb4MU2cJDREdu5yMaM2QABpgDZM2sL3V70dpqgyg5j5
IlzKK3+Ikl+Bkyf1bYuPwDn30A04paH43gzioMz9zJpmoXN5HysOn1zTugX3aGCd
Da38D0Ys+C1pbeguAGtuBup368UX1DDCaPDFzb5yxlFldhbGvvYbXT7iGbIeH1Ee
sD7GtOEZeEUHPYwudczDykQxYbslhzKtiMtS0WmZoB+QR6E/DsXF8SjR4QlJCP0G
XubiX3j0XJBSmzqnafjyboFPi8TeFWjnpoR01a3zgwle9pgkHwDooPNapcnBp1HM
K1OZkAI/bBFvXQHKsFNiNZ4G0N8+7I6OQFz4ksgLF5tpcOtpjT9SidoKE21RCXeM
/RooRAFXFRhnnAMYK+d1r6X4HawxvzwQMYfQLJFdDiTstRzJ6ZZe9NiwLYd1i5Og
/lqzOpKLnfGP3gnwTVWko2C4k6qJQp4xKHWYroL8UjrFc9Ypg5nGyky4OFfa7D7F
4GfRt3xa1/TTPeokZGD2A2BmNOkEsMbKALDonBdr2S3xuPB8XrtXAeU6t5tBlIU5
/oYe359HPYc0AveCJQhEStQ3wCigEv1LcJoCCirOpH4cGJehsjc+5bys6oRkztmn
Y3Oe2IxOH0lASp0MX7zoxzBG6bMEWUtfNpo4dbMTV/MHEindQj8xiBbWfKdSGk2C
hf+D2OMlH2mgLNy2hgTFZiu3kSb8nCfBfb9FOzRoBo8NNt2ksM2sywD0XjUE9/Lu
wWbOZYEAgyNSni5fGGkM3LnhF1DyaKZpRgMQE7N98DHfxyFy+LorRvT65+e1CHEg
W6JXd+BWMQm19LGa+N4BcZ4Tu+xKWokByYNCLlzrcXiKH2sjUEJ30MBJ8G+1sx67
wjdGmUZW15+DDsl5xHeqaVbQUk077k+sctWde/DbRi0aRFbj/FJLCBKrBgm54n0H
+61+QZwG0PmkfoH9oXl8FrqPgJnpZU++C8VYi8/wF/p3EEVB+6tvH9R8hOpzIB/u
R3Ksb3bBLaQwvjEA5bKCqZFsD626XCAtcw2onqxMaEWS3G1DhtNzzOvqMD1gEVz6
PhorIP/NO9Z7/shYAEbFsE2Rm7Bs6uf6NfMoGqnvshHVjQ1dC/smo5Q1uFanhrZT
xGG0fyqOBeBcs6+K4CX7+xm80tiPTYW3azrRUfCdHR6AffUINGVs5FSCKh9Iyzc4
OZL8UuxRroRjIZSWMW6RchDnkjAR1QxZaLnlJpa3uZ/AEfjOeasZaoxjEYcihstB
Evj9468Rvk7PXuzReuQejYq73YTyMukLXYGq7CW3SlYVAh05Wh6EB8CQ4Nogma3A
IUFC1+uckoL9D0AA2cU6+8gTOZroX+twUKX1W1AuTBaCsK2HnnVN9v9bbYrZgKLr
WQtT5ojNUGKmMoWluSnCR5YoL2UA7uN3FWBVjyKS15j20dTzIPmnt42kcpypNKNX
Q+uJtCGowVD54j9m6Sh19rSTlR0AH2drQ9e3F4XjOtN90lFrmTKw5p3fIVWuOTx/
`pragma protect end_protected
