// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:13 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HXsZLP+MEZMKYAs3i0IHuIbiZWPF1MWjlPAn2UpTIj5snZktFmz7gSAJI6FComhu
Evg+8BI46q6oXip7xnnacOhh8QR+t41GCP3inViwe0ywNH9L/eqLSa3u0Q93qxgy
g7WHTIEbzjOtIrn47mHrA/bBLPNonqaMR4FNMvr6adM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17968)
5s7nOxKPmxEDw3c72wq13VxloSL5EtGKvMW4aKXJQHWixR11E1R5rQg87RPz38Jj
Rk98jgpYdkv/J1jw4XXiLJoE189L/avAtisj5RUzzMaemisTL+3/belsapagInsy
tO7MZ8u0lkg6ejdHpE/ygmKbLEmw8gWfMyYyRfnRL3ypXKmwEjNJKxos345IqzyH
gMRxrE+LH89zbIutATH/SYZdoK5ZeGjY8byQ7XzOzA12IjgJZ8obIlBV9VV7KDRt
oFJKlZFJ4onXM/o4X5mjbxhN5u/It68MJ1AY00OW12xrKwESDa9mlBco+wNIjoT1
VFlz6l0NeAPynEARhsk6jmWM8/PnuS5f082dtOZa93TYolqxf2RVasFbsXjYQPCZ
DlwJNIYyrOFxC2Qd/qCoh+v1vnrO/DweOcvEj9jd6g1z1SIehkCZN0EoEe3OFs8W
P3Jx5sLXJ0tjYrBoFespq1ysnbYTJRqByYfJic7kzElHNuaA/qUy7OrBr9Z9BnPA
YPtlZ4b/bmGImmBSlnprwR8Wo0EQvyztF57yPZ6yGlYf/LTeiwl0chCjWhJuUb/f
VEC4gcBSEIUwUmnAr9zsjanltd0HEI0TcTLdPhcIrgFTsfcdf2eY0xHCRfnIDqrs
n3ithxAzAZTqCR6bQFHkoyGOT3PkOndNtDKRT3buv+HhfvB0MBaRtwJqGpsDq3nX
qpebgshrFChGLXG6PcycnV5SU/Uyc8AnKQDk2foUW7PgnEVMv8zK30hmX71aP4Bc
o0zI3veUqKT4Htvhypm5eCxrun9khmOzt0pwi/1OFG4L/EXHcpB/+OQNb+UYbroz
LibFthu/TmhBx/+rFMrFuTL7BXCchb1VWmlw8YryqbXPAK5NK9BFVfLDIYmubYGc
VOaksB5KzfR6swYWk5imog7EV8oBPRvad8BBU7wF7IjZxZvg+pEsSXihoSd00TSA
cnKAEH60KCRicOCsW2EXZM5QQj1wIBHLTC6BTpFX9Lt6X/JTAPpK7CXz2MTxT+er
2aM53kfVLcDml/3V6lGMjNup5Z1WRu3gdA57qpPdcIRbunuDqKcRrBYjprNwJx8O
gyGSIoIjlvF3cNcy2u9dcHX2/YP1JoPNDOcjm+1tAwqGXp6H25rp9WjCrXMtLwkV
z9WOyRfSPxi1Lzu3Jqs1om6OJEJi6er18ASPOcmK8AWyM1ucScuBvHuhH1eRpmjs
RoMvdSNJdjxlAJLQC2XA7z5nXzCP0c1F4kXj0k9URYMi3nYS1g8P5kXtaidlCHzb
OjmQrsVhm06XgSUoKvnxrIOd9kq8knCWmr4QstO7n6LktTJkXAYcUR/ZuTe2vaQ5
IMF2wgUEnEfwD2nnUpHr0JV9TvSC06NVFDoPPnnW5TMIY34p4bQFREtus3Wgqeq0
e6/MmCv2jjxNh9GPT2KTf1MnSkSmjwsKNg5YErP/1WyhH/3GJ6OAtBiFg3Jo0cgA
AJSmQEw+bukmf4OMNZav78BtZaE9c4q14AOS70PeNRQkFtqr1uwuvHMWJWq+DMhO
cYxuj7+hpsI4eoAc+q4JQpqdnG0V+TXwxoEC31rYfsdf8gGG2i+hOzkH/auQBLvD
mxUyNRm6Vh0/EuGnMt2oPMqq6EVQOEso1jruDnyLW09AyFF33GXpNtF157fH++wb
LTcsA2P1a5RKE3YevX8/vzsNN09TW1AIau5cwmArKQv1A3jI+j3st8deQNtsmQrk
ttayyMPo+cXRvkEUSoTxUbkg8Sn3rhOb89l7b6a4EURQXLkNhcCIQnLeBG3rmxW9
ceIADOZ0mhF+X2JZ/0MmAtf/UU01BrcYJ44VD3Rw2os+YwBNWnpcoRDzK7Y9GHcP
QZO5oH8dTyxFuJybJaQgVP0r+CZ6ILKaNMWiy71B8ZSLx+BD6f2jD9XBYrwSqcab
m81PNhIrxDmXy6kxil7iGhIkCYPUpA9pO1ao5u9zxJ2w8U3lolgqsj7FQjbJq/Tz
YTXw+jqCfobaKuiTc+YTYU2MfaTogznCTWqkWh7zwjRtIUyZV10/wtPR6kr5bAmN
7YSg0dcVkhhg9tyakKEOJQJ1E7n0CHFzAOUbd96Jj0+4bbmVLiQk8OMmsyWn/PMu
yFqchG72JUtu9eJZ4RztQj/D6PM0TotFB7Umx/ZYgqARyUhUgHlU0p0VLi+fAmi2
zJEf8iqI1/MxRDHx+5HdtDwBMYAWCfa2DmbPj3m5fYSCJ9kSlVAnC+WK0Sva04YQ
3gh8u1aGHl2pKvV1rd1iommmPe2VTz0g3aad5zyNlX0oKCp6BN44mm+GJzmKCy7J
ELJJ/hgbhdsTdfLXGNitumuzp+uXZPgoDa+66rdec0VFWgi7yTEYwy3IINHwF5bZ
hKoH748eWBebjpX0Zr92I9sSuGW8uVyysONLu+eUbFhKqvLTIjTqKVVdTSjobw4w
EPN2+939UEH6IifVPYBGJNNsIy0txvi/KRbeT1lWNQ623eV9mYyZjDcnR4BtQ7yW
2Z7rLeo4xNW7WRMuaAiE7yHxzQBToQt1K0EZwSob9pMEOmRT56gBCK7gSVzB1ecX
EAbVv/4ibiVXEqyiX+ovR18dfHPzrwzQYxUKCkhZz1g+FC3sC1s+fEgBDg0Y9sx+
reKxIuYlnIWGlchlhW7rZBDPt2klrLMg7YBD3MELVCDfHy927+iU/j/OQvGic/ku
MHfkqkIFCuDXkx6jXIEoAsKGKMkCpfdETW2dLLlVZSluqCE4Tdmze3aZ4dSu/toe
Cd5qbeYAAi/JpVU+ekZyMwFxx2KwEeXEfQbKxV+X4+nPI6V2/O2WhcWXPGFULgDr
Di2Kiu/02v4DJGA3lklM5Dnm7sre/TS3EozL/gYzllHA99wk+FSGq75nA4bKfo1Q
ZtOWSlNr5st4jXpyF3hGUQjN+HNL7jh3aFWa0jh13IUUqcGY9PEY5bR2NfmZ9fDY
ZeAWnyZmR5lOpjRCI9i//e3d9KHw/gnZqtdKUqn0/FCNlf9WY3GoI2bOAHswlahd
SGQg6zmbscv2TWp3Gqn3YDUftPV37R6LuhHr9AAWZ3lZWcZVkqvRbQEDWPp3S229
2ibv12FgZVTbXTaZ8PLhckHUZg3w++a5+pKejUSh1TWr6sZLAyJu1hUCVoEj7Xb3
/fcksuwmU0WFrmK0giZECCd9Wmw3L+UrwxPgnxs6vsgdU+tYVhKBPiMwJasZ3UTP
Fy3in6nElLqvxRETMaoNO+Fq4ROoDPA0W/oPSruJjyWWef+VZNJb/MJvOZB6P7rB
CHMW35JvMi+EQzLDIbxhsEOeGsZn9yzNDUjuQoplcRNowpOgdZho4s3Ne3eDXpjX
LzWgYNrtRxcMMtyJtkpHfARAAgPI2g5SVTPaZ666zOlxAUQvUOXWeS+N9zqtga6R
aIjGdMflvgCtWXYmlwqAN1dcKHBC0idspC2vZCJf7XZwm8LRRGyI76Uiyk9/jv+I
+QplDE6jZsW7e+fAOzBobwGZ5BzfM6UJ6RA1ddkNHno3J0wdlVP8aCqlPV08Uwew
ctzdJ0zMdkz9wgOeu0ryh5o5FA3Ec9hyJKqCbL1fMmhP9VM6MxVyduNYpTmKVfAM
za67GcdZ4n4+HsRa/wzUWlQfojjTY1WRCShzPTL6GRwkFp+widWVz+xaW5AXRPco
rJ8hmOihdnoYf1jjJTAkaN5Xel/wAqCR5ynroqKKJ0ERf9274baH4zwQ7Tkc8MYP
CifOsyHN5yNWsM7Wk99xvNVYnUkK9JNs7AlAzi7P3kTBaDr5SWA9kBrwoOl0SccM
UuaHZWb5tsBaS+c8MR6/0LEQ6S3ToU8s41kYDwiqsNnqn1Qry23O/PZqFvus9+D0
+7d7rQg7+hs3rB00ZILurgGxNF0cTJxEVdrH22BTC86DbV2bQq3tevm4CKsZQd1e
9O/iuHwq99LNYrhoNIHXMFBO7rx7viqbaHGKytH0WMZ0dbdFV1tyijo4pQkyI9oF
AL5Moi+a1nUIo3ZNzTOPJC0TXcedhsw8eDb0Il3aljtv46gUyuLA9LIwHDZn7xr0
vczFGaGvmmMQj9+3AOru6vF3arH8TDABrArPiPntGBBPeX3bacwDK4Cassi5+bjk
O3uQW9OqltTdKa6cSIejkfrMwzNYw0ld+5Vg0e8ZfSGX2++GYPAZyS4FCopAoprG
ecLFErYCY8b2ox0qHkamAoBiRG86+cMQouAE83TsU84XaisNMmb0rYW60R+3WClu
6dyILjb5f+OMHC25IgJYIjVoUfujdmXxgyKG9GNui3DLuywQyrw5qsk6q0C1wtQG
fNIpzFwqnYGBoDaMBMbyT64J+FJcJ9301MKXSeMct/pVee5goroqYTzjPcpKxBmr
9y79rpuYBT9PYOO3V0p79wukPyRQ1pWes5sEqJ2Q83zBN4cO14rdYbxuW/LE7/xy
6//2qxMiYq16+sROAgtndyKzJro4GCAMK33UDiBWtGIgrTMaxWzlqtsk21Z7Y94W
SJN/KXMkcVoWmRsCM4PiMQJVd1bciOZhQBA6C/N4IoLwyXvYSUEJEztM6xcRiyis
mU4mfhWWfO6I2c7MwtlmHwvC/NXvu6vDb4W66Uae1nrqd3ftBadMMZtdzzbrHlaT
WNaTruuB1W6IC+LeHuRGexL1NLTei/j3ib6H9evWWzSvqmYSl44FAk9PXy9xxNn7
pPqRCO9QtDx3pyuBNbAGQAG0WwTtiUZ74G7ilkfEYPAdgbd9VvaDuYABTsWDCbJM
kt6UDg3IBGjs3OL7ChQKiwl6jhbWD7OYBqpksJCz1Eoiwo3mXkZu5ibES903TIED
RYd1yn7EApSjaJJZdICY4Yo0IGtsl8kBe3f/fVG19uem5yGed+gryDRU3ILNlnf/
VdcEqvfkjgnP0Ec21b82LW2Po3bLR5/THSO/fV+Wrqx7TomDGKwNqDazTdBA8+WK
QhCH/1tWji7pDArFlhMb8uQ9l1JzCkJWfgzITGgqscom+CkKRG2PeRoSVve9IgIZ
ieoInEvlV9Bx14TeY2NOAaTK7hoDIGd/X8oXoAX3Jb4NTDMSeIghldq4dIRCGwxn
yTqGgaD2Jkmst/A9BUXfPw2bhMrwPgjTszLlswW36vhzJUILvj+82X0+pZqNwpxG
5QuB1ZPOCKxto9wZgdzk3qu6JVkOtOAtdmuFL/4AiN0AvkvE5NN50ks7LrpF0bPO
YDSBvamBqixTZoOoBcGfdt/T2FtKmYiOg5KW19Db69wRk9lsMuq39WpOwuHEUDtl
HUHyNN8M4JTdmcw5G3yYnMol1z9Oibltn5mRLQ9CF4L2a02kJ1CnNo36uUeUWmx3
xH8VSIVGFdXOqM9o/8U51as30SZs408eiOY1vEO+lClnCQXdn43ZOHZudvYbo/Rg
zAXVkVjKzqRg85+4KqMqBQgpUbvErl3IzXcF/E94fwmiFeBOH8oNtYwp7+SgDwkG
P/7PEdsuwD721cLIJODWn/cs709DJpqGka3FdW64y4Qmz4/01RiCydK/3wQWx7RA
XzkkgyoPoOboXl/7oY6C4umc3MgRG7hpaf2uHvjcmlR8TwoI5wUFYDGzjfRNccBO
2JGBBcCeicmFlBv8hCry3Y2HWYEK3dtpR4HolRHIVFC62zZfg4WJbK2o1FUkqjYb
r2wAq+RkWJP/M0q4KzXSIjc8G00uQimFYM/kAmG7X2SzMQmZjC3SWpAxhgsylRfW
ljB6+0Kc2uASgrtbu8cge4xZrhfOmbBoScxwhT0FBX5zSxTaUKwbkHsx9GUCmDlN
dWVP4LMhBJXzHcI6xcNl09J152zX2NIN24M8w9dx8S9KOHXnd8ufS3wCZ5RjhRzW
JWXfUUf+O1i+IAiSnJfy3BUWkFV3bB/bFptRCn2lENVmtvoDLVfKDqdEcFHkYr6o
bdGf9E7bfzlDY1gxRvXvGKo+1r9M9x/72Y+YswHG/5bxAZim+Pw8TwP8GC5S9mU1
atFYuG/XqQ3EVFYfYXmaCcV0bXUSWv51yaiZHaciDCWGacFsRDMcEtiP3DP2/THh
9v4JQLLatfNSdXR8dTlZcA5h3nTXbK4rshQ0s5OgKuzhMR38psjYN5essu7+Pd33
A9w/VXnV15Jerk7Y7msrnLWoPDsas52yDNyZmKWJ7ZOtPZi4Hvz6Khk5rn9YKpkc
ObcroZ+7PbiJr+YPG/mBbm7MomxLWSc464My/ewjGABhWpPbYXXXZaReiHz0OLPX
QF9pvgYDCSh3kE8rBdM7z6erfmz06WVlTPvFHyKq+XXXEbF/QjNNyishv1U7aZdw
6zYkCIsxNvsU9G69q2sYDDnIoHfEVkqokYLFW8Izr9dGG2d+2AkvWr9bV2eQbrOW
au6xxFa+DGckQ9HDpQTpKHQ1+sI3JcZoNzO4hq4S2aAPuGC/9E2SWaJ1omzCuVaJ
xb3NAXjWshcwJWVWO1NmrSPl3kWzDAJUYMpzLd3Jgfr5vG09i4E4g5t8GmFv/vop
HsxAjJDDI5mRhPuSkwzcVHM57swkB/W4AoRi5+4BuksPX4P5bkRJ41B3f1LWcwYo
EtFa/DNb78R9r3xMm9YESru+2TH531QjAqY5qT+qBTZgKZ9tnkkQUzxPsZyF89+7
KiUKfm931jDqcBq8Hb2NRKqE21uJ+8BNKZiG9O67dSRzGF2qca1V37U40u7/9Yd0
bimfN+lMwAG3imH7GDZS6AZpy5xm0PzKw/F2YR6926l/0pZINS6P+V5lOav0/PSd
HhHEtCLfKnJo0q0QrYRA+VE5cPJcrimL24jzu+gPe7SMWLdhqeTaZ23GBgF28tHt
xPxJmR8lVhgIn4NEaZ5prYubXeR2eHrykV7YGNLzNxPgrRJVw/F0/NUszO9T2aus
KvdZLHqb4PPY3N2sQ53xNCFpTG3cIKVCeHQ1/74sZRqxStDsXOk+oDMftM0FHYn9
kwLqXsDPeI92ZZVmy5zBFoMSh8dWs/L4M5gC6DN9XCRn+xmMiSXC1YIEi5zJX8lz
gts8NiMkSGLkiwN6Aou+MjkiYKnz9G5rgupsYvkBM6ta2g35/xu9j8Q7sX5PfXAS
Xe89U3WNmaEdN9lVcyh6Epwy1VChHgmYHmAE1mq4DDIsqn6W6grXG/G8tp853sSH
XpsKpXgQD6gCICrNwGA5szrrFy4DoJjI3/xdCwUh1uTBUAOeNmzYgVk1Y85CbVwu
Bz4YfTfi3SewhBHpDJrb3xxbjVIQR54BiyX/TKQz8QV4a7cdt3tTUfjzkG3m0fph
XNc1pgOlC3DT//1Cc8liyT0o6z2aE9Z5y4XiMPDBWI3qRm/s2dmBWVCMG6HVtIpi
wkv8UKqBHV8whV6kVJoTwh9IWxm/TM7RhNC0o/W25AnsguYDtrzeOqiKera8ZIvg
vZB8zQgfCTxfPFlIazwXdNH82Su64ncnuo8rpCrIXdbQZ25VbqGXLVnobDbfXoSv
D/l4/IW6aGGXm9Nu9Q3P0/T/giswXE1iOVpghu+aA/iAcGa9KRxL2LbCY1lPVZJw
vSZbiL7B0edQJs5WlF37VJD+rfxCfyH5RFSlkAQxpHtToGHNR9Mrb+jQvIyuEero
tZRbkBnn12hogTWkoA3krke7mxSpPl/FoF69FoMCChTXRtSQ693dDv1NlDeSr+7b
nsSX4fh2d9f4Ef9D3IDqVeFtWllkzb8qcle7SIfvkMgx1ovuWjlCcAaLSV5+IEX3
1E6BsvxiPKG2vBw8kEeSG9kKubL0OtYlQom2+IRvPjg0TIr4AfO7cRdwu+kI0cfi
BV/A1TPqacboT4zFVrYf2iy++kwoXyoAisqqMhL3vC07YI8gCnW1woMPJb3EzoV3
FUS7Go9iiSeo6aSyWrtwfHyH9oJK1jxfFvz4R2BUc/3mzh95cj0zwFZ1rljXT2qR
3ZqeKfRNpE27j+fdIuT/LNmmvUe2GFCYuF9sit+xlzH1LidCPEZlg1E6/DpXLkWH
HjUmKC5QZayWP2wcMCTRQlFxMI5GnuxTwcRgmRXBnr+053zG3lg5PFff9bX8rLaD
lT+i3kbYTOwJwhjCuTesDXprdzya8GBYSqRLwEW9zogGMs+9hCWcBwPxgDkVe+TV
txRLoL3hTO7i66UpTOnOUPxo2Zx6HeEeewHdlr12xJKT4hqK7TPN6I4Xj1ere4nG
xNRuwiF8NSn12NE9486ehoNvpPqzzIkO0KZOjFphGtRh/86um3CGQDjK87NxAtjK
JjGik2of9TDXMOZiD9AyI8ZYFFfm7dZyikianJsixR/J9SZ8y0Y+4MMVJZaKN/FY
eWXMlPxiVDVOhHlzeFNKVVoE2T28Xprc5oqfYMCIBQ5eVqoPwNaWfM5jkZQdzqPM
Xq+bGGRFHvu2THjIGNjXZZnVqCNnKAnp3Oe2OT30SShuQbuyjUJ4Z/JvplBsrcoI
MVmzNj2Eea0xd67RuIkqDowd6+t051WDLYE4krSW0WQJxyoy2Ykxuq3kPbZlvj3V
96PfTsAoD200OeHD9WThiAvAbDcCLr2YjoVN7So57CZmSezm6FqXoYohhC82fyVx
1MDEaGCCfvXoF1SS61K1aujD97mHfd9cAUpc980sIEyvKq1n9Qxk6pzU/lNtZiET
d6Jw+OjnYqPVJn+fdAh5Khw9kqJazLsJjEBOEPWDyA0nolAkGOn4Aw/6Ij8stBij
/d8FCV14kw7gfhUMJw9XKP2/GeYbhEN4seR1U8ymjrqi3FAKtmW0wCYw/sx+ayh0
wvqqkGVYPo31s8xVhF4dndH23TPrKttgeH9qhVCPcynTqx5T0d0pfCE8RK3+pjTl
RVLbMM5wayZuSj22klVIkYLCw0VW4APkp1pSlnsjSzFdPLY27k77fnjiG4KVKra4
Z32NfAX1OmDiaemlldw1sdDQBJb7I2gG80GVvA8dhMG+jpWDAfpl2IfgGwHiCObO
yIhcX0WW0iaA9SgE7P1Kl/e7xZYceya8XHGtYvbt/UH0fmkQSCgZfw/26hUM40Vq
ADtWYRI+Qxj2ymnmc64b/WzzQguDXJUjWaSczgQ+zlhZ1R6u1wGxpVoF/v5U+YN3
HAg6R2kXKEyrS6SRchL+XHC9II8qAybzty9p0he3xFlfh27MkIQh4VlQXsZsbuHD
YPTTrUc8kD9vFaQBZeTCf14psVGm/zGndm5KjSFasRVhTGY7BjT9JN16GmPAOQZ3
FS3fQEWUHp3z/KsuQOivmy7osxZxZFZd+jBNdT4Fu0Fxq/Mr+7OtF1+cxhadrwGl
mgTBnynOVVQ1AQog3QNtxoKzKsBGgZ12LyqdJkWMYzk2IZFZ1onmkWXt9UnBzdmy
HHc0UBoFTH6RJYDZlWQR0VdBw2zhrIMg7GspsalQe8+tDBleE/6aW7Ig0nZ3E7P4
+RNDgqq/YgHlj1R/Gtk9fLZWwCltLK9SOBxA/e8N6OhZ0eFVY1ZHbQHhW23XnD1B
gz/QLS26beeXZMx8QjBpp4MqaltKDiBtfyKXEvdkr/BJ8pxZ3UgbOnOesCBuGrqF
BCyv2SlBrzA/cNdTgDCk/SiZWkwnBHgYQGoyvglKJTHLVju9OBdJtI+qO9cIHuhk
NRxGJTftfBf9saM6drSgDuRaMi9FcRs4m7hlRMgO0C8si2leT0puB/RtrYGCRmAc
q8+L5SEtPOTMlNT5zFsoUXrYjXgGs+/5Euj9p5ZFlWLc0wBmKmb/YUpR/TV1Az2J
g/pUfO0rJWWbAZaOTMX8oQ+DZvcmFK9UxA+heAGjO5/UnUyYVTPb7bHon4W39BAe
kOzVA5FA/gn4lMTZRQ3Hd4hVoFY6GfgqgdOg3djFzVASNCMV6r6k2Clu55a2PRK0
RTzyRWKmQYDNr4xd3cfrGZlaADa7IzlurUdARrVRTXWcgLqEkKyoQ2XaAH5S+gZ/
/Qb3BpwPW9CT32dscpfTc6+by8K9oJv+nWV0TsVtvrzwVliXLYGOQoKzxzZekbS0
eX8Dscxcl9+2nLkTzWgjhLE3pKWCZk4JAyafEQ/ap1mdqGH3Dj8c4UY+MriZ5aP6
a774ISTofQ2WI5KS17rVZuZxqn0+Y1l3J2M4JZlTFTcVWr2P6poFvCBL+vOcSJre
gwx3KJ+yNcH7iHuiAt6XQIwoN9Zn9fNawn+5aRu0t/kheOwYk8maUij1HnOV8jDa
Nd7V9LnfbaO4MyX1G8u28MhBZvZvTuDQVXSNDpLGeSpRyq/K/xyQnbaVm6oIFDzQ
ppO1P0uPTen8d4lQ1LKLTi0rkHr2k7zvXHy6BfuSSTMpOb4Vu6VuFDnJdBY76BD7
Ad0yngZ7SCBPpanih7w6cho4w5Qj5Q67+5tsbhDe6gebXdj6313+BOcGPKgDCzkB
KrjQNBkmFMyVUY6LdlGg2ohjvWpKuqRoUUWnreE492ReuiRKSr6vlc75wWsdy0N2
o3bXsbxer1bB9b5/3ttTWCcjnd/bmbWQVJ0LD5rhTod54FTzIIVa77da87ZBcadP
yeA0ztwVqV8EyNhDxS0Cpdj7DvqnR+2UnU0N5RqOWZv30F+fqHctr6lbm/N+wsA8
YDtRipIGqDIKhiWC2VHcnwmVKUv8XNMzAwJIh9BNjDsWFXPEuZNeTZSB7wZovuOj
tCfZaS9sd1IHWhCElGhEpS3RZ8FdEtq7OVampnUa5rWqzUkyQ6nqZZlBM9JK/ldZ
FM6nYwT1O1/7z9Y8HPfNAzDHW6i7qgNh7dL8neovUkZ6ERtRr5BQWBkPZUse8TBk
4HTQEcg51UVqDIZ93pLUBjRhFWgE/ViVhZuH3Kbahk0cwtDb+8Si5f1mZo4v+uKx
F22ZS9ENpqJT11fuNXLhZ6NE+MlXfQlS//m22KWbnadr+m2+I5dNV39FfLI4Tv8T
/3M9yPsWPAB9I6e2g4X9eNnbx527mVMvCO6qsrZnJc6L7NsGFfyWhTSTP3t67Vxb
GV4eomCsIpuBD1PkPJ18WCJE1Kiwv/LlLIgH0UvAukK35L4pYpp5Msah6ip027ZE
qXD46PBPL/ILfsWv+5SEjNjTbDMuQc+h0SS/CPlfhPgUqUaJp9BVy6+TSe/lItG7
ouXOBu0Z9BSS53GhbVJl48gNtfkj3HPZC0EGQDd9XbB7NChRSebe/IKtsbvkw0Ea
sUPQtUdr3M/WKOgljxMN5UBFRvwXhIzQINQse2Ml6/PH0BshBQ3dUxTyUAg7Bmqh
j116uGUBSrascz1STZHeUJepLXhSXsAV7U3Ci1cvFzTQbuelX5OphJMRvzt2E6wN
xC/j/Zs3T/ExM7Sf3ZO4Q4aHsHO7LweXg66k6cYlEQyhDUmfV/hV5DkghCsvbQ1x
oWZUIoVXM0xYDUb+NCbjxriBBW5+ZOMv4/kH4fsGdxr6KeGiYvBdRINc7fXE+AQ8
5OqneUVuuWfLLcqnWt/t7DnJtPvmx8ULbt9UvqhRpi+9Hix6DGzHboAPHQ+W9ZEA
rYYgGhzjwBmqLo8hjw2jOx5CilDaMNxwnFg7RTN9cZ/8yl5Lanu/TOgiLrOcM7Uo
bYKR3AwUTzmqyanBiiUpjsuK8F2rwzIcTLTc4MPCWT3xgE6jnbljNKqXKwePe9xb
s6wjxgbaMtfHUIn82ojC1b1IvPge2jaDuRPSSNN6ciRJbjI/uKBj0NgEoE2B7oc1
lj0vHjez5PrdD+tYa0eJ0vFpfLU248bKEDCpFd/PII3VC0deiUWbqhQkQSSnmvgZ
0h0q138EZjpzV2Ux/gqcEg2bkQ7s7DKON1hfjapzQOkRwCzzQRQHwUZn+drWyHIe
x2x6HmrrKS7Tc3Lqf0H26oBxWAsPLplqw2Os6v24n0E7kiQXYoQ8yrwHZyoPm/gh
b6IUhgWADKiRvcu16NVcAo82guj1ZQ0bTiPGvUEcV3D43emjJ8+8mXFvPmIR3xwf
+d5BM2FM73tlDeB2Hbxuc5n4G78k+AbKFskh8rWVwu4KWM7wg1mcP/blrIoHYhga
nMC02joS6V7gLdbM3HxH1m11p69blppoLyBC9EWLD28HacPbeWDrpg/74H70I0PY
w/tj01NpROmMjF11LfGVBpDeK8C5vzAqjKI5A5NAQ4vtyCLU3HktDdtUHFRB8dxn
GeXM4AU8iBlp37RenhjenIR6UE/961tdHPSfulefeClkmyMbYpQK8pYbcrMHufZf
k2tqxtc57yo34A4fE5ISLg2SDRKVZrKGFLLqFIA8Vfs8fNJK3PMEPgg1uGKO2Jyx
Esk14PSPe7fi5hrzH4YIQFPT4RyfBD9iiH5+14iawhwUYeocWVRxlRjNLCOYp0m0
RTojVgUab2SvraKkqTWJlvfQ/3mLxbFygalsBgYh2Hng+hQ9A0OjXjdjE/CKT1Cl
Al2p76w/z7dOUx5nGXF7UBocIvvZGqgD60yt2ui5F0cISv8HBrZDpXUKdAciFELH
gs/8h/xRkndX6q5Y+4hpNSPZg6Gc5jvzis5hxFpHR0jldCRe/XCUgkezmJW/EpBU
9KHLLFOOwih15yups7h+4MfMzYMyicevb0bUyiKs2MVBsIB9uAutf1DnrLS7Lbas
wBPlVPev/SzVopIoVxiBckXtIjVmLJX1Aent7PM1oTukY1xW8aEWZ3BHeh3uFHM+
jEnH44Ilt/TJ+uEmQe7istFS0jaXZItrh+9lFacXWDpa+zGLy94FxFYEisvEvbW4
txnMK7oAulsEu2fKF8+U4jzjvehzJScxrFKBCWL660DUgqC2bPTwHxIEkV0mtPdu
PUuofXLDbYuS/GY2huaFyKB13SzQa8gTW39kwyuSdjo5gKfI8JDPrpc2tzk9JyIc
UCYvYR++oSGQy6vcYtTkDo4ijk2EjhyzSGmxRcVOpTO0BpFfE6D0CsK65ZeFamoU
DJOxN5a2MUcg+j68PRv6VN1FQ0dDb0BxOaP8VyulREPivIEWJHVn135/oGdztNcg
5u1wlziO4hUro/w8N1kYfEt0mmwZD1+4BBizuLXx/II8t0llLGt2gFgiCSBab7Cp
n9m9NN6J9kYViaX9rkAy7WWLEJn8D1GmY8zD6SvLuA4GQJlJcIvyTpkn3+jMpfaH
pMfwIbqf1gmbRXFg6lxC3NBHFg4Tg7/pX+DOKzHU/+D8nkcQ8Vv4m9rWkPplXTD4
PYQo8vgIPCGbrV76+ogThd3kCREFyQ9JzJM3LXHalxn38KUGsPA4zH9Z+HH7etH/
x7n5pD3pHgkKmEhE6559biGu2k+FxO1qlOZSU6usgRtciITR7YuYKh+cM0q7+jxC
XpdN0mkhZTThpd+OEyqxh7yP/BP4Y7KdMffNWbUTkS61NaHJfyFeqBRWVzF5vZE9
NBp4gZGR433XuhEUr6lbFwa7fgtHecDnnhwZGOL/dhsZaaLFnX9uOme0vcGY/HfZ
TafyJGt+6Pkqh2ZBIHy2Fp5jkXgnLvYG6QJ/9+Dkrw0UHK8pQqxa2LJdnhQhT/3p
Pse3eCvk9jHWmSXG8dhadIdulZ433LXas4PZGdHPqjSThu8RwXe97Bn2ZtLSs/s3
vukIvYzHXVmMOmVRU9eiqgHn/fqa1k0UX8bK28Mc6FnH4aZt4l/BFfarlhqb/ClO
uyTUTleKMn9ZISa36uBzRT6qQ9i444IPJlSbEzWExfgYGUYgpoNKOwVJfOSCW5Yn
//S9agI6S04chZ5zvB9gBQEWB01O9EzpebRxxHopjK4jZYQlev3oAXtpEFNlLoHz
85LEcSeDvlVUVJ6Wc1/CFma6t2CjaVH5PQf8ysypSwu2cpyp2s16W/TTqSR/tDSU
D4ELYmSSmmez4YjkT3rHFqvDOGpZD6dDsZeZYOpWHeCJqHSMAQKlPd4/+LkIvfFA
j4V6IAj6r36wz1RMRZ4xdVfkRfvbrSu1Vv10twTVmxf8refHX/lnNhDkQF4vT2oU
4zgguClFtZb1T0u4+JxuYLwitqoOkg9zgutzaa9LfCNJJQ9/brJY5PKO53hFbYgG
B9K7b4A6+V7QMJE3xuTdaB+AA1eGV78q4vp4NRcPpd9QIil+c2Bs9VhbzfIKncaQ
aeDL+wuqKp/t9DVZqemyWRsYrNPu+nVFj9pjjWF5kpO3Ak6QsiRl5a0SolEkR2/o
qqOH9Fcnxb7WGDAyQf0sWQbC5ESPsR+TxSOyHhwNgKWtLQ+Kz5CZSBjcLTjbx7l+
p5TPF52TYbUmFK4fVYmS8ZJ68GmMsnmToJVdZahXX5+iUjU9fBVLQ2updHKJjN6q
tLmNsKl5iWUTM/a+oaUly8oRvywYYQsPOzlYJk/azo+4XZwhaHYm7xxL1h6FWXzw
Q8HHahOM9jDekzoPZ4JKIoAgRyB8e/J4XRPFv3myfI8HK39hmIwvY1Wx20f8bosh
rYIZJl520gYMraUHmDmN5AoSpPJJMR5E4gR6eMeDr6FNGv/+9LRV8EG2ruspO9oN
cSAFxb4fAEHvR3AwXcv1u8x9IiGXKCApCiHBDnc/CylEic8aELeYVxpvBSIGc3lx
DXpQob0pRoM6KP5RGk2f0ti3x1jzGL/8oh0LM/ux0ZfDEU8frBZ7twSiW6vpq2qp
bK7AxMojo1cukCIjjv6W0z+ihDkXMo+j4fWrHcwzLe8a7VBRbwse65pnQrQ9Ztry
bOvmeIV3ZwFV0aD3mfjWrtQuQ2eufpgEcntzOt6IGwJseUT19rGsMd+aLOzC100d
YWIAG4bnnRBgyLzUEg6paq8jYIOhJXErVYQ3LMfWC0lQdLqxF1ITK3ouWxil1twL
KVcjGWqGKhwellIlR0zSyk9F82vIIrCOuP6F4OFR2lfpRtCsTlxpj/I8SqpbCr5Z
urrb3VhbIXLWar26DISd4UQZMmUnucZoix2zx1qr9fDJu/HgCU9CBqTgGIB+L9B6
umBIhmvytZPsRhPSbtIkP2e6oEU7PyrNPa5ydx52nkQeSCfHD6nbJCtW6cMETO6L
Oq390+gCqWfhosiTjydjkXNJSNMjjvWemQg098ul12zBb4WWH/+/zLanIS97ZmLd
ZPT5/e/wd/IhbphzVKxdlSaXnZpr+YLFBbzOIYwK0twyMIOP+OCDuiVLceVBcEfK
1FPJYFLzcV1W1ywjvmfs8kntmAJGrg4yGJqj9sHj6izr+cqzT0E9CZo4hE6GuhZB
3cdZojJ/IzSHGMOZowdlIOa/q1wbAczHc/EdaD74+J8y3NQvzAvWGrYRXNnfqqTn
AYnQ7Ez4ZHx6HNoxRmIRPrQZXeaVYU4yubSQxBhA/nJ8Ng3+5JOFzk0aGQPzTISX
N/V3XUqUvlsMMOsqxspp2JY9vrGfrbaYt9qAoNJgo8RZoA/os3+n7ZEg5SbiYmoY
H3BKN+VCQrSQlXIoH8SrT7KT5jDq4Hob0jSo9mk+qClu63D/umJSfCH75CCGlwlN
Ijw2B1+NyXd2bMvseHKro0Ef1JIfz+uIP8hTsZs3aQvrhlRk4gPAn9pRMd5PyOhT
XsJBiHs3HcKMZE5T4VIEEWEb8VSfhaoIdBEYCwVScfc0t6uj1F1G9ZyC9Rvht02+
gug2npHeK+sTnLzIrxE7S1CAg0/Amy73mP2Uh3K/8k3/mONRcagoqJy8870AsScl
I1gMWdXi7x0+7ZRf4QH4oHqwzsKaAsR4iC9MGLwA4eBGIX3GzqpEfwqx20UElSGk
AhDpJnNPpP/wuYNvABuGig6kc5juA8NBe6BTDIlBlqZy+f7999ORXdANFKu06bsU
/q5943XCcyyuFnCB3xMiBsjV8YUVx9E6RpzQ+k99HR5SbcIglS10FAwR8BMxksM4
/uTQrOH9u3hUpdYbgElQv0Ta6XXJUVyBnbDwvnVAG2OwTtNMz7efp70kqTfz0hjM
CXOzGlL4gaes1MuYpzZxXqBo9v/U7u918EgNgtluxHUQIGtFq3u/SPKH+xJyTaex
2hF/Nh/Pl0kCKXZg+zN4GLuzfJSxIjg8CugTuNAok50JU/40K6Y+GpwyGJuYxVl1
gxQuVOq7UFYE6EW6AelOk8JbBKcID+lk9yUuh9/gQK8Pt8apUafbUUevQ8Ndri1a
f727+2OijgAIn5xGOIc2SMoRJqk4HhileLuYA31UiIBZYxmfg7Np4mM4/et74A94
UIok8VDM+Msjg/QBbugJGmsp63wqViqQ75k0S3CCbeClcy3kWLBcr4etYDRxO8vB
xJk553fSoh8365jofwyMl2NhFdRzukeF01d+6lu4MnXxPNO2VOC+XmHHsKRzNaEs
k0qfL/YhV7/gw5X4tDDNtBNUnJYybydBlCvil2/X1AcJokGe77KF1/30FgmQsTU8
XRwh5qGBD3mKzgI17Pz4Tfg4xVgG4xf9rYRdbrDhxK8XF4mIS1fZXAoRRhvU9vby
UFfmQkBqGlpOrQzdyORxt6czE8rzrSW2vBq+tDZ0VDXkZBWvhJ1d1eg6k8O+xLVb
qc+30x9VqJbk97i9ufI1YgAvHOoNWR/6qA7TNPZmKat0km73I1ElLGmO8ODpKSXP
QBGLZWZVITigJBgmzQtC8lpt34y6iuOKsaGmcOc7Yx9M6Fo6YY5tvksAB0z6yKMh
S3YSCh46o79VXlI4wTKTpBq1VaL2QN0aPvQmjShe6B9HUS86zaqzBh1yEhnGZFPd
1QY3mN5Vj9u/QsSI4+fmuTrquuRm50eIoADwscGEbOMhQuMVBnkLd7uQ9+mCICEn
IBj9y3k/3W5mjlsyyo+4HtUUj2w0mIYYkc7Umls8geHne/ClFmjo//g2nRrU/K+L
xEjC+cmC2TZvC5Ld95njMvlUkBQUZXzeHUylLABdEG72sF0GcP/kiXzHpZhuhXte
UiTC5IPXQ9PctIr5x18hj9//nYBX0niugUEzX10+PR8Jmj0Kw5mpsOqgfrpKV/D9
MMfipfqat/eTuGgnOEmEG6tqEUQ+PG6u0xq6wvSA6/EokTuEuEeXNbNXJXUDAQUj
lms8GSfLv8sZdL0nv86tkvlksl1CHhiLGUYJgZcDoKNrJUl9KjwSqhsFiE5ESwoP
zf3D/Y/Wy/olqZPSjf/XFwSnbl2Jcej0N+unz/ruKBSzzR6oJVKtR1ErYYFofbXi
rIpTvxWSr3/+WQDBeB5jl+Y0ecGpOYVLAVIUi/krblZ84chjWGQpyMkqS/g0vaNn
Tv3QNM9nsrcw5im6p10FCP//qxvq79vcsJcfheRdIW8nX/MQJVuA+/ihXFqTs2kn
CGmQbGDOUuQbji0H+2mLbhEI2tsd2/al7swa2Z0+ooW9aBYPSxlfgAWs5V0rGc46
LvQbnKnHNDgJOiAKlL7sp5qvChoYsDBoNPDF0tVa+DBcI5RwdHvGnAE/33sKm5rI
nS2VCK6Rkxv/6GGFQSQCYWhGwVdFB1HVhfH6RNSvPd+CNMksQVFaUAx7RvTlmnuS
dv5TA5pwRREW/w7D2hlftbUse+9+UkGNyMvabvKD7p4pSh7iSBUVKQLvDvJ7hT9N
vVFs7kj2rnmKrMlooMebvn/spA9a3KxTkBjkEzSlUZDa/P16uOWu2EXw7PEYdtiG
1BxO8UkCXf1Q3ugW6POW9iPCwq2YXh9fymXxzy+T7qEVBD2nNmKjKIhlaLWo44WA
0/PF8i/X3BfrnnkH3KRxiTUUxMymYhI1eljV6cuJsZSD+BXSJmpbI3Of9Sw/vz2Y
XHabWYUEhn+xtyYeuma2J5LrQolwJV5kdACQ7dK30ityXfJDSAxgbdrZoOtLThiW
Ge+O1JihrJ1/YdYHhntW65lo3Ifebnpp81UPtI47ZoLpaNrdQevE9A9hoq/elfvN
sF62lAdZU4BLYa708dGLo9+MT4XPcdLffVIh2tVzjua50Sw+CBvXJOHtRPCx/WeR
kuF7JLxodFrVCJDxZFuApcJ6Lpx3UFZicWlR2gpDzp6zH0o7+glij6L1y0mBmD7W
wjJZK1i8YGndgzVlvG5inV4J+4o+Y1yPQQbAw1h6sIZkN0fHHSYiOFzEvhQbWr+N
lSAxl0HEV9xr3F1j7akDrhaw2JUZi5CiZvVPCD5+b/RamDtR1dVDs6hjEHcuzJ9K
JLHTrtzVjG1O+zhKvtmV/xG4gvIBy7VpQCwd0c5JeabzJMZpeT3ptq8vse02VOwU
wnu+2nT7fnlDDwKjOo3Rzlz8YGvZxDYP4TEnY0XMr4uspRO10V8Deu9cUjwVCTE5
AL11UaIkWC0vK5UhAxa8X9+KKJsz3/r4BvB60P+9f7K5a7wOvlR0GCjDMDwkXbL3
vAjqbxAuSGsZ1dZNbB+F2yTt5Vzvx3VnXKJGmNoKNYU9TEX7h+g6ZXopi0c83U9S
hutE0rRqhkZ3dYBM34aI95ja35YuAu0VWXuMdFHKPVWzqRTWgWvTgr3GrF19IYQd
kj2cJ/WSjV2Z2evz1tQdiA1tgyAKQ+AUPrNGgEXWmWfv8GJdAB27UJjawkMkg7s/
Wm/GWWJcPmfyHTEiUaXXseViddbZ15EyMMFodjDdVBHgGQfuSDLn+nf7BCEknF9f
biN/DUYvJVcdnQi68kZsMgXk+hrbJYhgK7WbH4WOH0nxp8OXt+vgk1QXA6L9dCbl
0VVPT6V3wXNciVmr2rz5psGB7JR4lV0TSQWsU8ZGru/UY97d62s8k5+y/eGXFa1B
hmhJ0KaGa54JbTtgCR/BDRlmr3EoMtQLIuvRlTkydv35/oA+6vlort+zd2Uy3CUe
DsP5yAaoq0rQQ0cTFv19czFjTLN/Hpg2prHhsVW7DP2QeXruyWjEJFZ43Cu3QIbh
AkjjFJHInpvAUfXRPtxxfwh16MHFT6lTVwOu90JjrZpl3gGtGfMe7r7CE2iI6kCJ
JeXM7txR3vIPShfVKLM2Y6xv8m0VMuDJsI9Yte9XLsObkMh66ZZBmAenECE7gEas
e53Fhzi5siYTHcjKiGyFR9L50TORn7uUj06i191aFleak3hOvUVoff2eGL7ntD4H
+9pw4BVQ7SiRmGTEe9MLTFkl/UbhqgS+y/5Tz3nOz+mTtCQkXW6lhaPX4BAVh0+I
1QYNyKLQQMXw9XbvKFcPKeWPfdMLJM3yRb9+ZLrhgMlmeDjJnxiY7Set3p0B3tUZ
coQ2uGuD2jC5bNeSyBLebKPrvaVitnyy3lZUSMNaQ8rBgHI3MRPCd+d17vxyPYpb
q2yFpr77+BmeRkhBKG1YGIzJiufMQhR1UEspOBvnNgXwTZD/gz6VC7b/wf7RQz6x
rbAdTJmJZB6u2LZ1xpRs9KdJj4QeYlkLG6kWfKuxasB/cfAD/z7IemGiDEPdpE2b
9DVp8QPXdlgAqxmhcSzfUBuG4p8AH4q1Sb++7qcJJaoFFlqSAKHvsARPzCYg4nlB
HdDuHexBjoWZLA+p3brGfrbu4XT0B3eOvog8IacDrdnb2xFahRF+oloClgKNcT1a
PfmBM3dVELPtKnhUcTaEKALbIn+EVjPs+pP1yv5/xCOne2qI8n7iw6SCzfjqvAfF
d6baf6Rv8y/Su3fpQgqOB5wFldc6rnSao3pLUYY4moz6yu1jdSdO+RCuEecSp/ct
J5bd7d9+TH5BT0Ds61FIopRPMQgmIsJHIcAgYZLz3El0T5SWqA9MKu8C+aUizn+B
GrB0Z0RCKQm9pwbsbLlsZ/f2HLf3slO/J4HSP/tRGw7OWzDyPgKVzahZUW9bBsn8
iF3BfrQ0+uAfmzXIQRcFdw6Lul+KkAPKaCWyQweoJ0AL6EG9NayKryqJVOmu00hm
Y64eyH/xcjezxRpSDFzwp9fqVT2NwCKtPrEO3r187QCU/RXjh3ovdSwF5RxgX3fh
qB7LVwjQbTUVC/+GYx5jgYAqMulHVwwTpS5aQYheA6Eof8lKXrQSxiR15pQaWAzy
rLlqNud9LLkFWAQciv62fDHw5/6w7SkTp597urKPdnwW2Odt/s0hEVpsSWADVyN8
zw3srIFq3WT3E1KXByfv4q1pVWyX88+rA0j5JAsDsi7xn92RV3OJwztpFdRUBJNN
oP7csn9I0WJpp4g0i8pztQzSPQOl2A7ETFa28sa01n14X2JP+SBXtxRYSrsK0qKm
A0d1MHAJl+nQe3yNR9tdJe6o414TmMXXYdiDxkd8B/uun85nw86yFU9WSMSToR9R
mEDjySRKnX3oOQFB+YhET0wNYlOrvMK+w9sdS2W3XqGpJE6r9ZaNLGAFn3I5xMwb
I+3D/8ZRR/bIYce5Gtpf+8Qtyz/+u76++xlrDox9mHFKNcz341vUfmFPhJLc8YvP
CpxBDZ5awxp4S21q8nPtv8kWw3tgM77pdGO/MeGnQ1hXwbblN2G3RmS1C3eRlK2F
oiyIkSSdOcsQVq5QHNIiJcDbMcY/2n9AovFJASg1gLqjuW/+hyjYnGuLHeyXxt4g
8I+5bY/+JWoHxsVXXa+8TK+kF8IR8x/KTrQ1DEppZfJeMQoJmC5iTMksy9Eb4nYj
ZBokKcPMQz5h2PKUT1XSWwfmpV9Va7SynrpY1hlNseg/aJsYlKnRWC7dk8t+7qf8
/ABvwL8LBYVvLBMlYQLuYYJHgOkIxrddc0NTaoy645fTZImMaEhkwjSga9o7A1Oz
rFnXXSsOpwOqRQelcedA1L/R07KAktNuX4fj/FBZcSYX8SgcE63DIZ5GdrO7cg89
cs4yiMSDubQ8qKDTnqEE4GXBCsiqsmDP7VhHXRqSoKVKLuqmCrOG9HCCMaHkpnIc
8EPaKrt7stsURNhiMIbFaA7hgLAPBxxUP5PtO42GC1H+aNVl2cmWm8ht2iu3ulTE
/OW7OwTEqG0c4v/hfkA1vnmlQMdNyCPZIwCVq9wj+uCcg/8SY4V/aD/SQySLNW3C
eboFCjVw3NbUata1Jt+8CPOn+4OCithh1KOSxblL91JEriplboXhnF+Um5edlvFC
63DaeyVKYhQd0LumfUd7p4mW0cB7iuL6yW4F9dIZ+jVIrbnNIFAH0WDWrNm2cCsZ
SV4wkP2yixfk3nhoDxxVtJYWpq1WE4A2RxOMjL5hqAw15dI0a40mpjCOMqIISdAj
4FqvSAn+ur88/Vl3sdr5JpxKkf7crARYV22/0KvGtigfh65lTltsyiGJI9kwt3rf
CQiflsmYRKmBuKS1j+1lijVBDV3OwRknGspQaop569ZiZFumzWTAyQVfOQ4paYOt
ecLiq/NNsMA1GE9fwNXSOx0abAPCYAQchBeHNcoVq84/UKKUKjFWEXdoGGFTXr1b
JnBi4QA+hak8e3QszIqhJzxhGJ0sQK9bR/8t4nxA/tg8hsgtqU7oZmWfoM6L4Y2/
AoRUB+G1M0XRRIPJvXHI9TNqMEzPopA1VlIk+7AOhQ1JvsiNQO+my2G8xLvU2Yiw
Mb/D3yfDHLrjMKwrcYomo7VW6LeiWiftydzBqiypAjFbLOxbZBGpMx7x40Czszm0
kgmq+D5csNu9LCWJraFNVkAX5DY2euH6iraIGuhNkkmA/Ag0xQwhgZE55BFQ8RGp
X99EdBdoiBP0pnv2+V+BCpE3PnpMOdSwC1L+zM9169wqrZoDwYwOEQsONPK33p6a
iHCCIhZnjDa6AyQkcaHiL8FUBVafIx2l1tv6G+ei2AZhH044Am1ylJ6IP+lJpxhM
UGFx0jFTkFrP+CYJCZnJs9xOPZmSX+2Kv7jyrsDUlEvXroCo0Pt15dvzmtjOo0bE
0W8zuZeJTZXKoE9FBVhtuuo+CX1NtnBQI11xiHQsK4HG/O+5JZvAyo3eix0+g0Pf
G6Ee5cs2vXgpk1x4KAd9IONMb7qoK7kr916lQE2iFVHXOcTqd4G7ZOty4CFF3cLv
BuAmeu0esMI07ebs61XTfey8IJv8NSxUli+e+7DiJoFvwhPdfjoTB+fNNi/Scv35
+uA2ANy3M3Ov1NtAGa9zbXFxmRuAd8Mp8h7QBj1UDO3dix2J8q1YYKO0m6REultA
oJP+SSPRKayUtPUmpTtqDejSJnuBZVOFo9oREHQuE6HxUuIdsaCOgVZx8A1lncPA
U1TNRYxk9VnS5TC6BZzeF90pN1E0wNohTId5rkymmuuULoHq37OXEhmUNLb6N0W0
R3wWChYzrZL1znIzkrCS5O2fccaN950HA0Gjvi5rfueEQDHNuInyV5SFCIeeMAPQ
/3qQV4UOJEYxmkI6uzpvTcE6XXuJsVFaKM/rIGUirN2cGavJJfB0NOrn6s6ttyla
BpOUA5KTz810T9UFlbHxRwHaNj0jPw/GHWmJCJE9yx6uqGMY8FtKhe/IzHzmf207
6KX+GjmULmy6zyCF5LWaEY/6VrguT8aMS0sX56H9aAHYTqiy0uBrpd3nUbygTcsS
JKrtez14/89Tcjlsfn3M1sYNqMb6S6tqgMa4kM6kb43+LRwhUTpGjEcMH6UzUFYq
MBSiMyqfXfy6ZW0HQgoMsw+1bQxKsl+R3nnoYvt0iaR0dTUTYSMBWbDWnhQwukCA
OZcDeHdvMfVI8TKBgeRk6hH2f7sDkOI4Ox/Wtd2l/sKWQFebSbeLV8wq7TDrx9CO
rmEiWGj8zfo/7tZIZ4mujbNbEhYOEnCbHCsPeeRvQQw2WdLKPiVNS+C8jrhDIyAC
yNHKi/7JWC/RkA588UIM6KV146mOV06gpW0Rn7we8LaLJA+oI5RVoVYaoxHHseQS
sjhjILPlGilKrwvrtQ/j+Antyx0ufwhmnnMdIVQmDsx3A4bvslHBbm+jemWSxnlX
FLYUTjO3rCJAbtlcMYpf6w9miyoBBOLdo/+NUhLv07W9NKemcOy4hYhZ0A/wKl3+
30HvWVtEjzIDBDBYaMDjSJtisPVUt/i1tc9B3MQ47YsYJCx53HZVVWdiFGTTwDLC
Vtpn+LJ0gNsTRA/FnLOT8eIa98KXd6gYkOiWaVo9EJlUkf7RPHdg9tGn+iQIPNj8
GSgWyLysnSEgrguN1jSi5yz36I2QYKIE7Y9pZJNsKpIJWuzduQk4eEFWD2mmL2cF
YMVJXXPxMmPbBs/ZRWsYFsr8h2WYSx1Vsbrch98lUozCl+uFMe+sMXYQIF+sq5E+
6Sk0gpmsl+SuhE9WNEp/jhyIBxRCCV+44WZm672JY7u1XHiYBzYV8cKjx6c4UeNP
qYNyYWLwWWF6bm+OrB42Z21lMcLhNxm27xhkBhbrWSmH6FTGpxAJmgKDNVRXoakB
RNztZEnQcuwTLMb4+kSuaJQChv2tsqQpj/5eCxMjzEL9G5DaRhXpdxgMuIgvMgUW
9Zy+dSQRANPbMV9JC6Rya1V0FaKo2+MA3928My1vy2ly07zkHuYXNxO2Pjg24TRo
wyeKpM4sZOoBY8P5ePg8sZV0TuaqPudHnEfztAPGoGbO9zFMwm4Xu6QG9jP7eu0v
lKtCzlLmyZR0axSP0vQuUAnhtujZoRUgIRcGBVkoJVYlvVpdKJU1MChqjCp1glfY
zqVdK3yciJtp6X+RiEW2ZCFPJ98ftL8DPXmdJdVtI1DBRLzyYgZUbgIPL9T1lhPx
y4eW8twyeNOWCu8u2RsTGoBcILEoJo5YvxeNd/It5RQUSo/G13YRsFKwGOiV9BlT
Om1Ps4ZEMUNxOUvPiSq21eLwWaIu7QIih17G4L+ZR1g1uSI5Ehy2LMRSCsBtu9SP
KlmQd8Uo/5Q5/VnUcro5zBwXBbydrP8AGoqLHwvrNfmuk/8yCJjxG+WvPL8IrduZ
pLt3IhTfNXOx3WedIBKpcRnY+rInmH90ESmqdxedS+2Tqd/tkc53fsGazXVt+lgZ
f+mWkfNf3FhUAWavHUiDcUPcitY0422KJrQZga2xumIfuObxd9r09HGNo7okBhdw
Pl32NYH8jEt2spYc1gzcg2bQXNh/4nsZ0dr4/EV4VRJsBeoV9UeCeDQVmQ6AOFLn
Ats7iqH1YyI2iwurVQG//14KsVb6LxJwA1QJSoNxydO5PWqhAsaQbmAtV3P2Xqkf
BIc8gvue6CDHponTtTZuXkS83scUGuzyy6qi4RTZylVkdXapP8Ueo6fuap/l0eIv
hjAdilgCKb+o5VZPZcmixOi7T7EKRiMGcCfgrmpJcLwWMKrmVrmJ099Xvqa6wg1v
VryhKG0UnbgHcnzDrQo3OhXY8HzM0eak1wXhhFC9eyrswqv5DnOChO3AhMF5C/6I
gOhW0maVbVt6DnefaO4iNg==
`pragma protect end_protected
