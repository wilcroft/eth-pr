// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:12 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QZ+PKxwU68Os1ia1CQ1ooz6o0gvsUskM8lB0n7Qtdfe5fLB3fy+RiMeEyz/pLAUw
KcgSTCCb2ffutt+F8ogWZzTmkRD5q9b2v62qgZopUi+hLlC1sIK+aSiY4DoGigRr
dgAv9GdLf2x7hFb9NMezMxk2Repz8/xpgz5czYR8qQ0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11856)
6qrjSEI6OdJOzkxFZsLeT1yD4NcM6IjxQYGTkeyUgbIhoeUBv9915I6mm+b4Fiu0
e/Xyar9uZ0QkEhP2FU4lIM1iDO8L1XVB+2VFw5Bun/KjWmVMjxZ6H+qEJQrFFdOA
yM8Yw9URBEcMUPHHXVue8To8dJTpjfB1Z990PeluwCLLm4SFsZ1zOm0u1gH7CRW9
ncr9pXNxPo7O/CuKlxi48rAkUpknMZyFnKEhsVMQN1K24fKncTbjl4cMe+fANRsm
xOBnL9P2uc7rBAEFZTgI/UDcoSvVuVRqvYcd4t5CaHX+90AePOs2sjziYElPmG4N
dEuNpCorKkcrRWQBIxucV+LrRmWn2HiSjs+7quDkPqv45n1x0P4S1EpL1AkzIPRQ
Woa4ERXVs8fTMRKCeTsSD+v0weNriEV6yjmvHyPW0BWHgdqJtRMp+mfXDDdDXBQX
Qa70w0VWT3RNDY8vrrDKoaLRD4W0T2E3jefP87bNRSGuRJdjiYYJeqC41Q2ftKdJ
ApoqXAl/iQRKifS7o6kqJxnGjMz4xrHpJEVUd40EnPjH5zEjkzAMgBNv3W8EMspy
Z0wD1i/n8WFMU3nBkCtUO1dnTTk+oDK5OntlrOeU613K81MRciQODPqZe/Ek0gAm
9iE6OMEgxx2XUCXAmu+2U6lfIeDrxlC21s1vE9jtHha/r1dbbj2EG3upcuGpZ6Id
BQ6lck+2plTRdX8a3dG0rqpDdjCfQY+CK+7J6nhjay2NwQE06MtdirObi3qrk5EA
ehbTkKFjHc7VAWrf7KTB/xr3jI+A9kjr8S863/Dbrj0vH6mC20Qi2oD0Orgive47
srHIG+Bt79BM86mxuZmgxBzGwGX0aCU17LmAvYlanRw+mchRVPLsgxASY+P93k61
Ook5yD/UKD7r+cOqTHq4KujOJrYJUPrCWCZbKLmNTa5Oktr651BL+q0cgfcf7C8W
oK7SYonOxD3mniAT43+g+PvXopNsAEGe8xezybtUB/dgjznw2G1M/mSKwvGzQko8
JuHfDdh3ZJjP2Fk0vwehrm5iL9XNcgyEgc0AlS0+oN8a7F6qCK9P/hAqe/fgSX8M
c+D8kqR9BSM8bltnUl7X4h4xJc0GTfSlTZPcsjuGCCaE70UXPHGAU5eapGkcQeXH
8lAbukd0IchMgKAWC+ofLZrPIPGWA9Fn6Bqll+xxnZiSY45LwxhQFLCO/zASFGBP
nTwvzIDSbcv+PpsnwZC4Efp807JMtuM5HM9sDQwOIa33vUTl/tRwxMs7ckntNXM8
1H42tmDwuD+hyY06Ny/lS67wm8gbEAL3KaRp4AyhLZWKYIByiE+IU/CJ8yaoHV6g
MvliOoi33VkW6efHk2FqFQlhe5LIaQ/TQj7JvIYKvd+Tn4PkdcbkJ3o8P4ReCa18
BJyky+IlMumVu7t38RkI3UASo4E0CRXyL2ymwyEKZvhbq949XdrBhRa5yzpWkOFy
eC0rZ9QyHJ5QhoPWGc3JsEFzJaAfwOi7mvJ8qE4WFsNY4NbRG3g2U9Q7YPcV4+xV
xfxzvJdLcGOcGHezab67YHCOH2/OoFeqfoPPauK/iT62yEBBJ5Gb3zJy2+Bxgc/k
TIRgd0+jQG7QfdYtIGCzxR1/7SAebom5JQrpttRaizfpmqKU9LT2imhmyPJPZM9e
3XsKGE4pQw1PDDAvg/D82Omf4voTnRCS/H6vrQDTuQg+2xfG++R0b3kKFWxA7nSc
fwDuhdvAeZKeadLVYKqyMziw+JknvDk+NAxV5ksFlBI96SCCQhkuZo0RQvwhS/UX
aXCFEhJgYNKYDcHyuT99tm4BWUkbeqhvA5jHAI2H8XivHYcIMfN8HbEzeqlY/b10
nevp+mYVdNlJAcgYCJ900iaGJ9ozJKJwKiBBOXjujA0ziMhD/snm/1bOL2IYdKDh
Fm4JT2yLdV19j0L+bIMedTyCLYl8VTzvqvYz1up03xXl6HbS1neCY2hy+OFDC3sA
aiRg2jHWdePsVjdFeqY46wMzXYYY5+So2w2SZrIwX7QcDPPCFvY8nlzh+9xFhkce
Mf0zW+3dHKp4YNkw6+jTqeXasz/26YHMfEi1LAIWcKh6C0SBhx/D1NqtH/7sn9WI
rGoFQG6Uf8QJQW0n6qFER820Uw0B2K5KHO3LkSchqAjo+E6l8z+PQo+zYDZ6gEjc
JLueIg2EUNFH1E9vuafArK4FWa5K1EWUbjnFii0TGP28qR4l6QiK8sIuUZsNB9wT
pkISsOoXrZpUocMaIgRgFH5W88HPEjixhGpViuB9jRJkdyqKgfJO1V0n3wB+9R4N
NMQGUrstGwgAluLo/Ze+cIxb0viwGLD1kmQ1YN7I8IHBE8MVKug22YBQbx1sG8fZ
23sBrXCoKNDv77daEqSjRJsiIU78i98qkLH2BaTcdGWpDqgDCwXkTTg3F4z/TDeL
euGGIK28NLLVAtf5se/9O5EdCT92W158uFZWKmBFA/aq40Hry/MftLRZogLdOQZh
ZcCZMU7mJXMp4q+8vmX/XrZOR697Wa0ZuQPkLiXLzl/HlPP+5tKwnxuoSeuUoRmd
RFKgJh8MzatTeHH2eebFzrIL9FAMVrlapN8PepsLc3Ucaq94jBuZ3w51T1RwliIY
uUpJKrgMGB+mV0T4BmQPXKsS9Be9248GGVdGsYwsNCemPNsk/oAKQt3CSR2n2YV6
vN78EPyjFRHitPbJHKpzSi3q3dnK/F8oEhrDFERkp0CrqT9KwW7U/oYLKeVVwrL2
+Gv+PfYw5+2RXtqV74mwrh2JlfuxzotixTnFpSV7OvfNUa6mqh06bzzaxzSAyRu9
W92+EyqGmdh+OMno08ZP170uhqxVGM22ssi0eQ0QZMXmFAqafhULqCCHlPAMIVws
+qx/ODBuLWzrEFHCi7pHspkYT1KzDDT+gNwUIQZKiqlwkzEk1u+U/6uJd9zed2HU
Yc77QuZebsZfvl68lC1leiXBNE7M1bzvQRrTvdcMcCghIpPj72VJHfoKuhcjw9dl
7chpR0EfVI1KLZ6zw8yzhi5KhyKLlgq5fBLxtLfu0ESVnjNaXyqm2wNR3qZV/kHm
LgFtInZ+zDgtdpI5mHXjpNAJtNASzrn1Qyp7bvLzGmuUWv467J4RqP1cub/pkLcj
86Q5V487cHtI/HoOhRkfE9b0fi0da5Ff+inRvDfZZP7djFP3kGNjZ7/O9rwboAPP
9ayM6z37MBIF1hLkqrrUReZVqLMqTiDwdSOL8CHJntkAqx7XaLx4igTCo0MHiZAu
BEJ7/uKW/Y9iiVryAsF2mcxy5aB+W43BcQk9+wJtShSyiA0OTW1bKTOOdnU1wo6W
W+Ia5y8a6nGbH3bREG4ngTYIXpSJgr6glVryZzRCkFizExsq/FNsJL9jJSzT3DsS
0hRjJyo1VlFvs0EjF/5GoSs75Ir3mnqFpOp2ybnHIFw3uU/VLnLLve4+NOWCYaR4
Mama25bZAKSONwOebqAzpT7fD0ECiCLOgE3EQIaI3o6i9KVEGcLf+j3tbs+JrvFA
f5VqxkG9C1vr2K+TKHG9wRRAGDiDWKlvdm5qEocaTjWxu1klHo/5yCIZulIuFdlr
vg4NLPnW7k1Jrk4Q97kpy4yC5iAIxEptA5Ha3R0MTUcG0psgUXPcLaEnXe6hlBjS
TZp7lcHIskvxigF+mAwLOEDAJsJqLUEtwinyO/nnG8Agl/deFHkSoXOP1vvHIBOT
Lo1OnKJN59jOycl+dTCwrg6BO/RO2MhrWqswlLuGBMzB6UJV7ahArzuwJzEt9jy4
UN7mfzEkgmQapgherveZ5QCEQzEBKszkgw3Qy3T09Zycj6QVUSMdDD9SyTLEXpgu
6d7wRm8KvowloA6AcKNP3fTOeM/MRjXaiFL5exxWDaj+ZP35W2MdSD99IoUomqO2
erpz5wdUYDP0cZ6OqazEW4P+juaDWofw/2KhAxnAdvmnVR6FRnwWKjwpJd7sf1PC
+1b0agzhBWDgDMtXeK4qQnigMVFSJ0o5d7zGrpFZ1dTCQ6G5VH8PpJpVQ6C19Flc
WiQt7lkWUr3ToLAFYyuipwWL1k8RtMf0O6vB8bi4WGFeA5dKXwCLO2M4KhW3J9YS
I5boTdDEFgHeJ+kQQfDzakWXXTt6Hg4OIatwAaBgFY1X8dKGEpeQFOBqb4NLCM3/
bhO8qgEIIsEnf9oeQPWW3Z/fKoAoYhj1crD2fibSRfYD0jkI70rMdubuIFlk6Zux
VTeXqWnoOmZnBmSgELRMsyPvMMPK5V9Mc6x4TQ9Jtn/Ms0AqwMZSiUKe0o6E5rPh
4nnWQvBubSoPaYdnL+2HPyqGdXASyDks2/Svw5HZXoskFgjkepJCCcPH9lsdDccf
sJl+qyphF+9jHUfX60mNZtTrLuDjXsoPTlLGnlN68Aw1+9m2LCxRRv2pdNNvYNP1
dqjqHqmdqZde6tZKxMBnZ/ycFl6J/Wl5t7yvmu6aOLY9C79KGv5Tv3rG4aM83dbQ
USD6Z/ZGujhaqyEiqJu1sqOP7PWKpgSZcg43JR4q47M25tY4bjs03prwDCLv3qxf
VFMaHOiaLYF8dkzs0/i8bnAsszXU3mcdALgeBwlDVpSIqVOBv4t+NVKm3mKRv5ET
6Hk3BPBb3zvkX/b+5RDW0bYcq0vMIADG+pKtWECqXLtFsfPf/EAYN1HPPacMhr1z
rL4FiSpJMXCL6gN2GuOBgYADoa/E0CCC2rAJ/FP0Dmn3Y4C2tnV15D8abTDBI2Hd
jUWEV1KbM9PlKAQXQ50dqUrOwapQlJAhL6R2n90c0dpXNGA801gYpoUl30n7rbRn
91lDoUrblt8Fpl+zhM/sp92za6ga7XM4rxKHtBjUc8QpEpgCq6npChZYtJmRQMxK
OxeY0WYst0oZmTUZIQvygQbRp9lAiN+7LTBR3r0Q2JqktOh2EoCnMXv4iYtIaArB
jFnlGLnAdEUgtE3gNw9zN4VGDlrE8Ogu3Ie2bzpCIEVRwWYR3ss7EL33qsh2tmLL
BiOdSWjAkQa+Bmd9gnKHzjaaQJBonei+eudImCyIrqHw28/yjy3mb1DikCrEvPUh
NhSFmRtK2IBrX3uAGZQ5HEHBnjzQqoAmqKGT5soWSulPv9HY02xmzr8rv3ArcV1K
h9I8p1gWJBgOkfAIMLogrCmBFV7cSbjnqCaRRFDH5p9TUp/0i0DDTlwiJYxLRCsb
OMmjS4O6gMAmXMTPGl+XIU3qle7Z+BOxyRYjI6oc7cQZmzVA0BIHNEaVgczjxJNs
GIDJGeN9AaPKUgq33SIwaikjqzK4DPo8pzrvwUwQW390NB76T9WfKvvbQemTdBD8
moAx5qGADleGzEeJ8FG5lZ/Srg18X6x0mwYqMRJfkOmkbUEO9boF2RO60/2Adai5
Bollm2G3clq8QZ1dBhfSMFsN6zpGa7hKtPFclDEI06DSgSqwLMn8FSb6gZZjb6up
4ljJzqe9aLhol61kFvEUKoO7Vhi9DH+poO+RYxvkactxKbXg48MRNHkd+jxUE9T8
Ui9cC9xoaDf4mKAOp4X6OpSpxy5w7WOuXRiYVemQ+X5NI8zOzeOWV2koik5WAe5G
679c6cB28JDHVGl6YkDTfZGZYcsDtH/6CCXoIq3jQYrixMOq8AvsCWHqRjjOOW5X
ZfYx65MqfMwmCxz4r1KU+r69wT/2OhOwS/WLsNH3Dg/D+z3juzAfX16S+/8t6FzS
5Ks4gMJBWKo5abeOdUrJFmODSSValapduFV3ER5GJmK8OYIE8q5V9A9xVfoz7GCQ
TnDQy4RuCKSL99K0Umb3TYOZofymS4G73dCBlhf6ijNUS8a98x/6YCRFaOIsUOLI
/TiVv/+gIpSVqOuYw8eItJHX8slkkSFhE9hsLFprrpC1E4TWKDuG1rZGmjea6l8C
HimhgxCkjAe5fdHqjvQ9ik7C9ETzCDjxf8r8iekXEJTc44V2NU/SrbkE5rvaNSOz
XtKRVFGyCzuxWkZe3PWqXcCsvbAzlSBesEMzqwlU39fXPi46/Ka3BNFxmjNwAhOe
Fb/D6oYNsJMDEVGX5EblFBO74ROr8AnkhNohPKhLXnjNlxnAzHs/vqieWvm7VexN
7/CVsVXbdKcnUN1bgSH1EVOBX+vtt1uoKurDyAoGJO/TMXy70C3Y146Pr83Bmws1
QH5XU9RcnA/pVrINJM+0VFAVxe4OVIicjwkQJvaiVMDVis4eQuuyYrVZfMKXGu5j
H9OdFaNwKXbrBVTLKXhoOFhd2rmqVIAIpPzavVYucjDTrMYMSzxZALhYY+OGtdji
b6KyykHZPcuoibNvJ1C+ly44OuDu6pMi4AIgKzD2rwAKJ/ztb+WnRm3ykjkhghzZ
d/bVagP63BYIQMASy90tjBWaHqx76lBtbDQvEP8SsvCjYoT2mSxBz3QD6BQAHVKe
YDIwW03J/bdpDBLUv22YGi0lb/Ryf7S4eBcDsdQ8cg0yREy0iIlVe3VyrMdEoQuE
VWaUD2+lY+1L8AMd3I6bvaDmjvf8dMvbSPU8/Imy9tajdhnC48IjmJzxIh0k4PqX
6N51f1XtJzbxkPNoWwKEKB0yJEUqC5PkT2GeY4r7MMbPn5AQUAoQlWKM3nPRqqTx
tp5hW/t5yNEBuEUBl56tgxu3HcwctJ+fqcrtTPQecmJNRMdwYjnkN6JBokdXL1dT
bHq3hm9VZPeVthMfJmJhdp5hESaRHyrqEqE/lna/z24yUGT6uH2paqjAnxlym06K
GaBEkb43upnUvQopCwEL6bpp3/NYzcfmYiRbYrDmZTwXzNl8ZVAssj3sH+yySz33
Mv1e7l/rtZBfVIgwz3Y7zUALRUT7OyCbCKpOWQJQilyRoip2K+6o0r00oZEDVFny
6vXG1LYwdSckaUbdXCBALBYOQXVTqajisGiKsd0jZA44u541eDlOXZakVZFoQhzY
l/IVSwNGm/LvfT9Re7k2GdW00GHrCieSUqp6NBUG9FwPhZbclltTHyJMGr4QKiQV
9p9Zvd7SnctKHP4C+CpBk3HdUXcphIfbLRLWU1lM/JAXr/0zGbvBRROtmZ8NU+0j
n1WYQl52XVK5dNin9116+MArWkkQFCfkgWBtvsOCQgqO4uOFWHAPIsGFWfdZoo5k
IPl9lNZcHp5aKl3XAm1b1sJKWlsordw1gfII7wK42GHnBc+cLnXNqa+OmrhKtbt6
ASkpAPvpWvquGmmfVNi8Jgq2f6OoBuWxd43MOfjtsxOdFPQkRw+Lsh00N+NkctZB
Tzi4SedhBQXx9t5iJqyXw6U0YDTepMFKwnFWZeGLY1K2vZr3Nqu+tvNRHaV5U/Qs
9tTCj2Nfvwf/m1oiRNm48kVBec/mhS8aZTuRKUtcghDsuG1qn5aNYura6ygMzOWJ
AayXJ7ViMzKFCNuPftXNd4TApLFDPAiwFnp6i+X7hGlODifUUt1WltXocfNe+JFA
evc3PJhALujlMSF3GapolcgARWZWHQ5Fok2aH4qPJGjEIOMcYHJ618hKBdwEGL7K
m6Qr7L2a6lRhi+QHoaaBB27UlRR0Pg/z9rP9yekmoaTm+c6X8HIEFc5Qjo9sDl1i
lphGBucLUr69btycwfDhNxp092zd4CClvDQNl/JcE7WbuSQA0/ou6+9Ucv9xbO7q
surDfJ7cpMZgRcX/P5EZ5SSu2x6YEINicEHn23CPBWRlnmFOnue4ADr0/dXItEVG
OSyWYA706FRieDBQq+PukeKfeExW8zxwKvBW3pJZHURxLVT0CxdfZJ1Czk+2ZxbK
3YXtfG5P4gjvQsiEaIMvhCCF1OmTfLjiEmGUOCPBSpeoO3OTLo3YibgCQKNrIA59
Ih2gcoKudPcuPwa9AMmuHushgYBkbYOT6YBh0eW4N7/wHnTGN4He3IuadivmzU7d
Hkowd3KsCp/gvnS7p+EWQT99TplIirJPHfrINvUTwifvVdl6PnOT1Joo7RM636uz
uzw2Hz8pnP4YxSPMlLIQwTOy+vov7uW+npWZPr3BOfQs9zUL6QudV8vdUt+6bT4p
QUQykb8LU3ym1ZOJbcq9uHimt6M/7WnpjCapig6kBltQjE0Y68UcoX14BKh49Zf+
TORqeUzYvOqHhdrMKuEFfZyWUmkZXTl5ucq+Z2Cp+agOVTXh1ZsoB8MHtQbAiHZP
b/yNDYrRKvHSsEALZo6TfDTTn/4VHT8EvncZU+6tg6B/E6WxGvF5GeD/YElzOVNn
Ku4r+VZrJZMl5gIi/8uc+kbZpEUe0ozUjFjtOA9mhaVkYSVO4y0P2TPlhHYnAR5g
Gwvtqo5Q+74U7zRPckIbPnVi1PGBh+AHKLxSau8dCyRGjv+mVB4Sxl4Td/cJpEQi
B1zMPTc7RUuPkOFPoMVswOzKZxNsgva/wml4oe//xTn4BwqNzW+7APPXXyBrV38M
uqdpAQGT61zk1nv8B6Q4C5a8LK9V2v1znRdtptHdzpqHFRZn+SMMRTBcnNQIWap/
eoU4U3qpHy+TACPKwAqrddjP049naH1n7pJb1KBfpBax9XStRZZ107nlulyHSR+m
Nv55dWofK5m4G2Xzhs2D61/cIaSIsSIaVwkCTtTEvdqXHYQHs6QeCWFT82aJd4jm
Bi0/iZPoJh+9usZbAcYfynNFkcgbkYQC4qLmYGSDBmRdrGNb121OnhFeVIbEX+uF
Gxr0reNwDL/05clCJM3Pr4vKmDCkzuxtY7gjZB4y2oo/mGU1FZOR0NsUOaaVSvFF
btltNHkI6t8u5e2ZlbhbONuVfEdGBkR4E9aLKhZ/jaX5Zn5SZzQ/7YRLyOPa0JM4
dxSOxJ+M7qbSp7lEinEAwssStlV/j0McNST4o81IAEMnqXPE/+1ay9mvM/oDrnow
+xEL5BgPZEmOhW7HhWV5zZHh0ljMqEYI5L1sONZBZWkuBZTgvsXv4tpAecIGz+CC
EqJhTnStrnu7cj/9dDLd/PcAzFQQ1m2X7Q4DOtll1VFDE08cPklEIS3djm76kRAO
C0gHLc9VMSgbo8i+fIezb0RCxFvzbi4QJI4EeO8L4xxurDc4glh3B6VvkLCaiAS4
qBhkQUWczq4RBa1y48pscUQjlvC4ajgxd/6/5cKC4G4FEv0ATDd8cj9CXovjXpCr
IynPnweJ3eb6jIq0Q2j8INR5HoXS6HYrDhkvrbehMwuNVMjxezWmFWTEj71QoEFn
3q3qPy0GqRGSVzJq1zNCGnlAATR3R4S6oZdppv7SO7k7rLOBaazyTMr9/hf11C/o
4feK4wWzS+eprmN2X7Hu8GjeTFxmoJjYuN/z7YqCAXvf0FaMUzqhISi0wosZHiFR
NbGW+eyTQngYs0iFOVnn0YH4Wx17vqnYgScwPYrz49fWP1jrg2yWW6b15Y98/skw
53TsyXAcxZcrXaaQ1EkiVq8QD1tuNa0tjc54SB089jKKVRbDqe4BizCI/uAfprv9
falLjdbc9b1gdCwdQ3tVbJbS52oIwgdvZacyxMup62vpdq68HMaEIb4PiDasakCR
qi+OMpyc2chASaeLLbbt8w5ShRK/STQrwqgr3DXgbG/un1AJUdeOHmYmtV9PMY87
D4G4hY+ylhCd0XvnUJidUdQjUPM+v+mAEPr5/5umxSkwcJJfVq1jEzE/cV8s7k1y
1Le9ZZlcLs7Ak4wkIOs3Bpc5Ff91eF61emdEYgBGJmuJcehJVQ7yBgwOBslRxi2N
JBLn+q61vHVwAUeBPVAyMCqNXAOd2I5jXCEg6BiUY45RjJ2llIgkuUiI7NCl9G1J
G/yYn9RXXjQHllPIwgPh0zLYcD/FA62WgRKDx5N4ZJyVwsoQKw2n+9oxyDVDWIv9
rL+YJz4yOy/wMsX+p503NEsKTwHdJiQtNKXIcGGvvKHB0siPPq6SGXnWTQ0askzZ
Y6mbhEDTSceNsNnCg5emXTIzkTYPcsww3i9j+aHEbgsJKYvqPJRV3VaYSrKM9TQW
lBBE/yAYw5smoyhuh0hyCFyxEgF2khhwkEc7bmI5gtBvfVvX1E/rMVO/n+gWtsJ/
+KYadb4UFro4xDP0C630DhVtDpmzH/Qxl/pC7SIFW0IUoJZUVdawkgTyM7YHEnKt
6soPPjtcDBlI7PkWcK4MkwWAPBc2eApTBtH/AA6j+mxJJDZ+rjd31gYvLFuXYYlJ
VIgGLjSnCxTqVLqRJGG9OZ2NZ6QQIPUaC5qNGEGjcLN2j/VfqiAvlVkiKyfeXHBh
cpKXqza5O8Uocl5DM0VyHsQ9XEqzrKxvwyV+GcaDyrDSkTTYBe+jqeDYBgxJXtlV
BVv7MbaLUS0Fh0gfbrYlTL/MbPyfYCZmytpOi0H3oXe/SrLQIqDrq4W5Wvms7TZZ
pWAkwekhDpq9l4W8MYK8KD+n2Eb3PLwZIS17P048nMqFOJIQS396o0RuBOLxWDiO
Dgr4XuuqtoT9NemEaQUvcFWn6v0+fF5P360ha4SNb55vvmbCARD6Y5ITdUI22kF1
JatkKDdMEAMS8Qk7CIdztoqqr4AW96TjtvZmCxHlkzFqBEpIQ9lk1fh9KcQKZNVV
6k/H3/oQAOpKF73NvJT1PD3ZCZmOrqIP7qbad2vWU4zrZwWDy6KgwNyPb/ApOsDt
jSdg/DdQ3GXHNltiyx58tbuetqg5tTGTg8zmokH40DM+tfhnYeAkqhO0BPsb7tjW
QRtDD5HChtUFPQmDsmjWmh2Obg71qJ/gcPhFGe7aMzq4jPi+DlU8FNwN6zJ9+Ewu
8uZA92lOzFPd8vQgxTNzDE3LfpZDzomU8rzUm0Db98sysTI33SK8zsK917Yi27Y+
wTaYEdypu9xWXMCwItyodKj/Wdui+rsJF6gja8hchtxUjL74ahqt+9vMsi9z/s9J
90pS6aSloIdcdgDezDLnJYbFFUMXMvOhCuNidU58GVS/e9i4+hSSq7bEt3gUx/7U
1l8qkjGAtLV6jMzIMx7d7YkkvvkBQ4q7wRUCg5F6AGziW98LLgJpjVSCHjj5ajv1
KOrCJpiRHN3tnQhoykFxztGSwTVw0/RlsrvY2qnJlBy3uYDE+HGIBgRqy4rp7pHe
gxKqwk/DK4AMs6t7Kc8HFN2cTk8fU8I9J0b/mAAtshGlMXZmk2HGDF6X1Pa+XXJK
AAnqQjYz7BCA1Juf2QeQL8s/Eu0f0bDY7ZUIYAaUfBoPTMJmMfbD7u27HN3MOTGS
VaZcaVlejtOi1oyHRMLUnEt4YF84lgTFT3UN9HrdCrxRd27drkFeK0dPcegAG69v
qzccCaryp6BD95c4aX8cGSyJZkPuGxzobOVBSsGETJndq9vJ6SbmQ/tI6H/+uhsB
fZAmJV0wYFbm9OjYigss4pkxW+NEq5p5NTfTVAgyyq1xOr5Md+7ByJx61RRwh+kK
9v++Ygs30q3X7RkpC3LXGg3q1pxJQmq96PZGUvEbnt1zf1PPsIuZ/LMN1bOWAJ1k
1/yjfGMkcd0u9OUacuyKGh7RXdde/4f4tqX5MiEkRKDFb8Dc9GQHPmCF/3QkX5dU
1iewyIKcQ6fuEsXhKO635AQ7rH/BHVekmmib6ISNwlqgCcSjYQsq+NGf12xcwnZg
d6199xYueaUUxGhSE9AWFxMkAolPgKkDNhkXX0DYGKjDrJlZkD6qon5kxXDnhkFR
mVFdWqEGMdQQMeSN1OhmuV+FzSxH932bJGC80Ket70Yf9FtCxlKaTQe2PHpj0BtN
IEKk8MWv08U70h8hh2OVkmBuNtNheNTnMkmK0AT0Rr4aW7fUcHcrb46M1UHEHcF+
szolYSQFt19FlSxaFWnwy7GhVoEOYH8gy1MWrG5eo1QX/+8Em+m/V+B+8nPrIsED
/hYf1Yz9/X0ZTmDGQ+mp4CEoVH2aanN1aCjYca5XeIlhfKYrORPSFZ3W4bJvcPma
yFpM8jsKEkaX5RG6PnMOCKxOikt2g2+gryN39jz/OADXL4V6ta8f17CTBz3mQBK5
rAk0TETXJv2kYZP7F1tc8JHsDWQHIxKQtwejpEpJ/sJkzfoULruoOsL5FOCaNsDB
5piFsiCbQW2cMKDohbCpR8oI+FoM9VSGp8qAA2i44o+/0i1V/caxxnSOC1QC+Mb+
PHkAgJwqUhWDaQHEEqLzYXSP3fsqC1L/Fhi+L3OcguGRe7RV+/bFIw9aulBjH9J5
yVmDKaPDKTYwb9wK9XfWoyf17r09XFbVYPpxIPh8QMzxFYm/UjGPSJxULwRd8ThY
w+s3jyIo7/F4M++Q5LbnDJgvwsYauvoHcWZDYjIugG/T8PBqw7mO1sxoRt2wvrIg
9YFlrptuybO+wC8fzMxMvd1eWWl6AyyDXgyPVx2ovuO+sqlnQwdSfvx0p8MuEYpc
I/LFcp5f70iPuOVHreWqR3eUTrtTV6mK1eGeGyndeljogo/HPcUGP68sY8MB+QTY
2bu1JBGoZtvwjfvknZXZsNFWlfNXukBUacjuMlCGkpE6H6nb2iUmHCxW1R0PrLLw
6hLyNvwHJpzrZ5r+GtD4udCGNj4cx/HqgBgUUS38jkdDmJY4g55Lk9+sXxjmSfbq
uC1wu0GzqmJD6bnqGyGFaU2WlQds/uQz7WL2dUKracDekm303VsIsrgzlqQlS/If
tLhIEHb443oWzBocfDFrVMWdGO809814F5qspXsOcBhSVzr46Suqx27+DCVYpm2k
LhVOZhw4nbnj98zBrNE8AlZtHxTPmlMDRAH6ky7woq/HJcAE8lsowJB+xp65iHM7
pjRMWM5UkAwNDXazY49TmLFjGG5cIOPzcuCUNhXahndQr57ckVkreVJpb3PHsidk
vVxc4I4OGQ4+0vg12kFoDJJuTGaGe68hCGwBWi2mYRIRh4QYi8ypaTJYqApN3wzV
i8s1PIbpkBmnuwZYLXZ6gBe6Hy/6rxAxkGG1K/jBqpIocpSxo9u3/S1q99C7q5FY
CYezSjJ3bA2U5F1GPogKvUpe0vqLcqY7AhL2CpybVoor0M5fVAcyHcY1qf5eo3k5
yBLos1XmaSXzHTzkOg/CRQK274U+sYxQ53YYo+vL7YyLMeetyQe6hui3ArHePOUt
LaICzTlwAs1mnBZaV2E/p7o1ygtvKd/c9ydgoH064KJ3enXVFxqDMecrXacz3pCA
/Lpj8XLbML9ftGQYkPQUWGiumt7iuWPJO1x3/JdsZUAQRlwHdra/2laDXIMirfVT
JYFsNS4NPtaif2p05xvlHOgm0lH10zfgdWY2go72CC6SfMR3HneaQCKegqGQCzy0
J1oi8vBKJWh8yOgoYOyV4ckK2tW0++AGSXQR3S4fmjDZNXcRBhJ8ZjeCgfxLYKRT
vcK8A2EXbgsDDldICP/4n036epHi4RVTMf/5Sd2NA+34OjxzBYds/r0cxDgpAXLE
/LhPrQ1hum0MZWkQVhsMfvd9ufRUjv/692db1cZgfomPkkrn2dd7cbTt5pjaf43/
52IXlv+p9msHMSLTJkICkHA4Idg35YpkBpFSMc7ZW0pa2rvLVlZxCXqFWUimwhn4
2tcHpNiFul1mqTBasq56OUhKpU43Jn5w7NNGIdCcHDcEpSAm/kvrPD+LgIfcGl23
ZROKFdydPEXuT4cudwUS9Pc2cOvZoruXqx+l2hAXSZBqMbmIHGTjkHSjwjAIKkcE
l/+/sT9l5AfO5wzFD0kdqUt+arUEDSwvMmkjk0SRtsk1xWDcckioHC05CaZuIIjf
JeluiW6hlM95b63U5cmZlxhk5ULjjBLoQKb/dxyXCnKixjcCe2hLlMXVPLvIa5rp
FgtUA+KZxIPrEkcZw7TYWKkqa7xTg4z8ahZc7++HogudCA4auC+A4wU+mB5jfhCr
mFm4bpJfTLF+CsONBuAyouG/YBnUl4NQemckP6ij7Y3m12Gc2KXinJWM4e+PZfEY
0anYbM17yoCyZEcIdexXfyUcbnk3IEv22AE6aPognuBp+fsCNaqTTht2Zfgtck0P
qAfXzwLBUc+a5c2XfFdch1ICh0ps/DBm+5TDIdoIfgPVO/uy3MdOSeh19QXpMqnV
Z5Q0+G0GH4XbCbsaZcUkdAuxQLaWk3XuSgabEWrsVeNVWGTNSbTuSKsthDrcyiyt
KaQH1IbzeaFPzFm1LLzAXXch5yRSilldJg5zR1NbUJKh36SziNwWecHoZYWi/W95
QhgOUNbkepEbvOeyfQCCgNxkzB/Dyq8vKV9KF3keLAQ3wo7CqW/sp2SE1tIuutdU
VBX7ADfouBo/7aFWclRQ62uVdCkGS15ixwgT1pBX/979XnncEavie77Q4x7vCKbE
DAZZ1I3hYiniQAVe0JMXKIQp3ocZrsN1Oyli8FQYiTJInqo4WXHVuI3tW7hB1E6u
UodFr6n+WzqC/e4s3b/GJr64mzc8/KED2QLSUAi0zyycDRi5MwPmqgRljs26iIBO
KyZkPEylruGB9g0oIB+5FJrzMGSP9KapGQN5uIe79LA2XDpBkV7IQhmm/J8ovX8K
Yi83fKXwtC8llFzZdCt+F1BUBeyFFaEtByPkutSqLDV78z4ep4B116+PbWl3oImU
gaBBEDIhdbmdAXanXNJJoTa4mdZ4YCt1dwkx4HDhOuC3be4W7Hn3qRq23Eh2xvLq
UNyC/+pYKxRM2IXGFoKXcvyKmWbgqylcjvqOnFVEjdofkWfw7caXj2PzxgX/Inu4
zycAyVb78JdTJc5+jKAHlHNNEQ9K/5GZzBGCpq7U/EEDPogb98jvr9lhKACzhQ/0
hl29KruBOE2dSCKEodJ/wsrM6+axP/ez5cCLWhAXSNRWN+9y3trnGc4gSax8zBXz
/wFWP/anRBtrglpzHQHNMhUngfghq+9Q/shFGmqHxR3ZjGq01CctdGhDmHjejk2/
l40nccf+1y+4dSQ+KVUs9EdMTG1Bzty0cw/wsxpyphQg7jBV88hwwjb1vlP1/O7d
YdJEBij67FzgqYmL3nvoehYUL4P8pN1CVHtfbvUQNjOK5xothl/XLSmesmLjS3/c
B8jdo+D5/xALjrcrf46coqnXe/edH/+tKZtHUmPAwtx9Z1huPN32/VOXEtQwhvMe
lXfhrY9jQJUNL+LxjeuWbZVD2dlmBXhK7fWQH9+5rxRV+VP1OW8/f8WlwcDSfiUR
8KHaxxI2jI+/ZXKyF/ON6c61kStNNufRUUH72sLQEugNXpdLGwUS9a8PLbBUf/IA
fByBoksy+GShL3GNPdRZ0wHOkU0M3cT6jx8F5kLFvxeEZhfaJ8iTk5OSdrUTyRsJ
Ata3ZIyy5SqnpGldZigNFSLdolHOfpr+4D+lDbYPxuVKwQZlGP10Wtq1uQIvw+ma
ASB6Qy/wcARTgIk1EiHB6PENcp/W5NjdlqYrsPJFh7BNsPiDParb4+gfNybAcg+6
AfDAd/9TrkJ6KVRuVGOL4Dy6FHh9fd4EmHLw3Mol7b4l1ZkM15PjBa7AAdZEuOTN
pL2nyL1EORTF2rXTS8V5u0uIwb8TiiLKicrXSlDOE2V+CPgbKRTh63p6tDjlkbUM
NZa1cg+MTlYAhvcLnO83HsahaEo45cAcw8hMwGpdy0kEQ6Kn6UO4Xfv5q8VDDrIM
6nqSrRYyG8wIinZaatpas6WIgOzV0cSzC9cZtUb0OlO6CCijXIlE+imulGeBHsi2
kSjaYUedJ9zmBQSglhFHR9oZyiNBILHufQB4QinP7eCbuR5Smossvgps5ANucA6n
3dMqJ7kVrWbIRy+22hH0uUWo4yJtmznbjGyxIXc8DB9hL4t5Ft/eyX1kLZ4CXi4K
CmzULxPJ/Lcmy65OvAcKptkhAnb6KWCA3kt6fI+w81yvy2wmPhFlOzPdmedfgN7V
p0fYiJc3KoSPIGp+R9VY0+0hS+ZMsohXTmhcon4LGBffKQki5A1Ul8PhZh1MjleJ
`pragma protect end_protected
