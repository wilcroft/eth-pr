// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:14 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lpbD/NCnM8rpkP1/8pNI3kSOG99tWPnPrbkuAhZDjGIeL01tLiMMhsKzZYbOF6Q1
UiXwZoDhe/QdcLjBA7K9KWrScpe9mzvhp7MVhBMme3ceH4TDLj3qNM05MhH+gNv4
lVJmn4+lTsJV1HE51HCq1+zjcO3Z1xttAwNbCrmYxv0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28784)
1nHhVVhLtRegpJ+aPqhuXM4q1A3iZpL+HZEYMFtGJtgqO9UmZnt7HljkqyUiCs9M
z5zR4ZcNoJGsT1DXrgnlOOhersjIJ/5E2ooaTtuyYiuhM79LvUEwx2FOTVE2rM7f
ybp8xrfmqmL5TwdJaN2UZXF/9mAx8TzPxjyDST9FW2o8HlUDWt6jpbOPgkOUMtUB
wtMAziWTa+BWkYDegkh6zZDzdyMxvfdJMT2qSe9/+WqJh0CCMOOrtKvWhWjvd60G
7j1vMNud+UWCJyZhZ6+NHxjEz+IiPSxvPNv84jdWR7U7ClL4tupWDMvl/QroigwV
wdK2hEF11NsvHJyq6s07eCTc/mScSFPuf2ZyPMH+JurSUTXaQpzy8urbyZFtGJDd
9nZ9Ur6Mbi8y5vIBlOCkeTiELsTS7IOOcvzF/WQmquVDQsStn97tkJ2a6d6PAYkU
Tnw4RDt2YwIjP/4WKmyDoCJJ3TsKgajhcOSfma2kIyazdXvzkjzqbsMv/IwByxAa
0tF4UjZOQuzkWJWE8ibaBhMQ9NhsCsRuYKAK3MJ+oY//zsz29q4e9SrtXWRww8j3
gfUajYJIbf9S4WP92PlL4N5sZi6SEJuQcWXLEOM4ZA3Roq4RAv4BhHprXv8n/GgU
HNzlfIU00pa/qLCFwshKBHDWv5fjodl5hCVMXBu7FzTbo9fYB3kkGF462DPprMZU
JxVXr7Um9Jj0NAdlW3+mwdQ5MgZQseq2I9YYAwlg2RcMrkFakKiFBhoUYB7IZYq/
sfArfnGlMfRibskdhzZBox6K3XDw71r5S8I9hEkTzPWMPodfa/bV3C9Vn4rDlz1Y
yFfB0bibkvUzzJ2N936QQUaL9Vqp4Y7usihH+Bcag4vQdfnK+XwFbvdEZIfaZpgA
90uxfF9+i84nVs8a26ag4Y1LjFNsYMO0dqZBzh7IQ8cHpUW660sndVFgcHFAxQrI
nokhgJGpyPVPRhBRcbjBelN80PoZL4o5I71wcNScHGuEsXnT8ShWW4CDCZbChrB7
yC23JqWn8baIzqa3iXQ48Q25WYierZOnVMgzZiLScGohkFkCOHbnT6KUuV/ue4yJ
T+qaBGhcHC0xNcajtRiCpsejOGuwPqrGWcVpIn47IJ8lv7BAm0io5FBoxuWB4hPs
NB6DmlUUsbyJvhY6DJipQRzl63YqvKpiej/CdKFjt5Rv9M+pri4eZPvfU/BQ+Tlx
CJ+jvuW28zs9UmaVm67w24agIEMLgb5KsU3ajdwr9bjiIrBWCVpGB1sFPswRgHYn
xm1cyNdvkmNn10wI8ZVIDqObQs1RPyh7lvbzw/3ztv3/tCShFXWdRRAFUwJWDonm
OoIttzJykhWyVSNq69g1m0L4atBjKIHBz4Qmtu88po8yilRXoTwhckP/IfaNI+5B
wMEqCbCMT8Cc5rM/KD/IurIh9Fyw9BFgaHedoUMu8wUuIVw70XHiUxbC2Us6giec
HqstXH4fHNcck2EBmRzFa7Pkh5wU1gcw4N63vlprm7n9AVjJegmiE20/cuTAj2op
PS/ewMoWfiEhh/KUKvzW2Wa2n/u5JmjyX+t0gAeU2Fm4vOEGJNmA6ke61tDigIhE
9e3XAEOP5tqjoeqMu/PBpsy0vKavhyajuhCmsBBjeeXX08qvgjIoCCG3kY5FFuHt
tdtK8WOpZd/1HuCuVUZ8gDzX9nt7S4YX8PkkN2sk7IBlcK2X+Amg/CuMbyd07spQ
p1vesGqxZsEaLXoEqTPSPpB834NgLzCcgFnMnVnAtwpI8euRXJBbiPvTyvBNSNio
DgIk7bVr1CpWKRuCiXgGGxzf+ADWwHOY4DXoKfsjB3OatTqwhRHvgnnDw74P5exT
Bpzfx0jdCz+zAlWhFX7h/fflneOGLLX22m7qs1JftRmFuA+slFWEn2kh9NC9hojH
896nQHu7Sukf1ssEKGMFjLILTd1O819Eh8xlTfGdk1Q8n5pPlAiu8I0G+6hqlzSj
EfntTaUTkCBxAf8Ppyl7cRZ+RX3X5XwFCzn2NKAatMrP2jCiFEDMI0iDfoeGDlYX
mWI5n8hvIS9KLVHEEBbKdevjjHwGGBekMQbM4r4/RW3pUU4k2yxbfC0f8mWchuCP
T/zVypXThohzUyY6iCt0idgMOHgHKJzS/dRrELQKVOyjSGX0pd9zfJeWuDpwHpMO
FqDUWkTlqFvKKLdYvQL+K/ajrJ8Xm5zqncKrhZlMER79KCjjpRHC0SB9IOWe/Q/E
yQrxy53LDjYSsH5HV6G0cKbGRZr7D6+ZEaFn9tfJSvWaQNZKh+Wj7ACJnTfFulUp
T8/AMYNd8RzPkqOZzYv9brEhtMctM3QbLnlPpX1jB6fpZPrs2HDeXehSBTlnWh34
KzbAXYU/brtPfQ3y/c9FvPdaBw7MvtYtqn88tUb9NOh/pYq3WLKDjeLKZsU8YoGe
e13jWBvSyvgBlrivzjORheCDdT+aL7+/OrtXjJtanlIuo+kR/FVB8bxFMHGGEHhC
o5+2OtZjTTQKN5zrg18XNM+JvM9ZL2MfX40/BdCN9+0G27ZbpE15k31NBB/qOcrs
bXfe5QZRnxBv6rSVKQaj6D/Pe/9cyqyXicJ1J1IoZadAhSt8MUGpi9Q7O4MpZ+Bk
kMopVwYxjbYqHLKR1m665PUjb+O1yn6mTsZePvUidWVoREyXFwjfglB3T5oH1khq
rrQ8pNMsRq7XIjnr9ZWqwzGib8hRs6viMxZSNZ7bh2kQWQC15U3t8Q8YbAT2Yvbp
EsdGaVw64Rwo6Lwtaw3nL1lcgtXi81ROzg1ibczfCQBti4ZX90HEv8kednOvOl87
0LDKVDPEPQAEu7vHaEsU0pv0A93VYDvZHpSHquSuYgL4+COsfs4CmDUkraongXq5
/DG5XClR1JWyOa/LLmS1+YD1CfG1EZpUDvMjjh5RuIkeAgSMZwyGP5XrZ7Ckql2/
2756PbMH32stFBNvbiAxA5BfqWqLJS38CAx8ia+6uvVyEyqLJsRqO2Zy3ujxIFls
iARzEsyHfVAcQy+PRK3XTM1knV1Fq08NUPKlEYBN0jlXQBi7K0508OQAnu1IebyH
LNozQHGmUCDP1P9yYrmjHdXcshFqIlHMXaou6GAD0N8SbYm9Dsv5NTf2Zjhx71Gy
3TS6Ggwte+rmxN7q9jFSZGB1vTiaZyk6zYcAl26pOvZgcTZCPb5/mGU/aKxV1lDt
PXiDDUWNpiGXe5tdGk9uhP5CzIVw5hZw6FgncHflu4EvOOsNmo0RhgQyJsMPCk/p
bodR+Jo8MJKHZ1oKGXx+kbQvgGasd9feZGAXaHJ/5rg6u8jMgVwpAlDWAL+wLMpH
xer02779zAwVPPGoLSK39mw0vR25KTMTCw4UiBMr899/xf7je2hIzFMQoHMn35Qn
qV0AbclwQ11vKh//PqVjYC3pJSXWox+wbDVpYeU6N+5CZW0bCpnzS4y81eHdK6eA
RNeYbP6oRGfd8EgJDwb2DT8YKgu/Ij0RmtXQX+zoX22A0IPYOV45X2G1sSQEe806
p6IM9SUgGal3dL4gZUGV92ryHo+C17WC0kN/xzSq+e2TxExQo2PuO+wqMl562EgM
3IvBwuXOjz+/4zSvez7jXylBX++HaIqONfj4leBuEt6jiUn/fAqYSQGkLWOy/hz0
qksRnZGe0mVYrt++6GigSg/RUh5CV+j4Fot27oJjxMxYVG/Ix/w3Km7Dh9rvRUpc
izXhc8enqpdF1wSYdkQTatpLZnkMLxGbQp+tGo8rkCCOW5QANX+hUxjet/ZTrw9h
b4oLvh0jg65PyUByYm7GsVigTfUE3ulkxaKam2b61FPvbP6SxxadWeuHsp8lS/nX
DhaBc908nQI/A2+30ncVFxPTi6csdh3we9NCeLYp52nJ2yXkY7Tt/r9cQP3JWT/v
ZVIIrZzX6zzfu0CsLk3n3FdWUedsmjqhAvWz+FcHiSE+nPAyW4h2abvfN6YqS5CE
x9/E080SI/AnuwjANLd8X2IqhIjqf6J8czd2B/PO4N0Ydg2Aiy4MYD2DxaP2A/2E
5fCZOM+alv4STe4ehkJjyc9OlQiGOUW6XwwR2Z4L+Rojsu+TawMvGM+hrofBoy0I
HOTKEV1dfMsd00eXD38S4E/8NeUZaQ6O8KFUmqT4U51XqakYgxP+OSFmvpO9SgES
kjrke9ZYGy+PvPgPP8Wzj8Qsnol1frtqPXh2MdMdTUYmV2p1pq+CV41Ungv6QMOB
ntf0tTLutb4IhBlZYcjvJ6FrCQrUJAlRb6qFohTNSgG2FbR4btumI+r/vH5+Hwca
0F3nIx3WjMFtbw2uh2UC3A5L7TW2FJtBnVrtjRAzZ3aqrS7uv+VuDjn4XME5h2DP
paZukNMGguOrdR7rRKcNm1WXzlVVCkDA+FSncc6fuoaPJ0MeijsGBVYXakMMPuE9
wvD63UioT2aLD4PzeI5rxlOIUOl9gPeX31HCxqjD52OmyLnHCwnSklqI74EMV73Y
9clV7rRh+txJuFQr4K69q3Mi1/UP8NbrgJDZ2SY0052ajbEf+pMcFBQIy97glvdA
/4bUAnYl0UUeEor/2Rmrp64QGILcKf5nSMT/Zgjhzt0iq5v1rRNHYIei1XvnUSZH
Mf/taw1JkF36o/PTipKA6U67Rbfvq64+9b4gpv1dTbWim8LSff/pvuUEZwR7rgVa
wXl9jC4z07yIvoXM3LO9alOYzNMv5+BPrp309MRGdBvOJ/iP6gcRm75QeZ902dIp
aBZTP0P5PIY+j8LtJVLIVsI/klnkV0/xBicdm2frdMKinPcIj12KbRvMDWUno6zo
J67S+NQxhqyJD5X8mj4nTuUmsBYfkCkbfv84zjerIBExMF1OAYEekdIfewK0Gw6G
BpvJYPqGbZUEaS6G3FKLojh+on7WkQAHTWMWSkMO+mW634gfNz+0X6HVORmeJI9C
UH23dmqIN3ob8WqOR/fbDSb+iP/5beXn6F3z9+D+YEh53GuY7wyh52ZqWAiND61m
uFObEi88OZ0KfGgG6xji7tOlnVAq/+tzSANdk+iREeYBxuHwrOti4pi1+f7l52hP
cYxzLXaP/gXwb1Cn9bfDXvFdxvr8B42ZTnBNWpYc8QK/xpF7r2+YMYjToopVfg48
dCwXOZJV2hJrfSOBu0CZcp55OMmpNoke9IWKi7Hi/nWLW+Ssgd4mxViP05gjNBB2
oh+/rLmbxTlYT3l5JedIBvIRPVipLeCYgoeXKorJecUaVVmmXOk3wQ/BQgG6GbDE
+/v1aiNrL542W2KDmDmyCX4/kl3NjgYHojAwqMri84TDXMPr8PiMh/vJNizgD17c
skgYiNRvzSbqgGeCajbr/zbj40xn2gs6ZoN2JjtDAUyq/ohIIFtZoGdi4RDYavXf
R4BmWuqKhPm2F3V0CW7iZMb1wFqReZk1a7HOvjg47+1h+tNaHELzMY6QHQaxTZgg
WA1X/+APCyGbfIoDbes2aF6KG7bqdEEc7vN1UDtRl2LHq/Zs2bpm8yVoMFCIen+N
6+msTAiTRHR/GZmCc8zT5w1JQaQo/O6DZgzGuyn6TYw2vUjhaHWtcH35e64r3yU4
1HkOa1PByAIzWATYl0LmI8DRRok1Sue+2o/qVhvGb06gxuWjNfSqfUQ2BIH18CZ2
NM5IEm0ipJu0CMrcKwa+QUjUMXsAehxVt+O28/G6B4dH+9jz0Xsfy+D0kpZw805X
XSitnjecmAz30cCep7ikqJkJnMeZi3uF+18bDsnRLfdR+331Z0p+EjJ0hj6cKUpk
ym9WLx+2/ZyVpvwvYwr+UMRnh/3kXBJvm8u4WMLhpsyQ3z1gCDWi6sekU/c8H5J8
yB+x8EUkIfjeTeu7ltHw1mqfRZqTSSe0r8WKZOmyXb33bTgJ+l5RL/TzoW8wPtPQ
CEfE5JaG0pOf3YumF3AF7yd+frWJ9XJisXkHl4uqBywB2MTsLiSion5wr6tpTsUx
SKk10+RcHQ6eYStnGNX/1/hHsR/+ey0OPuTZo5Wim5JeRK4cguqJOWDVAeJCjgks
KYpVeykcwkCyEmA/ZM0T1L5lwT3mUVOTk5RJN3p5snnDpfELI3aXFSvPpW04ab9L
6kOZoVEUL8ki/bKC2cwzBgNTZEnj6xhBJFFdVPihuNwG9o7VfAI/1LuqQdxoaHWz
aGsnR49flJUqwAqPr5TJ49d6hP8fVO6d02+Crnn7ryJ4AzCS2dQ/SLP8GBhuWUJa
7zgnsrFzJTDVyxTKwhG0wfSy37inQ4Y4o9bBk8mX1VhpZXeZiCHo22sCoAtFLsJ1
5WOSLSO27qz/Pjr8NWRAN2XafdDNgvCUjfpJSMQVdF7eUmqCE6/iYwt7A8AZrY+/
ET/pwxmD1NHvsS6O1JkDE0JLWy++JVSvK2ZgA7uhuoWWqbtcdYfXx6717gOg0Ssa
T0tx071xC0Gpev0F2nV3fu91nR1/q4YNqn1V7yeorDJhxeaQh7iAMosGGmm7C7+n
wOfuSB5lGpD72076tqLmLo2R8ynCK+Bj257wePE9SGoscSxEvxaAv5QkDmllNWjW
tONJAGjEQfTu827GQZ+XL9P+gwcBEXV1DzwwnSuXa/wwQMCrASyXJpw8mfhY55G9
ekdxNA2B4QWSxseUb+tleT8wInYWDCKczBTlRyU9cW8JgvLrVpMwFuWP2OB9JZCx
xvJx+LnZqBalPANGXYfH8wqghg19xCaaSElElmkCjeVZM/vE7YB4AFsx4ji2r4mj
uWLYC+V+D854EIPJABB8QsuBvOjguKXzUpEPpdBu+0bd8fmFM0xyGDKpMCvXqCaf
W8d/9+GP0mXWaW9wBS3gdSPdhtlh3kSfmbw9BAYocVsjeFHvFi2nRwKqaJM+aZeS
BuD47H+WkMi+JNfAw8dvEJYAbIWphJ63lKEWOas6jpM2yPvrreIZ21285luh/EbE
0FoOlWjYNgBS4E75ZiBvhOgg7nVVYnxONMta7IlGI+XGJOej1AYLzKzMsOCTteNU
vmooc9dAhQnxoAzE6UGVYJNqoWzoVMgbnpTLDfuVG0V/5cS8zosA7LKqqb2Th84K
PTQwARdRkITz3xC55md8Hwq+nu4tMO2BDF1hzCh6tqSzl0tv7N+Yb982+hGE3l1w
wJ/lnuyBPnn4+ZSJhf+AQe6J2mBwFgozX1c99uly/ALPewuGkwaXOOyvfqyCvyQg
Ow8+tEICqrTylXiQ9LFRKL4d1p9xbBUxoALDoLpWyYi8evhV7LrCSQtcbx7pzTNK
xol9JdnU9u13/9L1AjBMolqL5xKat5caq7KGEKifMFnK4Z1AbgMuRkn7jr/EjhhG
XyfnSxI5nMTLpKlA9m5W62s8HLSVE0m4LriTmgAcLYaLqUX1oV65VrEikqJsXyuF
kQoq2c/GobhH5B87YSwzHO/5e5YwuwCWS33oooNwLGo5KcbcMJ/qejKLRc5qxvn9
ei6mftgImiN2Od8hVQch3nabe+gBAWDX0mG6kpeKUzo7ctCbJTPTYLHWti9FzeKG
GsPpjRtCzYgJAVNDM3tbNxvhQU6vWY/fBi14eJaBEFZpxOHqOSMsKecZjMDgGGzn
dvOHFYCvqdP/HnqpZLDXSYXZf/wN6mQZFMN7geTTx/hzxZyMalZLvyP8R/Nsm4L0
5EJFiA1gkPEYBUo5u29v91A9E0MCeEJE0x+GkiY9eDA5o2+h+JiUJUee88/kDHoO
j6yG8oOhoh4qza5xkvzVzdibMycq1a41lS+dzTvliFQTePHukks5QNwe/U/XYlPf
AnB7VC8LupJoUTHP+e7UL1mJ4lAJdqIByREuv/z8YFZWtBfDXRydbvilxO3kgfuG
DqcvtWfOBcL0/2Yn75fBrvev31Db0mGoj0ZjuH9IsNIXy7+hzwko7B/s0RD4AA+r
ZrapgGqnOSf4fyteps34C892uC2ifcprMOnejruuYkt3KibY5tZtKcjGMP4ZzXat
g52Fu34dY0miGcEXoAS+rhfTKfKbHngLG4ROQ9rn7iHrg3aDAmnlvq3KloWOHie9
P3BxxdlbSvx3Kv/olzXEH7IiYuzY2mzU8LKQ5awir3PpLUqnccPv8cS4apUI0NFq
R9kkaOQYNyVeFfRNSgRBNxzltftbepPCMrFmL+dWRO+RrpjrPB1trOhWshGbauTA
/jFTIWUtqrkTWuj6bH7FxgK098vS0f3USS3RSJ6oxE7huTo+IYHi+OwmK37CQj5r
zyup4xk2PsdCI4N1MU2sZZ7Txkl+iqWXv5eRnANoCVO5T+q3WWawMC1B1XSKWPpV
tydG258wAiWhegyaHrEbqBO+zGEIYLUjQ7UgcWODhjl+w7AutTsdKKrJ/h4ytaeH
v/JvUi4F34ghU+pzPgfqvFUBoGmfGKp3vq0oIZBw2yIh6SGni8MlSO1YglQ1WzcQ
f4d5jLwQXsFb8YT8XL3BftnsEsPXh5oPmxEGcpp/3Dv0LXsD996n8pUNdCf4Kdps
txekgHPfk2QW92z9cJFwZRUrZy6RJAJjMPKIkxVUEW/AP9J9/bvMey6J+dvpM7gB
eIqImaorGbHhNL/xDzZCKp1zXr6Ult1Cb2KxtEjReUWBNkroHNshmoH4+eZkx+gU
mqrFZOuNvhzgQutbJCUJU4k0hFRaLsG8ra0q4SgbHf+HqbIwXW/9HufVFyur/Tc7
rbrUMPz16KFF43mzSrKECdsPqWEnOD2VSRGo49ZKRHZ1RQwJzYzWK0bn2G+M6bEu
ovqw/8bMf9aSVRxyGvUoQ6tiYDHS7Y+Qe60Y3gMuGYBEG2+TfmAAalKANFzjbw5Y
lajoRrj6eTSWcjZ6Cg+iL62A8cbwf0E0luynBZyOYwbh2o4RGxe3Pm0BUsuA/g+Z
xOfgfnyKDW+/nR25ry06hk1hdx8FcFIIKB/KG5y3VusLLRENgLgqiOr5OHjycz11
IX8n+8WWDBPs7t+CSKxaCp1LOACkJXHLrZS6pvEhWhUng9DVCPhs/N2KBfuhzxAz
aVCtE/DcZBP2oOfuY210O/NRHl/QP9MO9Ydwppkx365Dj5RstqvBNMLF1ap13EnJ
vNgzKRnTSW4boAXiighofqe6ykPneQoZKvRAeixoaACAYx7rN7nkOMfo7MKAiMbx
DftpcVkqrRnkX7K+qZOCb5E9cmEREi8bwAM4lI9PKcvRkft6DRHAXFeMl27vGWS3
k+UYEgay2j8m9OulEAyNlTpm2ucP3SMk+sOmj3CE23kZZNjPGdaWHD0hilCf5Sww
3ij3VVtOF1ymNwyKHfHfISJAT2UWmW4asfqMycNTn88rL6ml2B4nROXbZ+bFmB+n
nVSiWHOgf7CXH8kNZe2G6xVcflGYWGZ0HrzJulw6kspnWSExPkM/7Uc13CI8ugFt
Biy3EFyzmcR7rI4BQUeC/j8EIQs80lLE5sUa4YvSJ+q9yjxpSZTAYrF5Cj4j8yRW
D3MQCb1C6y1UQ1BfK6RocMUZ0tx0PQyhrbtx7N1g2EzTGmMJ8lqJpGA4VrQf4Nl7
+oc3onZuCIFc9fa0UCb7ySRpWeXUshY4QVR0w2Enqm584I3h35hBeGFc8S1/bUnz
pLAKQPfC98CZaV5mG77hEydqhwnxsVYoP5+7+caux62PR09Hi/QSTZIQC+vDOanF
CgG+w1MAHMHN3DV+BjTLJo0MIImhp7xi5DWoWwH5i+CnbYS9f1WbivOGpIeTRh7f
i24IB+YA/k807eygqtKMqLYRicT+K2d/o3Wq5rsCtK/26cIpGxxyG7uRjOZet5yv
GdZsS8Sx2rorQSBgYmYEfkHLE+uBTeaDqeTYcbvZ26CnerVTjcnkA41S7ItsHa7k
HOalsw+nz/9bK/Ev0F1iYC4bihSGW7BKuIn6Qzo7glrFmBvon14WCkBp4J09E3Ts
KslVHF+EvlbYLy6Qk/lelOqTa3YMNFiawjjb8m7MmTfrql/DYX55Uw7kFXp63G+d
APpKTqiVZBFxMbVwMoA/I66GJqlbdnHkz9NDD1S2TU1a1/acDNXyHGw9El3F3zBJ
tK3Ys8rLSs8312SxwndsJvDVQQJt95k2QF3zWnvmI9FIB7+QQGtTIcch2x0Y8XzR
HUOZl/6r3pY8YZDNpOp5KNfFPmIpQncGYSxFpHf2bF8/4rohYWPUpYf8zV6IDFdk
2NA4tVZ4+zPAn9uMzSwTAxFLYIanuSQa1yVI+iJXQrUbY47htylEAHg2+3eReuDM
oeKtpqTjqBH+hINp8ReKVTuFDyRtnNUymo724+Ur39hP1rE98jYyDpRWjqIoFOfU
lPOm7VfDGYjJ6FZauN9yfRmBdXnpI1500VsNTIgQ44op0tLwlaw/cybYmmarf9Jp
Q8EySfvNROraosuGqawv8CRyff4gtMjxkozBX4J3SiLiK8tIKVUTvxCk37Nwq/cx
gOlvD7NFffYJb+/7kNH1wCZXXt2awnIFZckVFmIeFa/sn3YNnLChDct9TXuHucbv
SN9ccu3j6w9a+Y3spRB+qB9M3ZdYL+cbefg/cFKSatVQ2cUV7k72LWFa5Qizq6vv
b/157eyfYhRw7RTCSxMQCbbef2yPBVMcYiMdC2t/1xjqmwj2fAbf/oHIxekzqJpv
Cj++bf6Jz1od+PJmdmQ8DR3cR9eWPyGDfM2cc86G7Qy4TmDhA0mQ21G+RJvjtjoT
R8SL1bu7ZdYxyjfmnRgDYDNS5GXzvD30/X1BwNEAPyq45G5VkvUBDDv5WTZ44j89
wCCduuH5oX3BBty9LKL0LLUiTyYLAt89t2hkC6JEpfMz8CQvhGStorXimu/gFtUz
V7M13r9zAtGsLycVGoEdWDs+kYTjRUiF1VmM8YzIsSJfI9kXBiVNWi9LJa2mVfQB
cXKeDKcY3HIvW6ZX8RO+LcpdCDu3HqPhrukfhWyBl0aiuKmGmD8R9JXMEn4wbrgo
x/Molw9hPpHSUnBvM9/oaXH1cOQGINahCyRncd/FHIqueqwJSO1AKeRdiPRJsEZt
Kjkyy4wo2jX19C9w54W/JrfFL4gLpfNH3KQPaXun+vq3e0ufHRGetSLqvhOE4XuZ
jyy8CSbYno4D7qXCAEQ+J3V16R5CPb8q5YE9FLqnI6/cc4vFkXZUC/pgOwg0z1aE
phuMUT/DBQ67jhpgLzgCyLlpZzG9SpNZLqn+iJv7KDgsIwKWLIWC6iBDNjR7ttLI
ki6PgHOp2vpODqORuMAoqulCMv+7yG0z0tu9f1s8nzEnVUp2+GqT2sGH3+lG4WL9
n7IMucV4KeaQ4QLCRyL++H95ETcJFVCTtfUNVDXED2pqPaeTISayZkdUUhbSgGy+
ClDUuv2uXkbAi3nAQGso5IfWWkz9gjVHm/9G/jDYiqB9Wi5b5JADJGon+VbN7DgQ
GsulsaQEJipZkOJN/Ehg/0R4Cr0/yqbYtGLAxB504HB9UejeVLr0cR0Y7HtA4zLc
iORaXK4qqlW93myNH+Ve08sHO/Pv793eFq8Pe5hGBj7Apfx8NWWSWZK23BzjrlpQ
r93h+wHAU2NBLjhhibowXdPNrfOK3dzMBYjoCn5wgO/gs6XJVQBtR/0svF1iEM09
y2lkLgOXXDRLD6uWJngNfNCwz3GBzK07COkb8x7dPAcOQFt/ZxvnsuwjFN9qvQL+
sp6SuHr7WS01Z+XQVo+4iVX4MwU4IW6mtK5r/cVKlCCLaGHx978M6lHNx5Uyepag
93OAdLptH2P+r1Sa0ahsuRSaTSWI4FAi6YVFvIuG6ZUwu6bqvzUR7UEdzRZYIke2
iS7X5qROO6/wQYpdQLV7jjNT2DxzmNr5FPdoJ9TupH0sJbTvVd2w7UYaELH9Y3Bl
h7crknXywkj8cVjGXbV1Xfc4Joatupd1kQkjLzmofIGy0Xq35cWtptrSVep5yRqh
K6Rg+8UzM+21kERAbGBFPRQJ3yHKN24y2fRbuGnFm5+Hieft1MVhUTEA6U3IHGKt
rhI7Fnl4uymj/5HudWnbDk/evlctFW/FfmxO4BtKZVa3tZ3JHEvJX/qalN/qRIyJ
jAgUUD8nj9rlYygirhV6Xz9KGEVPhk0SGVbUuk1hcI2oRKvc6f9gbVPpCvsOldzx
GKnOGk7y3dWgGVJDRfga05HWeMMVRONyhrz3syXwlPxCb9NrnbeiKpc559Z0ilNo
jcY7k3yjZ1qMHQpXxT/6tbg/G9bDQvDYNptzyw6adn+NvPGXdhyN7hvng2nRfKKM
BXpqM/5AWk0N1fiSiTJsF2mq0QMSt3PNQk8bSj5MgQoPmrFUsnFLzjpwqgs7KOCW
JUMoMVivZ5D+OH7VTY7862s4TUZwZBiUySa1d2lnJ0KelixrwbmjO7MrUCbqf+jx
Y7lVsmIbS5E46xNCRqT3fvOs0rwmz889E9cPCO/5lRh3TxghO+IfTRFnmFkNQDhF
/frNhJV+FP2fr9kZwiPPY/I5hNWHNMItAnSVqjABug3MMmnb2tsmaA173XqkH2Ya
E2Kq639bFJrfS6JDXebPXy4HNw/hUDBF4kReuWG1/mfhekP5ppVda7I4Yrjj2N9n
74J1ytl0HPbPYYPj+ak4SVse4E2xr2IxG8N5uuiAxW4G2yOT0N7TC4TDZbgcdHg3
M46cBQTZe78H1qU049P7iPQkgHsr1Qzm63hL0V75bdp1WWtV/UznYjO+gYH2i4qs
/qQiGwO7hoT/z70tnooKrgVFezIQdIOKktMJk5BytQY6s4gwocpONPhD5GALIifA
kbQ4evylA/+KhB2CF4P3tbmqqpugdJ87zm7nrI9GPnYEutueeMyUG5xtf5Fg+clh
HUfJxEbzXjV4yJRLdNqvrPFwVyA8eqB9TeJ1UzB2nPiFShKSSWgAcbCrduHP+Pir
slEuLTr0OjHmcE5LcZtt/rBIxmF3fwINRjBQRiL1CIapVpWooCSzPOMsozafqVAY
CmtsKemur1h09Ccumkoc7HL3oNrgXKIwgSG/ciZbjd0AG9OWbJAYeO08jEuApMxo
7FZeFI+j9OwXUwNCx7cLrpodPGNutHz0JqCNtdkIekT1EuNwGZOMak5Uem0isvps
2nt0rq+Uzuf5nXQDORfQOXt52qNtve9d1HrxM37YDL61mbaL449G0uEN102NcxAl
39udWB62jlB+R452QTOeggH6d8Y7+no7BqqhLutzsoSHNUoz05ib4V9xF1fkbiMX
EJ8mbqyv2/hVX3cbDPjaQx4/YB+Q1lS2LGc2J4n4kzzJ97pZHn67XiRnmwRDZ11x
aF/AAM0NBvCX29Qnd/h3K8XPZmNp4PQELwMmOSpc4VHCf97zs/rJIBno2RveUdq+
UzIo1El0+9pAyuGbABBP65WU9gazjF+jWBsB3Jynfvqu0JKjbCzlfDu/jZnjSSyP
YzKrO//it7Qx91K0dVFSEQFqvwf+gbdGUaa99alOqB1uLOO9ne6eWatp1DcSrsxU
iHqLFwn2iyHevR3N1VGg8AFllXCZic9gju3kvDF7h+ten6iuT1ZYky+rUPHOvVlA
zpWeJHJegpIe5whyrDCpD4AF628iqkJVRMqWybwWZvEsuAjU58sDz0TiKsGEuks9
mFe3Rr7eFoXKbjk5OWmPygjilnccUb1JqS8lubms90sZuBRrAUv+XiWubGbmfCd9
A84KeHsYaf9xUIs42BTUW8jgd6G5lEZLBrPp+axmSiq4m23Fsh91dQGG1/xVRZSN
XCFGeJn/J0L4X/dwdLCcKgdIcQS8yhrblcMuR3wUF8yvKVuDSDR6dVX7NM3Teyx/
OxJIT6K3vuXXIt1kL3eLw+L3kFFFHCdvQTrOdgieHyEmLUzafteRNu/FUfO5YFth
p25tucskb10g1ZCOh8JgH+oMRCH/aYW3mq8kp8+C24CAE6prTRJVHK2MkN3NwqQB
itaBtjK9k+VDH/YmDP5ZEuxqiIc/p6oYH0cyrNs+tNbRvYumBKwfey4vsGPhganx
+Q9KKL0kOLZzONdHA70kLfErpdEzIipD48tiCzFllV0QiUrC2RMyU72gSh3Dr4j4
r2nsfvnpenQ0VNlw4d3b/1JJbSlI0raIjxpkuQPGERG4craWre9iVfaWaGBDCU6y
7pyWSURH/zAUDdIR0vLX9/oO26C31Sw1OFsb5zU3VbXzyL05cr2FjkiPFrXvYLxP
Lzvonjm4FYPI0CJoKpbO9DdtNRJ4+wIpqeCvST1pv+KYoXXSpMylCI6CiqI8TVQJ
S1SncAT4mvfJBa2P01/C1cD2tnrgmtmeybZ88qoM0WPgvBCWR65R1jV07fgriMvU
KiijEwHYlCy5nnBv6R7ZxBt/jPe6YjBW/ctdfd56AtddLHMueUl2ypAuygujkr5x
UWMsznjwmGZ9RtRz4ZzGoSAZtzzPnFvkSpKWDfO4wUH1gNPvddPB6oPPsB6e9z6d
ljNfT1xLoVB7Et4qCG1f2a6H64KZ+5fP0dUHDFCQbCrfM+/WEeOVy4UBtZoxrOyh
uQoWx7PigFlmIwib8hUMktUssoCasSI7zE7p3mP9V1Ke/4tHkIN8i7hZsL3TRB1o
TobGHA6zwkokdxt0IK37hF3rAnJjS+gjeThUWd388GMEMokwZ/Jw+97hJpMe4bWn
GNGGx24iznArgKVOelRD0JkNhssmnSPt10rDmaPKzp3FFrLVzvOZs7r0KCqFrdoN
aCdcQ6iNvdRfzdsFqr529I39PUxn8/8eCOmEr+TF2L6EYPrXuwqUOGeVgtfTrNtF
wEn5XQjhY4WeAFxpb//YgAClz9GHFv32rD8tXR6to6hzAOsME53g96P8+Mchq3vi
S0uFatlQ/gx7++PuDRyP1G0TGHAFgkO4LjW9XwmzrUer0k8Cb+onvB64vJcyrxte
ozOBGTJHNlzVLILtjN2atRYcSvs1FTUp1RyH0VuJeVvjLynST2dtoigy28IShcS2
7RB4yq/iRu5RrQ+PmocrEWsEliQuUFa5oHahsuFwQ/7DltEkYh8DutkXsbBVwzyh
rbfzI1HNNmvP1rlw2g3xKHae+pRUNaG8mc2kDMvmlibMt98CgC2UGwWGLFMtjyZZ
6pudEP6tNIUoPHQLhc5+imP6DQa46eh2vfZae9lsEbyF1OrvixYP5pegdZ+nRYoT
EMtflbZlsHJ6dEB2xeTpOhTzeVYYMsPqq1SEohvf29W/MQQMQ+snVjWP7UlvDhIh
B0v2fKSTmLcfs4ve5jNBVS5up7riOWIq2Hq61KoRYbErulW1fzz/7tXraD0I/J5v
8otReUcXaWyC5fYZJYZCA9MPLrxRui0xkCWvkHpQSCUrLyqLLQymBzkm/LtMaIdC
GW2/Cl5GRX/1xw3CkpwiYIXTpB6foWWRdatX7cmO5vOz8swov5V/IGwlrcabS4IJ
6o6Mygr1daxCGnPb+Dr8/HedE6WIROVVsEqKPy33/4BKh3Jv6Rs6mk5X4iT0am0h
3gXEgD/bQ+BLPc1W888oxDM8wQDLMkccIHnriok5jjMJ4V1aZ1il23loBsUs9ezw
+WQm7XnqawOjbz2tj4RUH3wKzEWbwFhwZ5GH4w42ydG+60PjN1Ur+ypWdQnb4Lwl
NRCUQfA9inLMxrl0CNthAkAca75kN15Z7CaT/zBXRJyNUMePzqxUWXIBI7L0UWsA
A96iAx+C2KlWvKOfNT9MFj7T2x/w30ALTr/Czplp84ZqJ2grI6YU7w+AFlL/14CD
hbtgVfJjhhlTnvOViG7/5Yh9JLUeANAtBqDKPb6dQO6eFzeRcnWd+sDheZ8XVFFM
5xX/ZIgUjBH3E7sDRf0awEu8FpVp/Pbw2qT44DZF/beQg1/8KksGMx/Q0HRKDF+8
xmGdxF/JNBJPSK56wVpxFwIP/BRXDrLnGJ1C4WoqQ1yfwAtLo0b/Xxa0R/KT9Y+P
BPyrH9qOIbba9R0YXVibinaUU/hHtVcrbdbiikB1uuQ8mt4YXK9AGoJYsN7aKION
iE6Ph3GfCqVA/DrY2lKobmmd9h5Yevfjy5TEedSSZbg6acXjM6rq5XWtW22BIqRI
OBlxDfoPi1/z6BfH+aAYWQ9nmTxRyogQjyEJFPrcJMdb/lbb64JwzSKMm9y4p1Xv
Mbups6Kh+buw6JpuD3xEaybAB45DwwvPQkbGYSGlfCfTkpGCfk404SvWHDtGpKRg
iErOPYhNTnd5wFauxKv90IQZ4REIfDDlUQ44i6dAex3R8BJH7YrZnrUU3PD3u6+e
xsH9g+elLUao+rimIk5gdzgr6QspvY1No1lvBB4ESv1oAB3VXiIh6QolbBVfWd4X
DxeMOoqrqX1CdgDEetvg/9bvd3UGgnBpH4GH16L32SsG/MopLxRNwX4MUnB3m5xf
pb/w82Y6jO1EZiD7jKg6oGBwwIvIRAv7R80ehyzhhW9vchLrNB5yPyZI3wztzm5P
DlTXLzsJmbRkZrPMiYknloerDH9QmDXTvJ66rsBqqFqJTDTu8gJ6rP+ZtXC9BJH6
ajav20nRFSktU7PzskhWE1RfGkpQTtQAsZqPMa1VgRhQTaQnVw53y5jMzT5gouKe
aB0fz9Smoe33NRccgj/zixlZbN8FrhBczSHfxwcsbmisQBQJklhANmvz3gzgGR3h
g+2FWr8ewumPO5i2rFXmxKD0bEgJctOFqeGtwL9ZyOY4kF1xcVQG2ihnLh5fG+Y+
1PotghrxaQC2GsKUHG9GQOy2J9PeNFf/gPRy+mlGAfe61y/BgD6whvhIgbNuk8pn
TznU+7sQ6u1cN8fNN8fuF+nVDQh+ntvklvtBOzMEnw0eygkgQkGs0JOhBKlpQmXo
2i8IOk4XTZTErdK5nD2Q1E0EbRXizg1WgMGhzyqOjbrpGkhr2EeE7Yxh5uFMRlZ1
MLq9f+/JUF486IAhnkoiOms8vngasqhuqiTnw0bocv54o/dQ00zd2Gp9Gevj4aIx
eiqKgb1mVCPJUwKiushvtU/PNkWhiOw8/AfpVmJGYhy93dmvsOKpRgdocPVIgHBl
GXQn+uE2602wGHZ65jb2PKhKGAGoBrQG+6QuAB1DdgfAt0g8/5vgmebwnd4Hlr9y
r4CkQcVvqlw+AcZmBlbSkLLMdUSrDkC/uNf9iCRKwuNEbHrgr5eKr2snMilMYZmt
awQn8ck6EdIogFbKxHG0Ym+xLieocc2rrdYWa8R/8PnO6GoZ6AzwqAk+jwwob2lx
mUImbK1rW04F669N4PuqacZ/Yx166/u4oB3VGS9t/bVyB/ijVSrnPzijkmSlFLhk
aI4p0kCflK/SXeNxI7djnduydsR31DKSbmX0/hSgRj6fGkALQxp8tDQ0Ad9rHpzK
b3TX77yyyIBn+J+eJ4e1SX1H+3T3yXv0Zu1lT0xewt3RFYekXJATmi+hP6wz1Fvd
G8HCCyCTR50qUZxWD6J8Vt9JqNSbQ2krhuHCoJ4lKhj9vxe8pKGvcLD5vj2slRQd
3Umbav2OFvXJqHjPj7Go9lV0zxunuFOFs3IjWQb9AmVC6vgrJDalLH/x4mWphUi3
2h02c7E+1f6FiE6Ca8THOfa8LSDK53Mi5jaVorTXxUTohHV8lqm4TE4OEUYGX+WG
E/aRDjT3pYiOgCAfd85AJguEf1jfkABp/MjYP0qiTyBJ5hsJqaAPoueKUT+SApN7
2G038DfenVDMRtkMgBMRhO/73HLyNEiDtUAu96q47ydqXJTThs7m0GH0Uc3p7E7v
f4L9/mqvtyYggoANg+2jkN+5C4K1PbL9Hz2n32+yM1WUxtyWETN7INwRufcptT9k
BJ3/XIZd+axr46puI6WdDhgGan8saH4t8zkfBwPMekDI78ou3pTjoAXhEwYk0aMc
tFvNDnVIsuzsOsVVuiIqA4vH4w7v7TGEctNPKzKC0Fcz95vPa0vqirOPkOgQhEeB
GN1TUqVKRXYO+g391J+qpCY4GZRDs+wB/ZvqiXksL93MhwEIXr99Cv5k4h5Y7iwE
yIws07YKELvLXCJ5pp3o2OguOe232V9RX2u74GAIABpOyHeMEjr0jARoitgVbknH
KLEX4nQf65n2QmIrYycNkRn673vCXL6ju+j72Reic063FD/vtnD0ovnsDq3OBoyS
5m1803hni58KwvsskxLngU+P7cdiDVenDxO2zbEEe3ukksUJe9mwjCvCQA4b/vnp
IhxotV0vjI9KDACmC3SS7h/PBADnEfHZaQo8OWJUYCv1ZZM9NnHLs502miR5BD6o
dI802O6v2XXV2LrW5HK+w4Cnm/y0BxRSQMGI48ZvPpTz6WkVvHpJ+e2sHIWDz938
ifQUfQAsSySKzHwAHi21aMGkVeulfYAP8a6nA6hQK0ETacm9Ko+djsPAxDtGg+zw
N8/WYfAtcrJnpGn5eBybhRSGQrYiawTtuG3kaxAIbEDGGa+Se6KmsTnbYdqRRHjs
oKw8updvHZIEQoLDupJgpWPOm1OtXtepD7Tvxx898L99gJwgl0xQG+T8gjCt5wop
JwpumurXg0qy10fBGUpb+LQa9j7Z1ruMXjVmeJboM/JRUyjM/iNmW/zJsfcrgCWq
a1SD0Te5T8vh3OQ7tYuJ+VL0Wu7eYz6mNpg3g+4id2XxZFfwyGedT5z9vzm4lHKL
FQOu2V3C+AvTtWfBJV5e9UvZg0Ay/+uZyIeEpfdUWQlexb40VQTykzGJFNoLB/Ti
PvkchGhUVHds1nfiqZtxqMEdrC45p94WX7oC5XFGtB4KhZDX2eC5AlHzXN2i/t9M
uKFFoFDRuEtoS9Z3HJMzjJDsS242ZARHOkisy04cFn/mMDUw0DsMODXD8/V7rgCa
mYIvQOmRWzk0WCuj29AdKIv+NOeBUsJLoChMR5KIsh8Nxn6FE4nCH8oc7VapMlF2
XGxXAKFlvYajat5sBNTGTWzX3H6tQKe9/6EVQfMm1atbdfh09d/ra0IB3rnoodBY
i+AplcVUC2nQAJQDIMAUayXp4PDxYSA4ZoY2o9Vj1myAoIIcZbD9A9zUtWXPU8om
GdBG4zpLP/xhto6mlsaPrMp7OwRWZQwduoU8c4O4ae+gsZqIVj1Tghel8xUmCDiM
R5vaRW6RqO7D3ti8fpBilc/re64sWjF6QjEDJEo1xBw/OIcx8+YXfAnmy39wd6sC
3FRnGBA9X8o5c+Tq0qH45Zq5LdwodBjFFi/gDroKKOccB6GQrrj1Ud4DfB0LYcrN
5Grkm+3K2t+tKK0TGIQNjdMTbcaBAOF9c+5IOJ8nOl1B4ybeW2l7B3yfKnsH6lc3
SnJoShrtWeOVdAquNPoE9ToYUYLqPsH8uy74ZlhoEPoTQPHCa8OQTPXBTDw6I5DY
prsu4VnpZSBfnKGO1+RPjSbxpj20Ugme0Qs3HhEhf/IiZ84D32svsoEjuCC7OCbN
SJcNXCSKMC3qoOvonkvFbK/wGNRbZZ/49t0pHPrQ3hQhzh/vf49Zij+sdzL53EZS
WAf1ulFDJnWrSxiV8HcLZkAmz7MzOddan4MQ8eMp5trDDFmcS8konzjL46HWofpe
CMmgmD/IKXBY2pQtzOOLNZzl+1NryMOPlWoBfJedCiZ/SYJmgD8Vv3gBi6j2I8Gd
78pHdiuQWLK4QtRcX3SPp3XGrKYU2Go64hXSUUxzdRQP9MA1bZHENbf7hkv7Yr2p
JrPtW391LcfeFUY226rsEc2QdEvfHj8qYdtypJUoKo/SDz0LnoaY6PnYxteK2vXv
y9dTpDV+4qyooyWBDx8jnvq/u5Q2M/3tnyK6vSr0VpkO4V1LNF1YLGzm4GuOAqtV
tgRnuxAhYsEArUBbYIMfQ7PK5S9EojO6mhwztvEVrtv9mCyE4eBUKSJWXYLP/Y2K
3sd4txigpqdn+zkIVlEelWKBDvD87fBOSwHHPUnYIOChOoeJlw/5yZMKIECa7XjK
gROZfhI7QUBiy5I23NeFySR92kzxK+o3OKQz0UyaFgNTHQN6q7YebCoX4xsgTgCf
WygRfLtIUH3a4WeHE8RGhOf91mLoo+Pz/MTMrN2vNqM+ZwEhJFpAJ+RXTDsMle9/
zQDbVsDf6PKe+fgkf13vIVApucpfYZmwQnChs0ZfVzBJQz8e5WHYrFMUocqLeqoi
dK5oNtFK7ll7Mci5BkBCSkv4+ZYWZJsjKOTp9A8CEkmd67UjZEsBGyulzPfxWCeM
ahJLsE6EoLZYPX3ZhMB/e47Hf/Awhma9ZAN3+8OnyspRSsJtQBKNGabsNZgFocOA
RtO5nobLWQiejBD2JUCTGHCa3dBbFHuErIcg/ffHTgO3vPbN8e3z7ZaDT36G8aRE
T50ymjnOobldlKIL8+TKlY505ag6SBf76Ss+DnpZSd+OtZjjxewrNBvCSbAD17v3
Pq7K+rnk4rSYbR1nZlQHeNPWQPrP1x7yBV3gywVFqZzMf16IB24U7FapZIAgvPru
3J/lMcH3J11ZKuaVo6DzimraQGuILdwH1aOqpYBx/0OBbnCLzmQH1V76quh4mRL3
zPWwJgynCf7710Y5CUmSQXqkJgOD7dpKq9CxtPMJ6qR2SYdM48co5cvFl7qPGSWV
1kIJ/4KWIaEYdZgWnu/brzQR0CuyU4krSDMT9DS6/vUzjW5Zoni9KIznlBLDktmA
+ks+ZNnwNavV0X8ar7aLxJxG23BIh+HOl1K1wfV+IT9DhKRCXxftHaT83AIO7HbH
dA3osmp77onkc4yyzHB9HnKx4hFsm3giesufafo+dplkySb+c2NIOue4TOoOJFxu
wcdVJ6GsbUFWYV/ekvdVtozq9If8+7qhM1MS62l37VEuEObHUSjrOk1kbOuFhwb4
JJ0B7d5L7wy6ZKEao4pxs6tztKTsv1JPOyxE0waNP9W4vCjLeNQRz9PgoZoY2VQK
X+7RA2Q9j4Dox7oRXfIm2FjKfebC8SJYgiZizvJZ+A3IVAl+ejwgTX7VPrMcYgB3
S4CsLTr6pDt9TC9A5zD8Ptz9Mn8Vk8X8bxUaBYEZ/exHYkoXTBcSSs0rTBN54ZbA
Hbre0sBFHatFPMyehk6TKzSX6gOe/1dXxYggNtduiNy0kWSkh8yVM3bLdhTPS8J9
WLbaMZYh6St8l9nCGnMiiS0IYtu6mCDan/XmusfpBCvBIVvSzCm7kpajCFJ3Eqtt
b9Vt783uu5BkA0ZLRzwPptEUD9MNjIK/DWbN0LwGSE4GbQMbuXrOu1yxzQMxwGvM
PgEFHebAHTYNnEMA86A4HDJFCZ2vcuJwoufBqrVar7OxjK6Td6cfq1tzA3kv6TIv
rrDDwdmvY9Vp/7K0jORreoaS8CVnpZyPfF8zRbfBOyMZO+MLMlay39tmvzfGNtx2
WkGhv1ZPmLRusUZIPuxhzZaBCVB6kjGpVsP/ejrf+UuAGoV6j8iZo+lSZSEdhxNt
+Y5ougHgAui5YCwJYHcBgpheuqv6HUAozTn7jhAHjzKvQBJ+TsmFxx3s+Odeltmf
qD5m79VuMAVXENVn2a7AXTUI+xnt7pYSfQAdIlX8s9OMx7tUKtCh7c3f6atco8bX
R46DQUlyPNw+EaA5cykgST+qnJe1Fs4cgXjjs1IGWerCbIdziA4s5acubiYzqoJC
wjn67cSvnvRzLG8WLui3+cEDAJ+FPnYzIQzRfwck8oSDyUHE4sbcY2UoScp20f+0
i5odcILfTv9M+etT76nDLcn2LoA4G4kDfK5g0IbeabuPW9vTrYJ9wgqMmz7HfBbN
jyiycYlMoNfPX8RPsa1tVlUyNcffgXpSEnKfpoDtJUUOdhQbM1cqqlID1EeSP4fD
T41nyD86VdHQHDGyR7iNyaco7a3WusUZGOxF2G4HVrwRiGFOa73oZoGnw/3RvsxH
gZrNVqkoU/MoCwp8M0ce8dnW5hjJDG6HRTpViR9E6C/5Zj7AtigDVqKBNdoHCv5B
Zwk+alMZUuiyvHTixDTZVNVzvldB9W+2rZMYqjjF8xBKBo8cXUJKEwngqUdDd/Ua
931qvXUDpTSA6q35rj8ZwseqQ8BXHHDkiXc4IvrozpN5uAfAZ91MsxzqzXX65wIQ
qsjefHdIwFp1Jcwtm3AIo7ZMn0PllzJAgzpJptzVXjB04z/QyZW22PNkVVMki1Il
9O7+Hcl27aJJOw65SUZulpEuqTdb5s7Towj2b2hf1q2TaQ30AN3NynDGxYg1djTs
1JL9IL6YXbq8OYkvjDrcdKsks8ToYw6Pq/kbXQclFM8NN2xGtCRyUI/4+2vaGy75
+XuaPrV8CE7XKOvyN5tT5D+4EmCqi0sraB33zp5LwzWXft9TewRcoAVu0JR0MwBj
mB95tBtyIctWZzQI3tvUzbSBFvMHLnVeD6xRgcfG40e82qK7giLGgQ0CEoJDIvzl
uNmowZAA4yE5AYQ36eKbGdTDoVEgEsXU0hf2W3I7NI1cAicxIf4K9yudPcParDXQ
wv2AZ62nx/el3wtVmRKZZWruqJ//8I0GEp7PXwncSFO+r0XnUdVg3e9Suk3Tg4V+
PH/Fjo/KSYIJG7d6r8xWabIBkUe8GQNdTxOfQrVtGgcsJYBUh3+7jw3fIbjCeE/A
e5uEwEC0eo9yip9bjuPSfXg0hWb4CfvaaK9R/0PKlesDpnM4nxkwTXVC8ACiLDeN
poRoH8NDT6tBhDwTDfMVOgsmk4OoGYBC4Nyqh2KR3rBC93O16jJRX830L95rGMr9
iR+q6DjMMLrgo7tCYwicpgzONUvoMxWHP4tBHm9rCJ3ssorwpIgVJbMiDlCsojby
T4YDgYH4Bx+zaBE9Yd6MfpCVIG5druUT6WjRE3atQUy8YO2QH5BMUJTS3/8H39j5
NGBZzSv30VWX5eduFbrQwpyHHihFqmKjtj9NE/rmbDpVjwdLJo4cb3SL1j4h37/F
r261scpiSQM0QtY8A9yNtGEge2HPvBEWxTdn7NygLQQrhRLb6QD6WSVisMPlJnt4
pQgjElgs1DF4kAxst8ppy5JoNv+ksZIW1YlpC4keXAhvw2B1DESoU7gvFxzMmCPf
oG5xrDYwimZDVuGQpCKdHS7om7qo2i7hL1YFx0kZybbo3SNTG2kfEF/3mkDspH9v
stxBS9yLWawEb3djU4m8ORELfiRRu6a+NMOZjvCa40068eXpDaN05AM0NPtFg1c2
tYiK5vvdtmpvuUpknuD80qYgi3pHlnygnYI6OBruETQPzn/c0Vz6i/A21N0LUwrf
P1jundfMsRtPr05hsyMF9h+iGyqAm+kbSJ4jWjxiP8c2/YlXSyuhN7h3pQP+fdVh
XMcw30yOjulZmMjllMJPa5aCzPafoyRMBC1DtyzJNLngUkJ/SR/vqkLWp5UvjnoN
AEsGhdADBYbCwt2HIDLJIv0LHNKaBJG8wtzOEnD3QacZoZ02WyD9RpLqJsEh1kwy
9tlDRKk5M/4ggdjKW1WMb5mkkgGAzIMWwwaSnGlZiha12UQ74HJnipNap0gBG+0V
rXCutDaGpIomr+PVY9PD1td9gTRWOa1BhG5116BTpMokLIfhdVpWkpqnU+XSCV+4
pXPDdzCOJnfq35LcFqGOEsDWBOGIxVq/I7Z5hWuP0GcswhQEb/usVFzEUqxbyjO9
qVPgASREwJYXWlt5MykSs9RBoWkzMU5P0jEjjv2UvjFM1mIZ4PwstcxlNxn1tPll
Oo73vM1b6hPvm9yk2YpOX4TSzgY/TpzCd0VOLOuWU6TbqYAHyR2OTpocKHOUCQa2
VLwEOFjwuwgGACOCZ26EaXJgzELfA8pu+3UPwN6HRpk+JNSjGNA1GA1MMF5SHCp4
z/rRJ3tgDzjTCpJ386BUpAgplWWzwAi2PrtdAb0Q5/NyJtxPBnmNuOmcLjmqu/I2
y6xh+7Ex5nFIlXsnNkaqK7iPuF76BBactAXqxLyGsk/kxLsEsXnxch6j/0bj/Yyh
ySJcJ/P09WXdwUMV1Am+xdtvxWBEGXl+rFdvLYX1w0w9L0oGuUjTJRGztX1qLkww
ALY975bjd6SgNGfoHqdlBe+ZjjZqebKQugt5rBUbpzzveFqYVNuwwjUjEwPo5J1a
/YNtZwHMb9xTwpkisn1uKJYVXgRAK7WrOOOesXDmlZW7wmq51VEj4Bk4oOTLCMGa
eHZEIcSEQpPIfW3K1sYK5vB681vRLgAsCeT1vjgfRcLTmP2yNmDJuiPoVjKsu41m
TOeic6DWbzuyeKUHAl7d1lp45tbSCOpsicewFGPm1ghIxn24RNgOpXxcf7SCI5uB
lnGKfQsTeffeGrgrw2kCXykkamrX6T8ucdcrOadFxgEh0CV6Coz9FhfYawkiv9Z7
BthvaW7HAX1XVTug3K4WjmItaSgDnELJawpWVe5gwfcOLpA8MUUTJpEJ/q1grKZW
glXDO5abX6cLL11AfSjaNzelYXWzK5IPx5y8/TsSm4f2uScpi4Wpt0lQvPSX50wu
wxZPW18VBvqu8XbYvpP3skl9HE19AdFugVrZ22f/lN26LzjkogwAOMEtiD1FP5Xu
TZVikqLrWMkl5hFgFuMylSQ6fx2HwDnTqXLO78mRp6wHcYNDr2TbFFfHf6CQS5br
AfCJ/8/WhBJ2Gq5yImQ0r4jYYagxf/dHQ0aSf3BVmEg+WY4fVIV1aMRlue97Uq3V
C3cBvS6EN+g+AtFdf+QtUMpKGOeIO67YZh0mdffIhjPrWYWR/RoloihK0NwNT3J2
5kjCo0345t5/n2K+difacoTMhfS4A84qZmT9I66UnBcgjADU5QOHMeWSVVJWSFvx
Y+hXNSfqatJ9rAd97PaARAxe9+P3D9XzO8YthPGI0t4t6MZf+T5t/9InZtKCs0dd
IpLmG0RNbIKggQV0r5C062r0bX7qPZW4hCgiZkbNveKlyFO5JnO8MSYujQ/nIEhP
QQhLMIWYgrIFr6N/BldB4RJB4awSoxKwZf53BmRVkTh5zohNS6S1yR98r+5ovHh7
tz3do7hIfqniUhV6Q6b8v7aCxXX7WTDHLAKFMQdZLxJhgh1rVfJc50sVqkzztNDm
T6cP+nixjoE8lsDBlJGTckVKsOFH6c4UzbePnKxXk71oljt+YGeHdWTmCmRr8RcY
r3gPYTq1j3zL57yjFZQueuAWkdRKLEZkMIdazMmMHB6I8y831wMObSwjKK5ajkaF
nzp5BXws39pVhzKtFP1JvPJN1qcRv1/VfLtLPmG8vWZ275YU0gi9e7UoOy0U7/jx
Jhnvoqe1C6ejLOSPaN4YmZEPwf43wk64cQKnnPwaExtr1apRVyXh88yzIMcX4nZ2
FemzsRSXPWGo5LdCrSCgrc56P1WsrUpWE12iDcXXrAKzkwM30rnaU+ALLCE8cSfS
e7RoS9SZxV2uBPAGHIhdvb7YuD/OpTUrGb8/f0qaD5p6pmLFzI9iBn+Ciw6RNJuO
m7TPqfDnNW6DUGJ+SokxXBj5JPmvYcTr9ntR1AoQvx3/ye8nNm2elmJok691uvr1
BwA6dkptjZw1AzROKSBwhBbatBgINXyDEGbR0sc+f4ALjc0sPjEUljue41BQedRa
og+Yd9ltZqhw3h80MBH3XNS4Od1KINEjkvsYxhXVyHpIvH5grN4cv3kK3qOqA/Gm
t7dFvEFjhCEts5EcDvQroCv5RRc1yXXL/creQ3JdzlUp2N31W1WX9kwQwEhULbTw
ZuhRpwMKILFSR/kP8whk047irmYAechd5WkSz6z0CQMuPFGUwqCCGt0CxBCvK2aY
n2+GuCM5zdrtgR0B+mpHQ3IOk5V4rXvChjGDHh/i9xM5TWg/mMTfMkCwMY5Uctj6
+jtR8UBzhGiiOjd+vYvNV6JFmXOXW25PfladWepm/H525pNtqCqFzBqr63JWFqWT
eI+CqLWlFK+qQIUjQxzQ0ge/BBR4efd9bball7/LUCZ2gx7Vvi8dLTK0V6R6EBo8
iYTosjtIpZI5fW14EUl/VV+Dx/S/1gNLjihyK7ipFkOoYmP6B4pEPeWNnj8DiCzf
0JjnVQYgdDnDzxnjXJRN0D6I1+bYARY6MhCWuBkMaD0O0O431+97eHb3mdYMe+VF
F2eo+36Tb/+Q8tyi+lKaMJnRdYnFHbDEDceb24LLs4QxnYOYMqN2/S621eHS4goz
S6O3BsfcdbcsnukXjS9svWDYPueo8zMEcXCxWOYf0EqNzeYJWUZrBHCRHq2QDlW3
cME30/CPzL+iJsBaNPgtB4gNBJEG2KED03ElbGd9lmYyG2A+IBroei2P0VhlAQM3
P3f7lADn7ehljhj85fJNSm23C1vOA16CykRN7/3tX1JBn9zy5l01Ckbyfeybd6Sa
wiEGQZDtev+IcLmDRwmVaCDeYs1X/IpJVQ4luZexNuZL/D8DN2jqnMxzsn7aoy7Z
s4ZI+Wo9ybWFNZ+JW/tlV337jJlb7Ug2j4Ur4D18EslT8KtB6KD1nTQWdjv6HtK2
HbkdgluK3dk3gq3kYHGOw0vUwvMoxM5HLQqfevDyn0taoX7Rj8cOICRL521rXNkP
PGvLP+/ynBpEmkXsXLjlQNvb44iCrroAiaaufkq5rXxadXM1fLOOc2vQZfUUXpap
kCCW3zzr86j4lQ0nc/KRpOSKPy4RVp0++YwL7a/r8z2FFPpYDRhNhOJKWGMxPBMg
xRb97E0+xiK20ESeLER+nzYupxjHvGD/8IXB7IY3kiWuSv+tQcm2sEihLGeZYC95
2uQ4TvZZbKQ6yAjtzXO4RMFCcQHeaWWQqYgdHB/DHmpGx76JUV5hCcDeNVY5ZLp/
nGSZGBgYbNVsfLbyqngPDStaJ/v85BwIB7MfFjJ57GUyhQ0QWWxlXNMPEQcvXr6h
KRoDe4Y06YOkwTieCDasEp5R8uV6vwxbzdMR09tpaJonq8YuzVsMHWdo0VbHcJaq
mS8QOgQPIIN6brmM0M+e7Z3Eg2PdWIFYz5IVhpWqsWaZqB2EdzAVhaViQJj8cB4J
yYfY+kVH0n08J+C9K1i4wXiX4P5t8lGXPJZFk88MGC+uFYn3fKnDmvcnnJQCpLgK
xSeYwDca/lAIx57qetO3zYyTud92SwVUogN/xbCT8oZD2J5Ymx7/rMQrN/NzLsN9
7vMXF0A3BS/MuQ9t0eJah8HBALZBKlEfaY/YaEahKFMUEUmscBhSFt9/8zC0Lig2
4nrjgOCZ8RRljDMjw7n6Y4p+fb6MqlAgWWUbQjARp8tV+zKv+uwc7DCRIqe66yio
qK5ig++f0R3ujEoYHKSGcT0R/gwc8MmEtMwF7y/PY/+vIEa+FegowaRlUs0JeNYb
5dSfNX0r4cGVU/0yp1HIvsq5gRnNGDAKyXYrZiHQ6cXSNiP8WZzHsKoK6oyKv777
f0JaCMki7r64whk43a8Nbcu3Dr6gLEoXsrriRtZaPHor21BpsiGHl7w/cl+dW5D2
jTnx4cxioxcsfT/ZaIE0kroPHBTj3m+6C/FXY+n5XcnFT6WpR2jQ1nzUERtbaxdN
1r2ukYcTxItZC8XV/QiHIqlcrBc4gjecOG/NuxxX45h9RcDpL7QPI/YGVh792Yur
/9p5ka4OsB60TL/qMPMjbGWA7PpWHBVtL3wD+YodaHqrCiz49QZzOgd1YNa+zhzh
/Xp2hu5O5SnEwqSiy1UXQnFVbhTsLddjKeCMA1ZLKLAPNVQm6qgn4tnzvfYdmTqD
fHFwNXUO7OyFqR/aYKZkOCyplRCoYjrr7ibWZYB0dVikdFG4MXwmWQYLVuDwmRyC
PpDMQTPurKrZIe9mGOyi6HHuTRDtzb5bSfFu82lJZjaZbDbZLLhXv0zw92fkkV7f
fNU8bAwjAnFOCMYj24VlJiVPodcYAjmkjqO5OIbvcvIH2L9Rsl+Ejm/9CVB0ZYXG
hCf+/pK6BNCLKllK8lnk0uEl7GVAdrFgd820KBh2A1FAm8ArYDBgTw3jMQhDY6Ws
vctLq2QrQiCkgsUR4kIIvkWLJ9ybStFxMrNgUPJz9qrIpmDWyziIiIoONw8LIbc1
S40O4im/reSi5F1SiTlcvj1hfv8O6yFfA8zzdOIRkAHUiDzOd12lTjAMy7ellI13
E0Ad3sMeh4jMJg9hGcrUC/kB8zIeY04uzhx4xjnVvujT6sj0t7U95ioayPJRPhQM
qkk7oWwq3r9G9jtq6LLuWcQP34Dry/iVV56mVHxetr/UEHIfwYPbiJC0e9EP56WI
LpcsC7SMaTgRA0q19udmTGmT4DUN5mlyvE4Y9tQNS0I+JI8rsisT+OAc4VSiMgSi
zsuth1sQWneCv8LjOH8fZcAzMc3x9aZOsB8/n1mClODPqf0hWtPrVRVg5PVuLMR5
U6gZ+O7y7FauEHBMVY9S1y2fEdj+WhfAKQeZ9+W8J7Mei5oUaPeMeJtDhEYVZi5t
XN5Jez7jZRIxOds1nLfNgOxyEbsrxxe2oQOlRbCwpiQucCB02G3aWXEt2fAc6cA0
3DRgLy/9MHNCTjSunFLqjMD1zPjq4xsvadxy9b663Zod+2cl9vTiklktGWkvn9Tr
72wN75hwTPIxjBUnNHM44nUNubSPJOX5qvzjvfHeQzcsUixJ6rB4s9BxEteVSqZ5
YSVv519To/avMyoJuFlQ/mIGLCcAtBbeIjSIkYE0x9daUNjaytdbhJfWMMKeUB1q
mx53buGgburwvx/gMp9O/2b6sKrDbYLEN7W5QCZOHSxXSRbfgBzm7Lm03qj4cP9X
oQNUweKfQCU0yJmnEGuyNCCqdaPjXZn+pNFd2A0+s0QPk9tPKzdUjrMkZqGOSqTC
QSZWAitwqU1b19anAw38oXxB3zA6YH4FMfrzGyT+lYxv2PoNplAf3q9zEiNRS2h3
Up5NUhozAjj2vneWLKRuULj7V1Ec8gfiFkQ7px1BTFAaZfxN9kzDBMANEOhm6giP
7NKVmy1bWEfHsdxMEwah39BoS6DwdrpICYRYd5PBfOsJ8saIjCzA/RrOFx0nmH3D
tMkF/BN+nLQs/yKLQDTY4yRrgqtvUVL0pPSsz2oUxyKCsddsEQ9yKVsOQlWgvqnv
TauhHUyB4UUS5sNT8oaVAVfl1NGYjI8tzecyPYJmRLScYwf0b4ytOi6iaLNMVLnj
23P2cXKXySyJs4lhq+T0Gp6KQnfpenohcbtVoPDvbQJO3GH0sERbvlCVYjvt/cfF
cYFtyz0wGduUi/B6nVdLihtsVnPetzNiydWlfevR55/bRPl4J+1lc2mgczVBlGGp
bhP3dwK1/p27svJV/7J0aFET28VaU+fVOtneKMWH3n9GhOUpNXcK/ANCE3EuWZEG
5bnv3+YC5SqepWKaryV79sLEUE+ChVP0Qx1ZelnxDJhyKsU0UmBcyD2zBRfUDwrZ
/j81RWqtuVJwpkxiVkaJ6tXT16AFK5fZqIOaEcXIM0Q21MiZPKdstHDGVInWMVC3
Xrkmls1INYQCbm+TRNlKM8sbA+HCrwFdznvKw4zsJOCPNYq/fhhA2Efj+SeJshKq
Amm8QZsqHsO3thlGpa+ISH4YkGgZ2eCFjctQQnluHhos8q+w9Yj8ti6KdsaxhCZB
qSRPLleAIe7umdo4BJrMj7frwiUHhQE9IPebIMUK632ZjY6zvI0FVdPJ3J0iHmZR
ghJfFzRS2xWG3a2qft/rlpzODtng52adPgpgtgR4W4eg8NTAQ60+TLJajyjfMh0Z
ZH3/SGC1FJtY5Gs5qu322vtYTQNeYr90PwoOth3Ljy1ivGdJFn62cZNxHBnAkqr0
K1WWDLN0VBXP1YwRCeQM7zna2PetwTb50vKAgyCLuXy0gYJZcalwYCacnkbMrV2Y
0U4IT2Pun7/nRCre8sdYfaE5HtYiJ1j9J3fqT3oWAC4kmZEuDYTV1zDHlftafhbd
HqSnrO+3yv0UkNx/JNZcR5DuWnWgYIRU3rYQKn6mOLqSkWGO7h6CqvC5eT1y7iS4
+oe0bqfDp+agC4oPH0aN5NtrDZqOZuG4LOgKyj+dVNcg1exyhI4NZCEG4D2X46ur
2zU9tb1cZWlFRBkh/T2BIIE44MWX6mcHVJz7UXkLgFTFqgu6RPBTlFYWefPm7Nwr
5i3+kp2fVZ/zavLTrf6/VZz+N4bWDKBCOwiJsl0Wa18xHml38pl+nS889IJ9DMio
ZxLUKjbn43MoMxhzz+LzJtHqicLSVN/z5vUpHjQo+hkahkAjTnIoXhxVFVyL42kC
zAmqwmifIvq34l9uamB64XwHcVyf7tLyYqAqJprUSGo+fDudLr4JPm0lSxh5ToPP
fNG4wHjW9zi3neRfY0Un/xkQkDIOmHbq42T8BBMcUYrVZBpd686VmuZu2mrEqqrL
eajmuQDnkQpXytcWcCfLgOpl9LjlVdsdshNCZ+CR0AjJ1WbcX2a5n0FB8pku9si3
BUBHUthOomVHuBALechORlRNDZ+RT5nQZXiPFDpjFn9EtA3fMnWlI1yliAeKPN38
brDix6EVu5srCrYwN62S30NmSEUHGbt8kuNSmBtGiw/y7gvgnFyBRzb5V5cYYyJk
CX2Re2KxPvXVOupgQAmtNEcHhNno1sLA7HRLGhBX6X/cVFHlehefIPMVavDw8Sst
JthuspJnOYqeWDaEEd0wJoz4a60CIM/YU0I4O9EdCu78fifz306n7k9uS72CEwV2
UImplIfMFycpep1je8m/5yPnKGaFeRzezrLxxmnPry9Ii8ZzLk6o6p1Pd+ALkSdr
NRZTjcfz/IRCKavIpnX1ehhjb8evmzD8NhTj2hqH7jRyWVIclepehJenisUBotrv
IyE90Y9BB72WKRPo7ZlOJ5OPXejhjEONRqtEomIqZQZM3jkDLVtXrpFLmsxEqy7e
DyobsxKu8c8X+s6xlfnAP/Jpquw2U9chllJMPEXGFnaso47MIlykWHz1OCwHXRV8
u2aj/jLt6ib5lk7QhQb1QoBTC6QcYDp5dzIBnjXI0UtkCb5n+V5dVMlv/HXF/rYJ
QA7Qh9BXcd4W40lxdtbBab/bpAwIsLluy4Cl/oNhzGa7nFIPnnl7m1K3MmCuQFcI
YAnAnapAq51faBLazQgYPJZD11sxGxj4mcqSeh1xRD0Cf+/iLM2spcmkkH0fUIqu
q6tEbW1kAeBifqXJqZzEkElsvW7iLdR69TtI/juKbPlljMhyPIvAav3s2l8mzNAn
NRmXow4k/rd/PUH0kkI8DWBZETz4Emav95Uq36HzK01qDNgm/lzRqr2z8txeL3Jl
xr7JmGlh1LU4AaXbw6I8AhRFSw2iV/fu+XFUhQfheel83KEvZ1t0gg2TopND5o6C
U52zZ2MscPmetnwUevnOgP1dfaYFvwJ+tg3Mqkgjd57jPJY7t/AhH3GC/vm2qQPT
DftFe9JNaOg87SqzHjSAacznUMKepKxDT9MaXAMf8gOjXrEXtfazjBrhW/EksVvF
z4XXUdCfz7rRrJicdSMK6+kQn92J324N6i3gAF/kTpDWNymiKD8HNwQROYj4yWSZ
1Y5JZxN0QBz56wpPq62mUIDEplr9HZgwc47uxvf/hQp/7iUq0eDFw/EPNBwuOYgA
IJt0kBT7Pou+9b2snanULyYoUVTC7Zdu7YqTP1wg+QgyfC3n1T6NGunPqGSs08Zv
AjoUL0Ksqn4rCECMtlixfy2rm9gCiyT0t7Z+NvgRyZXZkq14TnNMccorHL4XhVq+
7cSPMs86l0gWiY5aaXcsAY4qGqtBAiQg7pQHe0VlykVy+2wgLq/g1s+BvlM/478Y
hwSlWMr23FtUXf3rNxHIl74ymX08KeDc0CB3tjiJLTXkfY1/7To0l1/ZE/IXaWNN
02I6i4raNuIda9MhRXjc1VRlaNKP5ERAy7H0oWVjXbxQCyKMiMKRmw/9sb96XcIZ
kfOVPby0miyGA4O5oUhKkh/pAxs7n1fpQtdUjKMPwKg8crpHhy+y74fwmHpaCUyZ
UF1gURoREmNdyX1wxvd/lISpohPwz7DRIcTZQ5t5HH28LFsIhoFshAA20+i9Eu8x
4BppR1YB5p6tpIilNSzyKcAVUCpSvHPHIWo1r7pj6oSBXioKyG6XRBycoK5Jiscg
Rjx7SGKRj+qxryOtBunlD7QUtWwU13GlPg5PLfdk8Mqo1oXDi/ai6fyiGQAEcTYK
U9ZE4qAi1iK3/L7xfF1OhHh+nJ3WRjtexswrsy+anRyLjwyqHsxx9F4TfJwfW1sL
BOraggRyJTgpcI7Xd9y8NyI+3/HtJdfHJFa0CRD2V06kTW2+Y3OonRH5Z8XsNDSX
6Aiv6ML5fVZ2sCW7aIBhxKDOqFSdslVsJv3ZSZ6kzQy3qYssMG4rV1GXbdlXwz+H
OHTSoQdxtQkmT3quXU8wTZG8vJJ/ygXaEM9Nk6j+7TPhkJ9UQH71VeyRMsLQzSwK
YwbU42Oedg1I9CDWQVXpZF5zZ+QvrsnkZGJsGCdXxTaXNcLhtoIEnXlAe3ubplLQ
hKP3JU3qwUkqN8T8n3FoyFEa3C9Y+RI5N1uQlSBqq+KjCHBBObNzM9VfhoumrULr
I8OXCoOG/aIHsGkejtHc0MT/E+hhsnKxbqi/kAqM35Q3qixS/ossZOZTCG2qYI+H
tXZlcBIT95RSWg3Kg1Np+tcNh0+9i8NMvTuhezZ/dPed2NN8I0nR/wcO5ehtDojr
8upcrw0yjF9mNFiSUfzYQQTbAKKrL7WDfwooNlT04gLpvoA5X8IJOrSHCeG1IMXJ
14rgxIg+xV8mwlCdY1z8vrJdSYBhJGVlzPPIr+ULsI8scT1ZaK0gvnyWPzKbM883
2r4hRv+B5X5Q4YE2YLnr7VhL4nWDKAlYa5zHmD9Mjri/ScQTuhrPuyHAgR+53l3u
xHd9FG0E3mfg53OSWHFu3hboOkZQyq8yGkRYZF0LIzAfe/GaxgABUCKGGra0Obr4
CJojByUihJ7cW3ILmp65nscY3n+96WtKbC63fTzGSAOXihuqhNujUT+4WEVszX8d
wWGZHL+IrEFqZYzxb+vVcwA2oydpzo3Bt7tWRWiuwb5mE7mrXz80onXo3pTEnKc2
Eys+lzUptAdK2nLv0d/vMd3SW183ojtThKMywI/W5aTrGHJZS1zGI7Gmt/D1OJSB
K0Mi/duOQYfquTCCQ2UEJw1JHO79sg+3Kt3uFzV/cyj71HHyFpg75C8/o07GTFYq
fD2dvx+Tf4TXrsVnVG/H3Y132kkL/Pck9a2uF90JXthHXXdDA7iGad1t1jaY/Qki
QNDuQ2sO7aaW5qojuUdXrr7+ZBoXNKVLLBAfq9lyqYcV7MGDifVBaXTuU+ieqNRg
Qvuc7/i6mPHhl/U2dsULLVTda9j+x0240beu9ZvRxNxdlwR/Up6hZq0BweftsjFo
3B2NF+kGQCik3fXznr7Ut3XsgTYWrXE+n/3lioWpOTBuk0wT04YTlFMqJlVMrj7Q
g6nhmiWBDa3JHJmqTx86586goQe7jRZhowrvsSkn/AJ4bxFa9GKaxGz1ElMkitCk
2P8rmTbxHjPDu7raxASKB3d3dh+yiGqjd4NQYas+PZ50KfUE2yrkxXDfMIcbERH3
jux+PmCEeOntGX4t8oy9v+HJFUi0/LdxOSdFX58fxzglgkquTumNATh87PNzzSmU
gHtflmjb98/fL74jqBv2pNNGmk8q2KI3gh9ltrpnLxVB7HSI8Dy5y8eEUsE722LJ
/qfVIUCwW3sbxSOs6caD8F6jzKLqrAK+FUVeVsq/zrOXRcfk7MoXo+19+aG//NoO
dr95ZwuvILqRGB7EANi15iDnONMVXMMOr7/7yS4gJw9BLFdGOoRKFvu+f9ETZuOP
dfkUkptpOzwRgBB+x890tjVJpZbg2HqvZcHd3+cbCPC6daujzA0MUKzcv6Dry1j1
kBQM0kc+NZbmtvZCa5EpmC6IUFazjkywu4B1Tx+Clb3vnPW770EuhTSUMoKseiOS
TX33CKSUXFcO+SKM11npWLrSgV8aJRyqsZiU2jnVDl2dCn3akKteCxLUlESef9Sl
izoMgar9KgAsNQ6iumOzYzXNau40bU6h510CuohU/3Y/qHhY3FMg6GVwxNx/VZcN
PihxkMEc/u3jCC43HFzHsICqFdclPld/1BaeOJbPSaGtxaQH8VeAS5X8fUAxsViL
EWVypjpxTtXKYCvNKvc2Jjx632BI4SYGWIVfYOB136gCdiEqdLSrxpYv50dkdSM8
iiYR5P9Th/QDzL6jlLes5Ks5L7VrKdIMvO9kfmyjipG5zddJh1r5cecxu3MK+z/l
7kFceusszVbbxWowwDuOgITaU2dmiKTC46FKxlurcDA7YyC3RLWSDC5c5UEz3iew
e9ON3Y068w7ro0M+LGO/48CCx3NjzZCFQcVired3P7x/Vsem17+3XN1sbgjmxR8X
u3mO14skTkTrRRuAS1cwikJaEginoZAucu+S/U9t8ynaPAaBSwKcR1/qV8UkXdvk
NNHDsytuG6KTfn5SgHIW+vmdk8PMa+lvR4/AWQuGeMg3sSmyrv8Vq8imyUYuMIXs
eYLm2vzb3lJ++xFdN+oofSq0OIPp/JcRv3mPW1H9tbhYYTA3RfEmD749hzeEcIqD
bU89gzINxaNKMrxEe0h5dU+zox0fxqRwfwm4bbNZkuTdkKyoYcVmZi20kgE8EX5F
kDhN9heRoE/5hfmbhPm9XuyYhGqGYN+1dH1cqZdw+M9q9ndo3Vj9d73MDGI+wy6F
dSiqFQbzQISL3SYLm2TPtVzx/nQ6C3oUQYu/6zZWJvcYoB0pweJfUgXmmmhp6pQX
VIZtZ1eSLfttBJvJwyWt0ctW+HhCbxmTSBCvsJl0ziIclgAnMMceRLYqgnBtZmsu
9fPy+qOo/GnOwtsHOWPFamT0AWb/dMG5Yipa2rVE8+9yQMQXxLvn24tUDa1/X+FB
XpNct33fauLPvlbGho2Aa2+xSms8Bs7G27/ds4vQZo+zH3Egf3XmjUMaVGUHvkBu
dM2R4PQeN3lMCf/Q/SSFORZ7YpkSeEZMVLr8qnfSXmlSjc+O1fBsl9GQLVz4Q486
qA3Hz6BOCqyOkcVB4+sws4Gx3DF1VdjEyS4h434yqvjv5dmjgj0tahbP6D9c7KYr
68zIsslH6O1GlE6acTPT5BhhwwL2l506w6/ydoiJIx6afu/1aFCraL5cbl73M1HU
4PZ6q8SxlmVR8Qf1WR4yN98qT8Ukn7L54oKgnOyrVIp84Zb7uCASu1h3hxM7KvS+
AwG0orHhZRfxePYkl3qIn3gg6E6ZY0izjXtmI7BkFzbzkJvQ4bnvWnNO1ZRR6/pf
Xfadt8S+Hd9693tP7avSxc7LISD0NvqBM4CdyNY7zL/i5CvHuWjGbbNGEJxfKZRk
PRUi7Qbd7t/xlywt9gTlUPgl/oW6h/SQ87Ii9KCi7Czg0jF2zZmzFzUXXT6gEruN
8DcyRw5bI731wV6R7SvSnqKgv5pmDAxs/PAxf9ycqv/QawNwuiZ9x9xcQUOIlzvs
i+V0+cN8Chqv08B7WDWHWowjy5dL1yuwnKI7ip65DTvKwV23LhbOmjqdVVaZaGxr
1UA0i8aLfMdiz68Gs5QXbrjPx6KqGz3wlTNe08ubiFE0O70kZ2e0Whedvnip5Eqt
bUIJ4mfpJdhBkvOjDkrcTKodjheDzhfQKHdymtYd6uc6jUviZEY3yhbBtleWJtKS
gzemHGncqiy3j42szDNBr0nOBzFMg7p2UBqbQ3LZ3xOuydG4lKsfzdNwBJebilcD
dhUpNJ2u987iFBLZNxw2euw0fDD1pWlOmCqbwnZCSmxydVHFU18EK60AQTE0SPEf
i6qHWvHOi89AnN74IyUFcvr4D1bVC6UGS8c+25GoRN7wBgr5zfwNkKA0/Ba/tGPb
XeiAXPVaqDZRqiKt+wqoyVaMJvwN4caq1KBZwbQZIUQNyemXvLNeJvZorLo4tM6U
jDMdJqZqUj3fd5lMDro9HEKrwL7D7LNCnNhQAiobNe4otYcGHwJrXy/oL98vK9MR
fvowkEcQVTR1E4C9sjS26ABUbNlMGc4D6H321RKevwKZvDPe+151IMS/gB1TDldz
C79paUG8tRQUMpMoRISLnswWTKftHuqKjfzscvt+JtKSCf067BicLcqj/niGkFTJ
NdUhLZqtAaV8PRfKZkMSG5QaXzND5iRvVx342Y9TIML2sJkT29oV7Cu+qA3MRB7L
wDRekMPJ9PnR+DUoUfCJhOBEbbPqRgED8GB4zGiLB8MSnSgJD4fuR5G0RzqyKC0F
UTA8yufJBkbE9oR6NrzCgwnMeEw1ZA79h22k3N8BvFygtbNrvHN5FXM5g1Qqr/kf
idO7ROTYFdK8tc8XMtvaRtJILS/1T7smYEsVYJmXOEfqa/SriXe4Yv84tWKsByr4
+M83dHyq3R1rD/s6UEP2aPHaJ00aalKek1PmIAWOPTkRnqW5awuYQvFVdavaLzF+
6Oxkrhl8kIbGthusUefA1baJF6xOrC3/mUyLofocXoyIxPJtnAM/MnFv5uABV4/Q
mvqKkfEvDtce6G/P1dsbdJ19yuaxtjhuI/OEcZxvuFM4tXoPNfgdzCJLDTwrw6vx
uwRCNzkvQyZUWtZlW5tCxJEngvPYL5iMeOCWKGrzgpcnPphAnSX2w7SAAF7VSFhb
kUishPQxRw5FIuTS3oj8qUwfCxzwBCOcG6j19TVvgz4pd0uu73/+B8Zoda6EdcTF
j49PJw/K9341LP/ny+QJsBa3SqOWMle3tZMEpMBFum8oJF1qB03jP3tNwfGDo4ys
X05xMAxQYzdapNtAw7ylBbRcEx+2t9Gsz7JQ/pp00sdxPBAm5aJp6DCvLHTYLh6C
cZni8XxBHIKMQ9YvAaEzdjWtg2hCHyRTH8Q76b21hvI1H6nMJDqld8jMlmlpESBC
j658W5cOIQNdXlJCKhWUuDy5XuhfjleGaHC+I+f+fLmZByf1IgezlHlXEuO7kTl4
HGrNdOzZKGQjcThwkx/Y0iFZUnIMNvsypiT/o2qEFwQJ2CSmAUjSnk8neeA/0lfl
YmUcwBuVTA+PbHgVmyH0UMqxMVFxrJ5juEkE4aVZxzv1kZfoE9Uw/m2iSHTMeXtV
QWoxA07k1lAKzIieW1tX5q5SSULvsL+FBQbQOCQ9Y/PhYCuBp8rE6MxpRzR8387c
JG+4i45uAmNSHfaSmIdBPzAlh3BBnvaMFwPJWBkGZuKRIjKtQqwjEa3omX3gev9A
lGBBv6sVmoH5pw1CvxitrvB1G5ZUtSWijMLk7XWBSGGVPrBeEUWT3XIn+EPvKmiX
HV3iIgsrc8sNnqowFCQbR/F3VpjYdAdUIbWh9SENOmkB9G8BgtuwkqgiaihAQkIW
l6poEdpOXdOQ22StWdwqhgz63OsQbx3SJhAJoOEzneDs8QWiSxsDUCyptEJRNA7I
1gBYxU8HFV7HtDFX1yX2FWehKjrP6RaLuEyibr0pN6eJhOQjDxdPOEqRdM9PUhRf
Z4wqj2XRhE7gLQrlND1pi3VXeOwB3RpMtV/2T8z/HJsM1arxTpxWtdE/PkeDD11M
ccirSV9z+9VoLfb8j5LVwv/ZhSwFr++epTXqijEyfZjbyWhNEwQnnRy7C8I7h36A
1Su/w59zeyI3yw3/11NKvL4qiT2Ri+2ViRZeIkPSbVht7TWOlhVAK1In5m97cnCQ
5ECoKzvjwNEKhINWGWL9Dq0h/YWSt7mzXiYFkAQJxDOaBABZgpbUQtv60JhxRcre
TcmldyohVSz0j5n6xvPsml9JdgHTcug2tDWU03VmThUOnzMlKkI17Cily4FNTBwp
cyGG6vDk0606yh250y48eMQvYW98wSTh/MO2GlajiRnL5i2MrISDQ3SDR59X4VyL
snC7Koxaf8nWGXRqUYDRgCxLlU+AUaM9iGBRYL0bpWNmcI70BI9QNMHqAbGlYumm
zNl+NNXDyMqU7zo2HAuTEuoTyy9Lbf+YL6mym6pIvJRusDoX5aLCSzTq93eBKiDt
7kS1bolp82GYLxcV2oZfoNQ7W13BbqYMinkASHzM5zxqvQL3H/bZ2DkUGDdGqzws
afwar/VUS7nVNxwOdcnPXPv+cLpHL4cxdrVSigDnVZOjMJbOnS6Q4yJ4AKoE6SRz
BzmY0PBMlhaPRCo6Z63JB8++nVwobKfzV6APiNHC9JI+viAjEdCrF95pGMtUCxTI
9/UVxxeVDjI+8O22e7TOinAknhHSSRTQnP0EhTFgpawFbIDEdlGeBp5nfhTXZT0l
th9SsApLwRfpZ5AVghUIE3Q+vw4t9rL4ASb+wwMkNZ5bH9+q9zbPAcGziSKSYvBE
t0sXkoaVaBVc7l4qBH7bnMyXfvMIyfrohgw3cjupniHpROvtE7idpzTrVn6vWFbV
T0AtXdTuVIyYWPMEiz4yYOFoT+l1gawEBSp369XAqZudmn1/k7qVTF08kf4e5OII
OgsykCVmdzNd34RSL6dVI6WH3NJvYaHBG4AetC0Uz6V42/3BYKSzTzEt3kp2XfR+
dExd42bnK0nWryLObauav8l0+Zve8ghcPmcWzW4yW1/8Wv/c9VI+gOJ0fARI2cur
gEwVSDcaUkXwljmE1/uSRMbHzbfQvS/z8pVot7/BhTKfaZtBYnEr+cfWNyu8g/bK
yZbiPDjk/jv3U6ZJ1PpDHTkutpRBDGnoq+4KtysKn9A=
`pragma protect end_protected
