// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:08 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tcuFwuwS+s7EKE+UyZUlAsciL4ON9ghcAjUrKcTdrFneF/1aBnM+g68q4yG45mFG
qaMdl+VJYr0i7o3wzFv8pmlmpbibwaSx3oLZfe7CVOtjCBNbwgtx89Fs5xGEexYz
jnWM8ExeZIQegPU4wRoHOxVy2MRZGIAFQ0u/Al6ypRI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9840)
zxFLjFIx1nHfA8ontf80qWEhKI/ZG1MQhx6gypuGxtHDBGG621qb1zuSwbJAbNvF
8Sth+tGynpQu9CVPHOJEgVOI8G1jqUrc55khl/YL9aPuKTCzqEnsM3a1m38wPTmy
l67RYeh+TM62gix0e5ujw41MtBIfO4ie7QRMjaWISsXfCL/OlWPEXvNt/V0F1FEL
XSsg9qYc+g2WS42Ky2hXKe4LVt21iR0ayjkNb3qV1bU1Ow6gSSLkJe182fHX3EEx
TGz7xiZ8SEt8gMCWHBOuMFyXeq6fJFqxx0xeojhM6hOGiTnR2nETkwK9JZ7+ZvWa
LgdHFwHlHVluq0ZY1FfOXfI7OYXhDMFAfpswiItXlQy5ainUctNunVACwjLFc2N9
o0RDmxlETunoyCH5rs4KukdqEmwK2dUyZNslAqNPBDckOOc4MxDLTothkLEO1lI/
3vkfnA8Hsiz8kVyvfZ7gPXvZQv9ZwET+LeuM1nuLyRf9exjxcTs3bxNhBgRNyRph
5dAcyMNfnwNkMOmxqcrKr/m/U2veRFHpxJNSm01Kythrv77XV2vc11dPHXnnQPqg
p1jxQHsq4cMN3PnGJs0o/cnHvFVPzIcvqPw1Uqh2/LxJD5C150F6X2jvtwGZoebr
vCaMSkwpok4+LcwxW6GcwkLJuyPEKxiU7ULqa8dz8l31Maypd9UxGPeizMKXcJng
dhQHwCK2L55xo6Yf5IMUxkZtn2vy2HfksrFs88VbNKtI1ZqtRNXJfvSbqnsQdleF
wMtK1reQQAM/gfQebYMCvlC6jXFZMsP5OY/8qrJnUER729DSmyxGgskhkKX+zvK5
1o9MjiY4zzqHRrLLvAMv3DcIj33RJC7HeG63aXpsUmuJ4+Z8Hk7E4St5S86RXDtE
TlqkUYvq/yca/lXoxmWd3Cn+l45lRoeqwTkqCfbXle8KZ3A+3DHrbjX1+i6LnP2r
kvSH3KES2viuwnI2tD1KWkcpUfxDUARo3Exvhk4kB/nZsp5iUXMZn/3tvsJru9iB
tE2fP3lBZ7Og40d6BeyOzIfZqT3DNJG0DTko8xDFOB/RBs3fmMr4Nurq+9wM1pQr
Em4819RrmUU1jmNAP6eYJTLttJgbFUiOWjk8lcf53L405ql4UhX0RABSQHuv0eeX
PYSzX9LBV3ZjZ1g/GU5uAXTCIZ16nsy8UZLiXzA6J3I7ZebJMHpnhS5Oe8wYgDsL
eGeFyZypZj5tyiuZQuk958wvibs9Utmk2kq+K+wkWCkTh5Ona5iI+hdji6XyBFm8
E7YQt4B8BSAKMHErrg1lUmIYnJqP5vjtxqGWOBtbNNVPDoNfWtnb5HJaxn2V3HX0
cY7oJvab4rjpACE8hggxB1oFEGzGY1xt43lrldYm2md45qss8xgpc/gp8wubsMLN
PmpVmbXdR4YUoWvekKk4gNKd09IeEs0jKwBvDTL19aoQ+IT/TXWE+pRuT883K9hc
Rfj8YOv3igoxcDfx/ZNzVfZxTA5AFJ1JBBCyoSPhh5DV2HTAfEz4UkkeeeHoPSnB
tKcG5LVJrZl8VLu/bY/qEgflJlC4tRvedhSFWC+26j13c6G+/IzOPeZrqzeV+t6T
8dJ3EBXWpnqJBhsex6yG8shMSFq0lNbmoq/FgCs7boxEIO9O2BAYFpeM7V3DaCRn
UyXzJgYGBuTbW7wB+2Xzj1415CVIHvn1UjyuAKe9dY9F051cp5S7r7YPci0c+5Ao
TcLqqidI/4nDbi7wwGcGimJlN2pjE2GwO20ItosOq3tXXsBSC5demsNCqrz0SAzc
XCYHXKPeIQosBH4V/w4dxr9EbkviQawysvBMctGnrowF7XGgQOda5g53dTAWQQhN
eACKkopH3lbhFt6IUH16uuOJ19Rw+kdpOzNWQIAi/VhdZh9yOhHWwmId1hqVurFK
zaKwvkTQ4R7lTsSpQxjH5fpk+iNeyxbfIcna+/S5RkFPHA6C1njnGWgTqo3PewjO
fE4/b1Jqh/5ZGeCRhvyqqYXb0b9ODS09hrTb9wFQEf4BmCDAup8H3hR9mGFJ8tIA
yvEYwRt6T5dTQEqPHAIhc3Votm2Wj5HOLtWpAQHWPZNP95Tx/xKqFh0C/UfA8QZ5
K7L6MhncllmUZyVTN+L1UfhRqA7kKjmiOl6osJaYvIAoGKzfvenAtF5/0CwTeqau
ti4ko9iElMRV9woAfbfHNsl2o+p8vHldkKCOZep2to9flZuGwBO0q1dA+2Kg3eAV
o4JFkxsknEpXI26pQGXjKehWee75NoIcV90CMRAEg9EU9YsaCQD9ekYC2ZtG1W8s
JXpn/lwDub1TGskYFiZM/0VLvOzXKCGdfg0J+zJO/9SSp9U9WyNMHG83FIL/AXhp
mZYSoyVwaUofweBPRDFoDWqpXeQaPbvxoV+ILC4NLS1xvtazJ6IU9LMyXRRPh1re
6KAeTJDP4ZAI/fMQ8mkcwgAXFYiQ6FPeaX1xO0R1Fth8yaeYlnG8MbzGIi+nYvPj
rpOhaevZhbdc2tHuunLotx6iNz5/bWV6ILyVrnAEyPNeFyU8sApToxjBlPK5J3W2
InDxhSNizU39sOJfsb2+IG+RKKc7XTK3IHOSiw9jRCNwq0sW+BjBg2kT+ebKyF/N
CIob3ogAmHiDKAvg9UxGOUZ1HIXPRgPLDfOk1UbLLgP3w79nhNIty6P3bWxuKLew
v0H0BcP7ltGMkp2BhcN5gZJKfYPMvcmFgZqUAroNqu4iHFg94RKRn+9y3RdGwJjg
hP1b1mwis6dtfsgaKYaGt/Q3l1DmadoGYceFoKB1RV2IiPsHGn85nmvIPVEqrKoY
GorvU7pz2cc2QQzCNzzHG3K1TG7rooBm3U6XsY/FtWbtjxX9RJyuB/OewspMMxJm
IlDy944RVXhL5jW+JwzyS3Qjqag0rw7NxMaSD7eFiJ2EAKWU7KCKzXKbUMf2hZ7Z
WlDx28r+uRfmMcRCpllh0VLHiywYsfPt0jTA6e8HS0Y+4JsAUwimrMyDAEblBxH8
kp13r2oTgdKj2UYSlzP6Wrq4J7oKPiJgYDS+uET1sTR2hoLRt3LxInco+1cwexMm
v5FopFzKoQALWPQxsiyvJkh5tVojLobYzlBS0TJIA9gj9Au9PJbAzSI7XSf2htNr
du/73ObJmGI0k1uyayz83e4xMjMm4zbgIoI1pRA7yuQ022P/dl+BPhDRvbYoaiBZ
g1uyLBAxbftg12G3TOE4KR8jpcL5jEVzUsPH+ow3txwPmawS6/voh4cgyul8O7bW
DS1LIE95tqbzr6ULFojQgD/TleUZiGjGuWh25qSj4oezyv243v10FbosJ6HjBfO/
1bCbTkz5ytJv2vNWSow+i9WUWz7uMXXTLMkZvMpWFJqzKRn3Z5B0HABVIh0yQKj1
0viqe5+XG9CU09LNzmiU+N7OgrJN5rNu6W/rRmmhKrMXmkcakfFoNwi/WP6sl1B7
4w/oSwvpW0eHQ7OLyBSO1UhOggWTyTa+H7WlthI07aEcfHF0kPMN0JwBeJcu857X
Yy6DwTdYZf3xAN6IInkSjIh0j7DPaK56ps95bh442a0qOVCT5E/KxbYZQBRHZ6No
3pms6lQlZcXVi0OIle4GHtZERebCT5ScCgEbHJiCq7aCMmayVmVbopjyFo9NyagB
B6jjXL94ndQCNsQWUOj7LmhsLuOhpNix65lypsawrnWHUYBZL8+qEYkRXXheCzAt
dUqYgAdJpK+KQxRVrh27amtydo2YY/7dKrWP+JZfBbdyiyv/f+ocGg5b2HVxVQEp
aonjKxHTp/8MeYqCSIcGHL7IfzKctJKUae0BqANoPZXWhZh1lZ3tvd4qLkV2S3eR
+Vt9aTjX8rC+MUEzwo0BULdd347nwFyONe/GVJSWoDbgJkmhBr7n/dMcuIv/f9Fn
4F7FbhCU92aR5nO83LmKxZv2NvnJ4HOzT5DLvCYkj+bpPsy3Gv0IkkwGRtehQPCD
w/kSlhC3n3YTKb7OYWrP1HnkmHbDsVGytUPyaDfAESOerIxBm4umaa1HBJOB9X2D
cHarvUmF8xOfs9hx4FgGSSl5I8I6y+s3qnyb1kdPd7QRA8iox/u4JOwtyAMaMTIY
2cRX4/RD5srAj76Gj3F2qM3SzRct9iB/ydzRqFDb5H3uYsZEFqH5mcsUdcykj+/B
0mNgQ8D0Z275ipOM3IDJUSl7BmjFF7GO6L0h/JMzGKae6rHgjpdFg07G1IZbEUhd
b92CUG21FPBvCSWBRNxs/iU8mke4EgD0StetUm56DMRBIT/sT4L4ianqTt5y3XYU
1nxtGccmd8oxGIgMVMXJg1jZIyPQGcpiE2m/4jpRK9Ys9nXdkhPui669vrZm+K1j
tis9LLcoqtwLe4NfWnIUzi13o9Ku74Q2p0sq925W7I8aiIHUVwyl4VDcShxKq3IR
6lGgQXg+Q6yOne3UqCP9RZUQEMMUY4ZhMKGFQuZJfNrZPr28GKBh+g6eOSdpf9+m
RJ24hVCLMiJMiCAgl5jbOUpdcofib151jzCk6xfQYvcuFix8xRu4h6D4chMlCyLI
kesfib4smnr54bC/PYVldLwkz0/jKm2BKUOBBrSR3LBwKnXFVmHOYgg7tb+Xkaca
SIGJYt+7z0CoAIBKEGE+RY4zIFop5+lvK/925IizJfq1FIAGqz5sEuqARQOFM+vC
OWLIYxjgg2hS//eRCQawjmEMaTcH6StETPLfO9m8StDcC/TNJr9UKyci+n+kcAFP
z8wTR23PQ4VmPfMw4gXfDkqVlZgYROpyxapVxT4gkj8D3j669CTv9RMXmgLYKJSJ
xRqP4Fuv0PfXGPPGdMR5EeFUosUztKqWnTWOS0UrQxlI+8li9goq7X8t26wymGUy
84kjOvetWmlVYCKnB/mL8qgxi+Y9Nq5thS5GSDFRXE3bCCFR1ImyoqzIE4swXrVv
aEOF7rk84+5hYMaBJs7cQ+Zht45rm98OQFZX9/IC48wtOyvdAOlFmBXN0pDCmYqA
kfjzhapCOymoeZ3UTXnc1aSpT0MV+ZiR0TNI0r7eXKkoS/vBswQ/2svKUg9dbI6l
uQdsX6CJKGUuDuIHWaW/UwLDogE7JVNyNm9CwE1rNpZd0hfbPq4w4d0c3SZ5wYiD
GpmDIXRHwb6N+G4K7XUXMCYpE/mVX8xgC9zKvbQEJhJGBL/HVZ6fHyQ5HjWpWKyD
OpRTgiMjmqW86KHCWIoOXVs/7qc/s0pxYtTXHrKZ3JxDLoy4+7HpVpxtorBp4dTs
OakKtt8hWGtYU2+UzNz3WKgccPiB+FnPByhnQQ86K2baeczPDVUT1N0kA0IAh0fV
BUNu8T5d8/4ZdjExidWm55WDAd+l0CEvF1Xz/5SRbs9o3ojI6i1DqQ7t/CQhNFh1
c5rocpgDxc2q2la3hxSNP+edmYgALli57aRN+pBnI+yE/1VQLbhxqS8+wyURiA2v
z9buQVOTIGGa35sgK8x/EI8dacwqm1LmXuMRdduW0JjqVN1Gq5O7FHAvRKy9RQnh
HZxlrY3cBwViUSDnN8tKtlb2lq7fy7FEcMp32KRXLz/Wx5KvtpNUI3m/IwrDtJDD
6YHa1uF5PWNB0eQoBE07BiC1aZAMb+T0kAGTwGJzS+eZsbBuXKR70idpDoD3mWWx
qCp7zLh4GWd3+/wgjVe2A1PkRqr2mXB9iD64lYWRd+YmrvyE0+OAEJYo3CcU1r2K
9U7RepMkHmvgiCWYT2f7xpASDfh2bdLnrxdfk/L4tLmZI50l+NN/tMojVCe+LyX0
t/CManM5vN42/1+1RzufvjaBZuD3pbTV+8EknoIGKAuierKT1FGxnNSTSU7jLluw
AlT9rj5EnUefIm+kueA8tY5avRL59vdthi4uV5Tufq1ikwiCndHgYOnRaDpUGkCq
sd7LQrrEao0kYbCpOT7RVRpDAuvSHy/XbXLV6PQMqPAb31HGGDFshlm/AZWINLYX
yfxClRQGRZ7aggihUaR1IU3ZpyEAl+ZcB/mN1JhiCbrOgehW6tz0VBAKKpTRSA3Q
NC6aVZIuSBwtQNSPAJJbRxXiurstpTfqDbyZwLkl96eqVRxlru//9KY9PRfnadP2
udbjbcM/Z1pPAplf4RIPbl13N84D0A5arAV1OqYpuY2NZEfBy8ziFp2Cx8KZLUR/
zBD9dCLvMiRWZKzytzwZLu31RZp75Fd/dLY7JRhREUzh+1XufMVaU3GE+LHnciro
DWarUno8W5FasFyZSdeO2m9rMdrsYXDquxPF5VI+WzPtRThcwRJQPOrBJgjwODiA
5uWZskCIlD3Aq+T6qM/JTtk+XKcRVQ1iUtlXsP65V+IsZ1e61XoVxx2PnUHOTye+
RIrWCQFtDBAd9BNgB8aVvv7NXXwDzFBA/qM+GJZt1AiC2TtksM75bRMgviiZ3WwU
IEoldLOVaPKClzCdE61HnyvbGMbfjKQVjlptTxJvJNC9+sPDMZf6jk2aYdpz3m4s
rMrIu1DQ+U5H4ib261nx8ZKMJVi03YLUhQtcMmPnDfuWIf7mVUS9JxjObJJO0WqL
0M7OYfgJr/NKLVbiOiCFoV6DuhS8EAPA8egmzfgbyzXiRPnKKT6dNheOT0PiMwhv
t0VRkaXSAz9ChuukegikiK7hGWuPkY73AUCy0XnkD6+Sx2mXJoqUsWmPlUpBnN/w
TuXxF0m6LZ+ougL55px9HuenaChygrsjB7SBmvI1P0AugK72IOjiN8MtUyK6qZgh
3E61LmPJ62OX1yPJ6BcUtFHwid2ZbcqfeHm1nP9wGp6HqHbD/ZsbkTfYFU9vHf3D
085uE6E7BR7egnXZ9DBHMKE8MZH9QyLvC2Gh3suUWyiB/YVnwaZcfGax0zzeD5sH
vKqxgi4YzrD1f2cxL87eHYsKvNR87+cKV9K2wOPWl+WhgH0Bbc1Fg4ILMdtri9sf
xzjBWpuiMyM+zCpczloknu1vHK/UYj9KEuia5hWu+pXwcx5bxDcgCO8FZ01LKSUK
vvlKGrEzg4HOFD+H+tWBDg1yJWFawBigrG5kZo142dUY3QmkRYrTSLi54nL5eOhQ
cO2EJ/9Gb7kTQOCqopmp+I8/a5ma2Tkx2471YRPMv6tNSgWhYaP5uimHPIl2vv7H
KjGqlRipnuDtmqqwJETwRhtNmULigAQXUsxA7j1W5o0GGQ3KmMIOgGIdw15gOfsH
LbKHQacdGQlhyYN9t6PkBBLWnD4KgixUPUIoDRo9tbDPjChTUmjQzxAKEzRJQB2e
AMcuIWjXj9Lr24wjznTw2iHYN4PzdyERMDdND3hweapZGHbW88gfCHW4Fs/BFdiF
dEQbv6yK3avOEvvzYu81ivXRuyeiUbwxZ2ASLiHOPUPmkaegNEDHstufd11AgKqO
N0wjkw19IhWAKOzMyVMjyBByKBsm94sF8i/wLobSANh3A9YaRxDdUqaFjPxMEOkf
c4yUld9QwpJFLeXseVV5VF8yuvFp6juwDWP6tAj7iAOAHFwy5hB2JxGp4Aeh4y1D
KGsEcZ+oQeM6/XvSuOTh7PT/cHIYqF44p2UesG9usFMTt5WQHKWin2iXXKslVMax
huwug7gBy1TsFY/kDtyDg3+il99cHWW/00oURNaNQAxn0kcLGBr0bUl6PencqJ4c
iTC3qg14DtiB2DkbUg9AmPbtrcTLVUqELliDh+cH5+MD605SiB9Frd5xzxNxMBAJ
f4D6R41z34Zs15/8wGbtyUpLK4bRFDDOY69LSf/86hDW4T3hgSI8T318gx3w0msR
DTn4VNiYBmAmtjcKAA233hmku5fHehnQPIg25zOXjCqkkpO6ml6qjQFmVK8fATLW
v+lQlMqtTqZYoiZLHnEfi5pwYE2eqJ705a/f+o5szb8AAjf40Kwh3EeVATOX+gML
U7hM0DoxPETwvmZlAUisSEZycBAmOWBel3QDR/aHZEwRyAT5Q3FG2cRwl8TsPXro
N4x2MSFEtANk3YZHUJIw61DUG/cUbRKTVjQgsr8CMfwJ4BDMLSx8qLEM4rr4Wzz1
HllSsDFZfTM6EewA28D6/uXZH76Wo11xiiDnuxaId6AK+HBhPOqjiP7JQ6yjCwVL
tlJDYeReOSTdugsNll17Q/mmou11F5+eQnf01MfbU5dtIbZpH+JUaKKZWwEO0R97
kIiZg68GpX5HXbAdiKkSU2Ux3hp+JLWKo2s6IcXd7QPp433h8LVr6LTjEZ/qoVm9
v/l4tY9dxgLb7LLOU7TKggg4hRyiSzThee1/r7mEyyZIg9dB0yTpRMF0QQLJgnAO
JvXoDHuoyld1SvllLdpY9wGPjD6CoA24vCHkaWjbKCfle/MG0g9bxCeKkSiESdSv
twT0gfbn0aHV2JtL1Rir+wL94IP+sFR/Mls6vdptV0J7QLHvzMQzDgfgKF7kiiGc
OD0Pej7s7Y8OBRrNq32Ppz8qqRrC+MLRfYs1cp/8jmW+SkykcEh2vPK/b/vzjGAb
dcCnf8HeR+FRMtN3Aa52zFzljj4SbmvJOo91NFXD97ICck8umcoHutLAtzgzzRL3
CivSV3dKpFmKY5IZHrpP/zzxSdlRGRydZpxChquYF5Rr3VdfpKk3Q9ImX5kY2mdn
TTOuu17gUnhmWRM+rMvPs+Y6lvBaKpeMuf1awc2XU55Dzlb76hDgqm3zLlgsjTzu
nF0aHLRYdAJUP5MdSL/fBWXh/2ug0hFxghEfZ1ShqsskX+xRiPgka9Et5zMNliiG
166nugb+j5yHuBz5Kd0yShhmhTdfjUNZq0w/OTYciUvvnZisEKJDP+ECQj529jhs
n5eeu8wUPVNPU7qWAajALPB6wSl61Tna49+JVuR9ER2hWwPvejrVwTM8ZrJpQ9rp
ZJeNMXxAv/G+gBkm61jmybCk+24PSTCG0bJiuH3ezrDY3GDlRmwNMNrFItOU9+0N
ouweDWUYN67lnQOtY75us4hWJkeCcoJ1lgGZ4m7EeYvVzfRYEjJK8/nuQElwBTM1
lN5INRqjP7BwgvOaCQTtNNCOpPkEwJ29qIpsqssmFeJrgswSSq+1KMo58pOZXnnS
bsyRuOW7TTQYHdWiULIALtY9VMq1irodBtgn+01Ty+FnO9NWQmuf2jb4KQANLaWQ
/fMqZjWxDnki9AgU2Zr6WOsjrfsyhoYiNqpQ8v6u9S4Qb993Ph4wwL33N4e3DVYv
HCF1hYjC5+pdCnz5Cq+ufXB46+NGv+TAB7V3RlBF4NcDtJT21aCERK1s7gw/6XCm
tQ4pw9o3l9OK/auUsjq3mfCZ94YyG4DVPT6h4wGNSolyeUWm/2ZkKagjjzxraAai
JBPaleEW6xo0cKoaOX0QJNY1Yf+/bIgD0201hhWaNDud5T6H7mHqM+cNpFXRhNZ0
IxEWkmiSvEPP2AwcokpRjQ6K6x7eoOjhBOtFeWlZm57LJTUBHoTB9GJfgNtid9ea
TWlxW6YEbxOJvHpRTlTt0Rnz4ZpAGZL76ITstTs8C97MAKX/Nr0dV/bgwGBnI/Eg
q+R8I+th9cEhEiJcgP96+mIj3vIUtamm1rTQOu2EjixxeRAdWWW3cE26pC744JA5
4IkGuZ1D781b2r205btfV0wuYm2j7C1uC3RjGzaRaK8hNW7aCyzPHIUje81kZ0+p
JjMsupj61M5og9gRCS6bgwnl2xlgPSqcMo/18QSjWpNBwnAOJyZklcO4Age6II3g
7MOoG+ZbtcCFRb5Xw0CaApJA3RuXm4XkotGHVqIhiTsZd81pz8DM9L2LehuGhhoq
p9iIsTuWLX2Tn8lKjrP2/wPJ/V/Woir169cZtu5rTZdSftRY9ji1mh/YtQ/Z9SQl
Y8umyESh9Ky9NuFxMkFGTBefp2gvbxjL3YwvTCW3NGn94TxssIIax+1DrbmGJxfL
xheOceh/a+jbUjYOA2dlaS8/qGeMS4DptYSTgIyl6do0HofPAi+penQGfbHorFNJ
Bs8NQ5uk0+yJePkrNKUw8mSmX/PlRGUhnX+Mv1v3BN09DIZAASp3Hfzi2R4zH6Ue
JopnngfR+xmy5/iDFEdJik1DkPaB3y6U+zHKmXokTQCxDMMZHPI0LXuaimt2Gle4
0z5vkTvVPKpnuXELqySiW7NZ1gk9+PJFraEvS1d+c57DCbJr2FpOlWtWcRnZjMpq
VAaN+siPROAyYPvLsdix6dR9ubiNy+W1tQ+DH0cdwqcI810cHWX262AW2yTiNkTM
KnucOaBZcbkiDhcUWRuaosbwotG/dz93ctsOcZ78IT7go7UjKDC82a4CCn/z4Fn+
+GJAOXoCuTTWierBysSsNbKH31+/l73Arf7CbjTGXp3E1Crmth9aYK3cceGlMnlY
RrbV3XXLlMvO4z6nplDsklsD+bEkB1Pp0KRqZClgT971ZAzFHTxxHCK7IHYfnRu6
2FX0VlVs/MYlUFgq+nyiuR1hYNgwEzCeOIdfCfgxEAZoQl3MsSwz8tdf7tMpOjbu
GcDGQP7x2IIQXOO/y7XO+NO0Vt2fD9nGBiwoGMrFMzF9RoEvpKzJJTJv6Lgg+7E7
LqTMc097Gb3vS1Iw2MoYzJXo4eMKxKoCdLs7nG/Qp+nd3il8ZgfbiGpv6Q/vSIyL
prOY1nD2r5Kc59JD99jJpq98/8lRdanoqBZPVKJTLhU1diOOWWj+vsUvt8DnTqpQ
I/QejuZ0aNtJU8kAQaVt6l1NIEV4gaCQYmGGZ7Ss1QRlxjtji1Gg3onsmYJJfH0a
8egqyOj+e6nrLpMyl7gRUMm+405rWocbLz+o9yu0H8FHBLU11SW6jtfN89GNK0A/
ke1DMdSCT6zNFbsZq4jti5fa8Usa6DQoo5dU7fCeVV+2k8K/kuVtWYA9ehZMHJNb
/e0zeTHCj6Vv2RjHoVmN1jVnjIjapZnCXEv2PevwxupXveyvFme3GeL6Cg+RvPxA
aLAUqTrjlI3jI7QtmInNrWVOTkDXuFOoWCm8jHGJaz/ms874OrRDbu3xLD7x5qc0
+abMh4dB7C3/PG/iO5dKssfDyg4cTtCp/OVTuTJFzGykBXtkPgn2H/PQZYJ9X7+q
xwoqxEHKn3Hioghk6oIOeH9wOyqwBzIxsqaFNBRj+n7MoL9vy2/PWXIIQVJWUPSz
hocalKtH/LT8YJV3E84aKeUhsSo01RtNjQep1wdoqrld3cmIoYvTu9r0eZVaH5JU
fREbJrS1K/3lrdxqJoQwAzByowxU5Zd3W8oovHyRSxDdCNJSAh37V+Xc6xfwKtE/
EULrGZIyawQTfkePLFnJAFVy1MMJAc2HZxyF233XXw+ztejRkTex/cGPyBm3/fpp
xyIXLgJjkmdwYNZBBOcydnjhiMF3oRpDWAj8ob4I3CnkAHuFxLiGX6rCXduizUNr
svyBOx2avLXLxuUEda4WjFwuoTWp0Fc7aj++lnjuBB86nd8l0ztDk7CKZ8UJ2qiv
iPlEJrz4Um7Cgcbt4EjbPrJMUaLU9uHlVCs0Uuq1DCw63UYcG/gnTT7iDC4eGduc
VtyXPFYXczP+Munj3mUypdzVTZx7H+JevnnIJUeLa0Y1AiAFuGG5jNRSXNjxjt2H
UIhIx9Gh9HLRUaqY2lx9QuJYhN+yCHDtP032Sn2cNNHHrwuRJeEYuNCzU601L9+s
OU6bwxTL3+BrqPfHMvSEqLb76L6KmJNDkBbZW2ZbESwZN0uYBISE11rm4lovQ/MP
kIujtd5wz1T7TqqWS0LevLyI83vtAnWlhWTmcKAjmNM0CrBPEeS451U2ahs6/ffJ
cFdpIGLVijn5slP//Oqo79/tO+O7H9CDCzaL4hSTP71t/OxbuXn8Ko966stoybTi
adfk5OjtLD6Xx3aQ9Ug4rRfbkmM0FMynG0aV2Z8aNdwtT6drYdDJAH0lsEFNenvm
n11yX9jD/6ea6+U+iYW3yQ8csBBwki6UOF9U0svuTFiI4uAMEGRvpmMW6cd86txi
vB4Mh3W2NbitsjUvOJcLFh+n0PNmgO5oRO0EULdekKy7tBSiZaeVlC0KF0rBN7XS
5ZFdLdyM5VwF5vGKXUqqsKvxUOCNoZHPAClOAskVSrPaq18Kq7ygl5dfjYdGrO3D
pfce2TvzvEiijZ5PPFTzcTG00oh0l7HOEG35Fl6u2BpUwMIqP1u/sYh6YNafTT4n
+6flWs5xy/yzuVOQ/cHpd+OL4XT1yLcIk0+QHxmrxSpO8LmQYT19oKwJ6tbkpP3z
W9zsW+osQQeT7LOba/QH0u/sleanRf0abaO4MSXoRRgG4G69NSidzwoemxeVRGU4
BIeMKP393TbT40wP3lXwjzLpWpmK3yFI72Cgik33sE1zg1Gthh1y/CtEwzpv5W05
0SwKwq6Z5AZ6UM3xWbPcawbJsw4vzyTKAOASip/c7ELg5LNqsljdjQYMjGPzf0a7
NUz8T8f4ckXUNKF9AsjUesZAvA4lMWMWO1l9RkbOAmB+Vwn2s7s96xwk/ZVlu8Vy
WHTU+Z2rM2caPXFgDEgz9ig2Jc5ErA1fRaYYTo9ABdmvKp2YhzzpiL8VM5NZ1n8w
VeLzCAB5DRWOaFp+YL0JOByK4oHpr8MshYdEh22lD7IFSydIWTvNBiepf4h8XGqI
yhXCasheMqygBwqvQQSZUMlI659M4VLpmi4ilcuEQqQoNpAhUcG4PtQ1ohtqYyWA
mXLlLgFS1XHmZYG+ucwG86SiGJjEhJ1+iRXblfNueQg73Q/3cSbXnkkZcRnPvs6+
itD2JkpQPkZwo/3ZQZH19agtkhl1x5v/PYyWoISVtZSj6rLlGLm90iQaSQ8LPZnp
mH0smyKQpxCI1qFPQzNKkUHhyF4CerboUB8Us94OCiBpT0Wr1HLUee/5wz3iNhiS
C5tdrdkX0rvf8yPoT50c1SW0CFJqye4rk4sQSliWRcRHm9OjuRy+bvMsgpe2vo/5
kqmL9ZuZYUHtQ9Jaj8SO1xH1sxj47XRtxRtj8yctImmsRhTCobkBME/5Rt03t7bP
o+p1VaXJm3O/S77smtiD5kN8UmblCjPjFiZVDt+p/z/2AgaofXRsP9nY+EufZRfP
6jQLHABNG0Sy3slm/WPyComwg1J+H3mSttC43N+r/9rhiuMIuE/tGiPlXcnD+T/4
ogPuAraFEARNsuxX8DWFBR6N8d0DpLyql9GDqMFEHAcG1BOi87zZl0lsCZOLBQT+
`pragma protect end_protected
