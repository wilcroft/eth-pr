// Benchmark "../allrules" written by ABC on Sat Dec  9 21:26:39 2017

module allrules  ( 
	xin, clock, z0_reg, xin_valid, z0_valid, z0_ready, xin_ready );
  input  [119:0] xin;
  input clock;
  input xin_valid;
  input z0_ready;
  output reg z0_reg, z0_valid;
  output xin_ready;
  
  reg [119:0] x;
  wire z0;
  reg x_valid;
  
  always@(posedge clock) 
  if (z0_ready||~z0_valid) begin
	x<= xin;
	z0_reg <= z0;
	x_valid <= xin_valid;
	z0_valid <= x_valid;
  end
  assign z0 = 1;
  //assign z0 = ((~x[034] & ((~x[032] & ((x[039] & ((~x[037] & ((x[043] & ((~x[033] & ((~x[035] & ~x[036] & x[040] & x[041]) | (x[035] & x[038] & ~x[041] & x[042]))) | (x[033] & ((~x[036] & ((~x[038] & (x[035] ? (x[040] ? (~x[041] & ~x[042]) : x[042]) : ~x[042])) | (~x[035] & x[038] & ((~x[041] & x[042]) | (x[040] & x[041] & ~x[042]))))) | (x[038] & ((~x[040] & ((x[035] & ~x[042] & (x[041] | (x[036] & ~x[041]))) | (~x[035] & x[036] & x[041] & x[042]))) | (~x[035] & x[036] & ((x[041] & ~x[042]) | (x[040] & ~x[041] & x[042]))))) | (x[036] & ~x[041] & ((~x[040] & x[042]) | (~x[035] & ~x[038] & x[040]))))) | (~x[042] & ((~x[038] & (x[035] ? (x[041] ? ~x[036] : ~x[040]) : (x[036] & x[041]))) | (~x[035] & ~x[036] & x[038] & ~x[040]))) | (x[035] & ~x[036] & x[040] & x[042] & (~x[038] ^ x[041])))) | (~x[036] & ((~x[043] & ((x[041] & ((x[033] & ((x[035] & x[040] & (~x[038] | (x[038] & x[042]))) | (~x[038] & ~x[040] & x[042]))) | (x[038] & x[040] & (~x[042] | (~x[033] & x[042]))) | (~x[033] & ~x[040] & (x[035] ^ ~x[042])))) | (~x[040] & ((~x[033] & ((x[038] & ~x[041] & x[042]) | (x[035] & ~x[042]))) | (~x[035] & ~x[041] & ((x[033] & x[038] & x[042]) | (~x[038] & ~x[042]))))) | (x[040] & ~x[041] & x[042] & ~x[035] & x[038]))) | (~x[033] & ~x[038] & ((~x[035] & ~x[040] & x[042]) | (~x[041] & ~x[042] & x[035] & x[040]))) | (x[038] & ((x[033] & ((x[042] & (x[035] ? (~x[041] | (~x[040] & x[041])) : (x[040] & x[041]))) | (~x[041] & ~x[042] & ~x[035] & x[040]))) | (x[041] & x[042] & ~x[035] & ~x[040]))))) | (x[036] & ((x[041] & (x[035] ? ((~x[043] & (x[033] ? (x[038] & x[040]) : (~x[038] ^ x[042]))) | (~x[038] & ((~x[040] & x[042]) | (x[033] & (x[040] | (~x[040] & ~x[042])))))) : ((x[042] & (x[033] ? (x[038] ? ~x[043] : x[040]) : ~x[038])) | (~x[038] & ~x[040] & ~x[042] & ~x[043])))) | (x[033] & (x[035] ? ((x[038] & x[042] & (x[040] ? ~x[041] : ~x[043])) | (~x[038] & x[040] & ~x[041] & ~x[043])) : (~x[042] & ((~x[038] & ~x[040] & ~x[041]) | (x[040] & ~x[043]))))))) | (~x[043] & ((~x[038] & ((x[033] & ~x[041] & (x[035] ? ~x[040] : (x[040] & x[042]))) | (x[040] & x[041] & ~x[042] & ~x[033] & ~x[035]))) | (x[035] & x[038] & ~x[041] & ~x[042] & (x[040] | (x[033] & ~x[040]))))))) | (x[037] & ((x[042] & ((x[041] & ((x[040] & (x[033] ? ((~x[035] & (~x[043] | (x[036] & x[043]))) | (x[038] & ~x[043] & x[035] & x[036])) : (x[035] ? x[038] : (x[036] & ~x[038])))) | (x[033] & ((x[038] & (x[035] ? (x[036] & x[043]) : (~x[036] & ~x[040]))) | (x[035] & ~x[043] & (x[036] ? ~x[038] : ~x[040])) | (~x[035] & ~x[038] & x[043] & (~x[036] | (x[036] & ~x[040]))))) | (x[035] & ~x[036] & ~x[038] & ~x[040] & x[043]))) | (x[038] & ((x[043] & ((x[033] & ((x[035] & ~x[036] & ~x[040]) | (x[036] & x[040] & ~x[041]))) | (x[040] & ((~x[033] & ~x[035] & x[036]) | (x[035] & ~x[036] & ~x[041]))))) | (~x[033] & ((~x[043] & (x[035] ? (x[040] ? ~x[041] : x[036]) : (x[036] & ~x[041]))) | (~x[035] & ~x[036] & ~x[040] & ~x[041]))))) | (~x[038] & ((~x[033] & ~x[035] & (x[040] ? ~x[041] : x[036])) | (x[035] & x[036] & ~x[041] & (x[040] ? x[043] : (~x[043] | (x[033] & x[043])))))) | (x[033] & x[036] & ~x[041] & ((x[040] & ~x[043]) | (~x[035] & ~x[040] & x[043]))))) | (~x[042] & ((~x[041] & ((x[035] & ((~x[040] & x[043] & x[033] & x[036]) | (~x[036] & ~x[038] & ~x[043]))) | (x[038] & ((~x[033] & x[043] & (x[036] | (~x[035] & ~x[036]))) | (~x[040] & ~x[043] & x[033] & ~x[036]))) | (~x[038] & ((~x[035] & (x[033] ? (x[040] | (~x[040] & x[043])) : (x[040] ? x[036] : ~x[043]))) | (~x[040] & x[043] & ~x[033] & x[036]))))) | (x[041] & (x[036] ? ((~x[035] & (x[033] ? ((x[040] & ~x[043]) | (~x[038] & (x[043] | (~x[040] & ~x[043])))) : (x[043] ? x[040] : ~x[038]))) | (x[033] & x[035] & x[038] & (x[040] | (~x[040] & x[043])))) : ((~x[033] & ((x[035] & x[043]) | (x[038] & x[040] & ~x[043]))) | (~x[040] & ((x[033] & (x[035] ? x[038] : x[043])) | (x[035] & ~x[038] & ~x[043]))) | (x[033] & x[040] & x[043])))) | (x[038] & (x[033] ? (x[040] & (x[035] ? (~x[036] & ~x[043]) : (x[036] & x[043]))) : (~x[035] & ~x[043] & (x[036] | (~x[036] & ~x[040]))))) | (x[035] & x[036] & ~x[038] & x[040] & ~x[043]))) | (~x[038] & (x[035] ? (x[040] & x[043] & (~x[036] ^ x[041])) : ((~x[036] & ((~x[033] & x[043] & (x[041] | (~x[040] & ~x[041]))) | (~x[040] & x[041] & ~x[043]))) | (x[033] & x[036] & ~x[040] & ~x[041] & ~x[043])))) | (~x[033] & x[043] & ((x[035] & ~x[040] & (~x[036] ^ x[041])) | (~x[035] & ~x[036] & x[038] & x[040] & x[041]))))) | (~x[043] & (x[033] ? ((~x[035] & ~x[040] & ((x[036] & (x[038] ? ~x[041] : (x[041] & x[042]))) | (x[041] & ~x[042] & ~x[036] & x[038]))) | (x[040] & ~x[041] & x[042] & x[035] & ~x[036] & ~x[038])) : (x[040] & ~x[042] & (x[035] ? (x[041] & (x[036] ^ ~x[038])) : (~x[036] & ~x[041]))))) | (~x[036] & ((~x[033] & x[040] & ((x[035] & ((~x[038] & x[041] & x[042]) | (x[038] & ~x[041] & ~x[042] & x[043]))) | (~x[035] & ~x[038] & ~x[041] & ~x[042] & x[043]))) | (x[033] & ~x[035] & ~x[038] & ~x[041] & x[042] & x[043]))))) | (~x[039] & ((~x[033] & ((x[035] & ((x[038] & ((~x[041] & ((~x[037] & (x[036] ? (x[043] ? ~x[042] : ~x[040]) : x[043])) | (~x[036] & ~x[040] & ((~x[042] & ~x[043]) | (x[037] & (x[042] | (~x[042] & x[043]))))))) | (x[040] & (x[036] ? (x[042] & ~x[043]) : ((x[037] & x[042] & x[043]) | (x[041] & ~x[042] & ~x[043])))) | (x[041] & ((x[036] & ((x[042] & x[043]) | (x[037] & ~x[040] & ~x[042]))) | (~x[042] & x[043] & ~x[036] & x[037]))))) | (~x[038] & ((~x[036] & ((x[037] & x[041]) | (~x[041] & ~x[043] & ~x[037] & ~x[040]))) | (x[036] & ((~x[043] & ((x[037] & (x[041] ? ~x[042] : x[040])) | (~x[041] & (x[042] ? ~x[040] : ~x[037])))) | (x[043] & (x[040] ? (x[041] ? ~x[037] : ~x[042]) : (x[041] & ~x[042]))) | (~x[040] & x[041] & x[042]))) | (~x[037] & ((~x[040] & ~x[041] & ~x[042] & x[043]) | (x[040] & x[041] & x[042] & ~x[043]))) | (~x[041] & ~x[042] & x[037] & ~x[040]))) | (~x[042] & ((~x[036] & x[040] & ~x[041] & (~x[037] ^ x[043])) | (x[041] & ~x[043] & x[036] & ~x[037]))))) | (~x[035] & ((x[041] & ((~x[038] & (x[043] ? ((x[040] & (x[042] ? ~x[037] : ~x[036])) | (x[037] & ~x[040] & x[042])) : (x[036] ? (x[040] | (x[037] & ~x[040] & ~x[042])) : (x[037] & x[042])))) | (~x[040] & ((~x[037] & (x[036] ? (x[042] ? x[038] : ~x[043]) : (x[042] & ~x[043]))) | (x[038] & x[042] & (x[043] ? ~x[036] : x[037])))) | (x[036] & x[038] & (x[037] ? (~x[042] & ~x[043]) : ((~x[042] & x[043]) | (x[040] & x[042] & ~x[043])))))) | (~x[041] & ((x[036] & ((~x[040] & ((x[037] & ((~x[042] & ~x[043]) | (~x[038] & x[042] & x[043]))) | (x[038] & ~x[042] & x[043]))) | (~x[037] & x[038] & (~x[043] | (x[040] & x[043]))))) | (x[037] & ((~x[038] & x[040] & (x[043] ? ~x[042] : ~x[036])) | (~x[036] & ((x[038] & x[042]) | (~x[040] & ~x[042] & x[043]))))))) | (~x[040] & ((x[036] & ~x[038] & x[043] & (~x[037] | (x[037] & ~x[042]))) | (~x[036] & ~x[037] & x[038] & ~x[042]))) | (~x[036] & x[037] & x[038] & x[040] & ~x[042]))) | (~x[042] & ((x[041] & ((~x[036] & x[038] & (x[037] ? (~x[040] & ~x[043]) : (x[040] & x[043]))) | (x[036] & x[037] & ~x[038] & x[040] & x[043]))) | (~x[036] & ~x[037] & ~x[038] & x[040] & ~x[041] & x[043]))) | (~x[036] & ~x[037] & x[038] & x[040] & ~x[041] & x[042] & ~x[043]))) | (x[033] & ((x[041] & ((x[036] & ((~x[040] & ((x[042] & x[043] & x[037] & x[038]) | (~x[038] & ~x[043] & x[035] & ~x[037]))) | (~x[035] & ((x[040] & (x[037] ? (x[038] & (x[043] | (x[042] & ~x[043]))) : (x[043] ? ~x[042] : ~x[038]))) | (x[042] & x[043] & ~x[037] & x[038]))) | (x[035] & ((x[040] & (x[037] ? (x[038] | (~x[038] & ~x[042])) : (x[038] ? (~x[042] & ~x[043]) : x[042]))) | (~x[042] & x[043] & ~x[037] & ~x[038]))))) | (x[037] & ((~x[036] & ((x[035] & (x[038] ? (x[040] & ~x[043]) : (~x[040] & ~x[042]))) | (~x[035] & ((x[040] & x[042] & ~x[043]) | (x[038] & ~x[040] & x[043]))) | (~x[038] & x[040] & ~x[042]))) | (x[035] & ~x[038] & x[042]) | (~x[035] & x[038] & x[040] & ~x[042] & ~x[043]))) | (~x[043] & ((~x[035] & ~x[036] & x[038] & ~x[040] & x[042]) | (x[035] & ~x[037] & ~x[038] & x[040] & ~x[042]))) | (~x[036] & ((~x[042] & ((x[038] & ((x[035] & (x[040] ? ~x[037] : x[043])) | (~x[040] & x[043] & ~x[035] & ~x[037]))) | (~x[035] & ((~x[038] & ~x[040] & x[043]) | (~x[037] & x[040]))))) | (~x[035] & ~x[037] & x[042] & (x[038] ? (x[040] & x[043]) : ~x[040])))))) | (~x[037] & ((~x[041] & ((x[036] & ((x[043] & ((x[035] & ((~x[040] & ~x[042]) | (~x[038] & x[040] & x[042]))) | (~x[035] & ~x[038] & x[040] & ~x[042]))) | (~x[038] & ((~x[035] & ~x[040] & x[042]) | (x[040] & ~x[043]))))) | (x[040] & ((~x[036] & ((~x[038] & x[042] & x[043]) | (~x[042] & (x[035] ? (~x[038] | (x[038] & ~x[043])) : x[043])))) | (~x[035] & x[038] & ~x[042] & ~x[043]))) | (x[035] & ~x[036] & x[038] & x[042] & x[043]))) | (~x[043] & ((~x[036] & (x[035] ? (~x[038] & (x[042] | (~x[040] & ~x[042]))) : ((x[040] & x[042]) | (x[038] & ~x[040] & ~x[042])))) | (x[036] & x[038] & x[042]) | (~x[040] & ~x[042] & ~x[035] & ~x[038]))) | (~x[035] & x[036] & x[043] & ((~x[040] & ~x[042]) | (~x[038] & x[040] & x[042]))))) | (x[037] & ((~x[036] & (((x[043] | (~x[040] & ~x[043])) & ((x[035] & x[038] & x[042]) | (~x[038] & ~x[041] & ~x[042]))) | (~x[041] & ((x[040] & ~x[042] & ~x[043]) | (~x[035] & (x[038] ? (x[040] ? (x[042] & x[043]) : ~x[043]) : (x[040] & x[042]))))))) | (~x[041] & ((x[042] & (x[035] ? (~x[038] & (x[043] ? x[040] : x[036])) : (x[038] & (~x[040] ^ ~x[043])))) | (x[036] & (x[035] ? (~x[042] & (x[040] ? ~x[043] : ~x[038])) : (x[040] & x[043]))))) | (~x[035] & x[036] & ~x[038] & (x[040] ? (x[042] & ~x[043]) : ~x[042])))) | (~x[036] & ~x[041] & ((x[042] & (x[035] ? (x[038] ? (x[040] & ~x[043]) : (~x[040] & x[043])) : (~x[038] & ~x[040]))) | (~x[035] & x[038] & ~x[040] & ~x[042] & x[043]))))) | (~x[035] & ((~x[036] & ((~x[041] & x[042] & x[043] & ~x[037] & x[038] & x[040]) | (x[041] & ~x[042] & ~x[043] & x[037] & ~x[038] & ~x[040]))) | (x[037] & ((x[036] & ~x[041] & ~x[043] & ((~x[040] & x[042]) | (~x[038] & x[040] & ~x[042]))) | (~x[038] & x[040] & x[041] & x[042] & x[043]))) | (x[036] & ~x[038] & ~x[040] & x[041] & x[042] & ~x[043]))) | (x[035] & ((x[038] & ((~x[040] & ((x[036] & ~x[041] & x[043] & (x[037] | (~x[037] & x[042]))) | (x[042] & ~x[043] & ~x[036] & ~x[037]))) | (~x[036] & ~x[037] & x[040] & x[041] & x[042]))) | (~x[036] & ~x[037] & ~x[038] & x[041] & x[043]))))) | (x[042] & (x[036] ? ((x[038] & ((~x[040] & ((x[033] & x[041] & ((x[037] & ~x[043]) | (x[035] & ~x[037] & x[043]))) | (~x[033] & ~x[035] & x[037] & x[043]))) | (x[040] & ~x[041] & x[043] & ~x[033] & x[035] & x[037]))) | (~x[033] & ~x[038] & ((x[035] & (x[037] ? (x[040] ? (x[041] & ~x[043]) : (~x[041] & x[043])) : (~x[041] & x[043]))) | (~x[041] & ~x[043] & ~x[037] & x[040])))) : ((~x[033] & ((~x[038] & ((x[035] & ~x[041] & ((x[040] & ~x[043]) | (~x[037] & ~x[040] & x[043]))) | (~x[035] & ~x[037] & x[040] & x[041] & ~x[043]))) | (~x[035] & x[038] & ((~x[037] & ~x[040] & ~x[041] & x[043]) | (x[041] & ~x[043] & x[037] & x[040]))))) | (x[033] & ~x[035] & x[037] & x[038] & x[040] & x[041] & x[043])))) | (~x[042] & ((x[043] & (x[038] ? (x[037] ? (x[033] ? (~x[041] & (x[035] ? (~x[036] & ~x[040]) : (~x[036] ^ ~x[040]))) : (x[041] & (x[035] ? (x[036] & x[040]) : ~x[040]))) : (x[040] & ~x[041] & (x[033] ? x[036] : (~x[035] & ~x[036])))) : ((~x[033] & ~x[035] & ~x[036] & ~x[037] & ~x[040]) | (x[033] & x[035] & x[036] & x[037] & x[040] & ~x[041])))) | (x[033] & ~x[043] & ((x[036] & x[037] & ((~x[040] & (x[035] ? (x[038] | (~x[038] & x[041])) : (x[038] & x[041]))) | (~x[035] & x[038] & x[040] & ~x[041]))) | (~x[035] & ~x[036] & ~x[037] & ~x[038] & x[040] & ~x[041]))))) | (~x[033] & ~x[035] & x[036] & ~x[037] & ~x[038] & ~x[040] & ~x[041] & ~x[043]))) | (x[032] & ((x[040] & ((~x[037] & ((~x[036] & ((~x[042] & ((~x[038] & x[041] & x[043] & ~x[033] & x[035]) | (x[033] & ~x[035] & x[038] & ~x[041] & ~x[043]))) | (~x[041] & (x[035] ? ((x[038] & (x[033] ? (x[042] & (x[043] | (~x[039] & ~x[043]))) : (x[039] ^ ~x[043]))) | (x[033] & x[039] & (x[043] ? ~x[038] : x[042])) | (~x[038] & ~x[039] & x[043])) : ((x[043] & (x[033] ? (x[039] | (~x[038] & ~x[039] & x[042])) : (x[038] ^ x[039]))) | (x[042] & ~x[043] & (x[039] ? ~x[038] : x[033]))))) | (x[041] & ((~x[038] & ((~x[033] & x[042] & (x[043] | (~x[039] & ~x[043]))) | (x[039] & ~x[043]))) | (x[033] & ((~x[035] & ((~x[039] & ~x[043]) | (x[038] & x[039] & x[043]))) | (x[042] & x[043] & x[035] & x[039]))) | (x[035] & x[038] & (~x[043] | (~x[039] & x[043]))))) | (~x[033] & ~x[035] & x[038] & x[039] & ~x[043]))) | (x[033] & ((x[036] & ((~x[041] & ((x[035] & (x[038] ? (x[042] & ~x[043]) : (~x[042] & x[043]))) | (~x[039] & (x[038] ? (x[043] ? ~x[042] : ~x[035]) : (x[042] & x[043]))) | (~x[035] & x[039] & (~x[042] | (~x[038] & x[042] & x[043]))))) | (~x[038] & (x[035] ? x[041] : (x[039] & (x[043] ? x[041] : x[042])))) | (x[035] & x[038] & x[041] & (x[039] | (~x[039] & x[042]))))) | (~x[035] & ((~x[039] & ((~x[038] & ~x[042] & (x[043] | (~x[041] & ~x[043]))) | (x[042] & x[043] & (x[041] | (x[038] & ~x[041]))))) | (x[038] & x[039] & ~x[043] & (x[041] | (~x[041] & x[042]))))) | (x[035] & ~x[041] & (x[038] ? (~x[042] & (~x[043] | (x[039] & x[043]))) : (~x[039] & ~x[043]))))) | (x[035] & ((x[039] & ((x[041] & x[042] & x[043] & ~x[033] & x[038]) | (~x[041] & ~x[043] & x[036] & ~x[038]))) | (~x[039] & ((~x[042] & ((~x[033] & x[043] & (x[038] ? ~x[041] : x[036])) | (x[041] & ~x[043] & x[036] & x[038]))) | (~x[033] & x[036] & ~x[038] & ~x[041] & (~x[043] | (x[042] & x[043]))))) | (x[041] & ~x[042] & ~x[043] & ~x[033] & x[036] & ~x[038]))) | (x[036] & ((~x[033] & ((~x[035] & ((~x[039] & (x[038] ? (~x[042] & x[043]) : (x[042] & ~x[043]))) | (x[039] & (x[038] ? (x[042] | (x[041] & ~x[042] & ~x[043])) : (x[041] ? x[042] : ~x[043]))) | (~x[042] & ~x[043] & x[038] & ~x[041]))) | (x[038] & ((~x[042] & x[043] & x[039] & x[041]) | (x[042] & ~x[043] & ~x[039] & ~x[041]))) | (x[041] & x[042] & x[043] & ~x[038] & ~x[039]))) | (~x[035] & x[041] & ~x[043] & (x[038] ? (~x[039] & x[042]) : ~x[042])))) | (~x[033] & ~x[035] & ~x[038] & x[041] & ~x[042] & x[043]))) | (~x[033] & ((x[037] & ((x[035] & ((~x[036] & ((x[039] & ((x[038] & (x[041] ? ~x[043] : (x[042] & x[043]))) | (~x[043] & (x[042] ? ~x[038] : ~x[041])))) | (x[041] & (x[038] ? (~x[042] & x[043]) : (x[042] ? ~x[039] : ~x[043]))))) | (x[036] & ((x[042] & ((x[038] & ~x[043] & (x[039] | (~x[039] & ~x[041]))) | (x[039] & ~x[041] & x[043]))) | (x[038] & ~x[039] & x[041] & ~x[042] & x[043]))) | (~x[041] & ~x[042] & x[043] & x[038] & x[039]))) | (~x[035] & ((x[039] & ((x[041] & ((x[038] & x[042] & x[043]) | (~x[042] & ~x[043] & ~x[036] & ~x[038]))) | (~x[038] & (x[036] ? x[042] : ((~x[042] & x[043]) | (~x[041] & x[042] & ~x[043])))) | (x[038] & (x[036] ? (~x[043] | (~x[042] & x[043])) : (~x[042] & ~x[043]))))) | (~x[042] & (x[036] ? (~x[038] & ((~x[041] & x[043]) | (~x[039] & x[041] & ~x[043]))) : (~x[039] & (x[041] ^ ~x[043])))) | (~x[041] & x[042] & ~x[038] & ~x[039]))) | (x[041] & ((x[036] & ~x[038] & x[039] & ~x[042]) | (~x[036] & x[038] & ~x[039] & x[042] & x[043]))))) | (~x[036] & ((~x[039] & ~x[041] & ((x[035] & (x[038] ? (x[042] & x[043]) : ~x[043])) | (~x[042] & x[043] & ~x[035] & ~x[038]))) | (~x[035] & x[038] & x[039] & ~x[042] & x[043]))) | (x[035] & x[036] & x[041] & x[042] & (x[038] ? ~x[039] : ~x[043])))) | (x[035] & ((x[037] & ((x[033] & ((x[036] & ((x[038] & (x[039] ? (~x[041] & x[042]) : ~x[042])) | (~x[038] & ~x[043] & (x[041] ? x[042] : x[039])) | (x[039] & x[041] & ~x[042]))) | (x[039] & ((x[038] & ((x[041] & x[042] & ~x[043]) | (~x[036] & (x[041] ? x[043] : ~x[042])))) | (~x[036] & ~x[041] & x[042] & x[043]))) | (x[041] & x[042] & x[038] & ~x[039]))) | (~x[042] & ((~x[038] & ((x[036] & ~x[039] & (~x[041] | (x[041] & ~x[043]))) | (x[041] & x[043] & ~x[036] & x[039]))) | (~x[036] & x[038] & ~x[039] & ~x[041] & ~x[043]))) | (~x[041] & x[042] & x[043] & x[036] & ~x[038] & ~x[039]))) | (~x[039] & x[041] & ~x[043] & x[033] & ~x[036] & ~x[038]))) | (x[037] & ((x[033] & ((~x[035] & ((~x[042] & (x[038] ? ((~x[039] & ~x[041]) | (~x[036] & x[039] & x[043])) : ((x[039] & (x[036] ? x[041] : ~x[043])) | (~x[036] & (x[041] ? ~x[039] : x[043]))))) | (~x[043] & ((x[036] & x[038] & (x[041] | (~x[041] & x[042]))) | (~x[038] & (x[039] ? x[042] : (~x[041] | (x[041] & x[042])))))) | (x[041] & x[042] & ~x[036] & x[038]) | (x[036] & ~x[038] & ~x[039] & x[043]))) | (x[038] & ((~x[036] & ~x[039] & (x[041] ? (~x[042] & ~x[043]) : x[042])) | (~x[041] & ~x[042] & x[036] & x[039]))) | (x[036] & ~x[038] & x[039] & x[043] & (~x[041] | (x[041] & x[042]))))) | (~x[041] & ((~x[035] & ~x[038] & x[039] & (x[036] ? (~x[042] & ~x[043]) : (x[042] & x[043]))) | (x[036] & x[038] & ~x[039] & x[042] & x[043]))) | (~x[035] & ~x[036] & ~x[038] & x[042] & x[043] & ~x[039] & x[041]))) | (x[033] & ~x[035] & x[043] & ((x[036] & x[038] & (x[042] ? x[039] : x[041])) | (~x[036] & ~x[038] & x[039] & x[041]))))) | (~x[040] & ((~x[038] & ((x[033] & ((x[035] & ((x[037] & (x[041] ? ((x[039] & ~x[042]) | (~x[036] & ~x[039] & ~x[043])) : (x[043] & (x[036] ? (~x[042] | (~x[039] & x[042])) : (x[039] & x[042]))))) | (~x[037] & ((x[036] & x[039] & (x[043] | (~x[042] & ~x[043]))) | (~x[039] & x[041] & ~x[043]) | (~x[036] & ~x[041] & (x[042] | (~x[042] & ~x[043]))))) | (x[039] & x[041] & x[042] & (x[036] ^ x[043])))) | (~x[035] & ((~x[039] & ((~x[043] & ((x[036] & (x[037] ? x[041] : ~x[042])) | (~x[041] & (x[042] ? ~x[036] : x[037])))) | (~x[036] & ~x[042] & (x[037] ? x[043] : x[041])) | (~x[037] & x[042] & x[043]))) | (x[037] & ((x[041] & (x[036] ? (x[039] & x[042]) : (x[043] ? x[039] : ~x[042]))) | (x[036] & ((~x[042] & x[043]) | (~x[041] & x[042] & ~x[043]))) | (x[042] & x[043] & x[039] & ~x[041]))) | (x[039] & ((~x[037] & ~x[041] & x[043]) | (x[036] & ~x[042] & ~x[043]))))) | (x[041] & ~x[042] & x[043] & x[036] & ~x[037] & ~x[039]))) | (~x[033] & ((~x[037] & ((~x[041] & ((x[035] & (x[036] ? (~x[042] & x[043]) : ~x[039])) | (~x[042] & ~x[043] & x[036] & x[039]))) | (x[043] & ((~x[035] & (x[036] ? (x[041] & (~x[042] | (~x[039] & x[042]))) : x[039])) | (x[041] & ~x[042] & ~x[036] & ~x[039]))) | (x[041] & ((x[036] & x[039] & x[042]) | (~x[035] & ~x[043] & (x[039] ? ~x[042] : x[036])))))) | (x[035] & ((~x[041] & ((x[042] & x[043] & x[036] & ~x[039]) | (~x[042] & ~x[043] & ~x[036] & x[037]))) | (x[043] & ((x[036] & x[037] & (~x[042] | (~x[039] & x[041] & x[042]))) | (x[041] & ~x[042] & ~x[036] & x[039]))) | (x[041] & x[042] & ~x[036] & ~x[039]))) | (~x[035] & ((x[037] & ((x[039] & (x[036] ? (x[041] ? (x[042] & ~x[043]) : (~x[042] & x[043])) : (x[042] & x[043]))) | (x[041] & ((~x[036] & (x[042] ? ~x[039] : x[043])) | (~x[039] & ~x[042] & ~x[043]))) | (~x[041] & x[043] & ~x[036] & ~x[039]))) | (~x[041] & x[042] & ~x[043] & (x[039] | (x[036] & ~x[039]))))) | (x[041] & ~x[042] & ~x[043] & ~x[036] & x[037] & x[039]))) | (~x[036] & ((~x[035] & ((~x[041] & ~x[042] & x[043] & x[037] & x[039]) | (x[042] & ~x[043] & ~x[037] & x[041]))) | (x[039] & ((~x[041] & ~x[042] & x[043] & x[035] & ~x[037]) | (x[042] & ~x[043] & x[037] & x[041]))))) | (x[035] & x[036] & ((x[042] & ((x[037] & (x[039] ? (~x[041] & x[043]) : (x[041] & ~x[043]))) | (x[039] & ~x[041] & ~x[043]))) | (~x[042] & ~x[043] & x[037] & ~x[039]))))) | (x[038] & ((x[037] & ((x[039] & ((x[041] & ((x[036] & ~x[042] & x[043]) | (x[033] & ~x[036] & x[042] & ~x[043]))) | (x[043] & ((x[033] & ((~x[036] & x[042]) | (x[035] & x[036] & ~x[041]))) | (~x[035] & ((~x[033] & (x[036] ^ ~x[042])) | (x[036] & ~x[041] & ~x[042]))) | (x[035] & ~x[036] & ~x[042]))) | (~x[043] & ((x[036] & ((x[033] & (~x[042] | (x[035] & x[042]))) | (~x[041] & x[042] & ~x[033] & ~x[035]))) | (~x[041] & ~x[042] & ~x[033] & x[035]))) | (x[033] & ~x[035] & x[036] & x[042]))) | (~x[039] & ((~x[041] & (x[043] ? (x[033] ? (~x[036] | (x[036] & ~x[042])) : (x[035] & x[042])) : (x[036] ? ~x[042] : (x[042] | (~x[033] & x[035] & ~x[042]))))) | (~x[035] & ((x[033] & x[042] & (x[036] ? ~x[043] : x[041])) | (x[036] & x[041] & ~x[042] & ~x[043]))) | (x[035] & x[041] & ((x[042] & x[043]) | (x[033] & (~x[043] | (~x[042] & x[043]))))))) | (~x[035] & ~x[036] & ((~x[042] & (x[033] ? (x[041] ^ ~x[043]) : (x[041] & ~x[043]))) | (x[042] & x[043] & ~x[033] & ~x[041]))))) | (~x[036] & ((x[039] & ((~x[041] & ((x[033] & ((~x[037] & x[042] & x[043]) | (x[035] & ~x[042] & ~x[043]))) | (x[043] & ((~x[033] & x[035] & x[042]) | (~x[035] & ~x[037] & ~x[042]))))) | (~x[037] & ((~x[035] & ((x[042] & ~x[043]) | (~x[033] & x[041] & ~x[042]))) | (~x[042] & x[043] & x[035] & x[041]))))) | (~x[037] & ((~x[043] & ((~x[042] & ((~x[033] & (x[035] | (~x[035] & ~x[041]))) | (~x[035] & ~x[039] & x[041]))) | (x[035] & x[042] & (x[041] ? ~x[039] : x[033])))) | (x[035] & x[043] & ((x[033] & x[041] & (x[042] | (~x[039] & ~x[042]))) | (~x[039] & ~x[041] & x[042]))))) | (~x[033] & ~x[035] & ~x[039] & x[041] & (x[042] | (~x[042] & x[043]))))) | (x[036] & (x[035] ? ((~x[042] & ((~x[033] & ~x[039] & x[041]) | (x[039] & x[043] & x[033] & ~x[037]))) | (~x[037] & ((~x[043] & ((~x[041] & (~x[033] | (x[033] & (x[039] | (~x[039] & x[042]))))) | (~x[033] & x[039] & x[041]))) | (x[033] & x[041] & x[042]))) | (~x[041] & x[042] & x[043] & x[033] & ~x[039])) : (~x[037] & (x[041] ? (~x[033] | (x[033] & ~x[039] & x[043])) : (x[042] | (x[039] & ~x[042] & ~x[043])))))) | (~x[039] & ((~x[041] & ~x[042] & x[043] & ~x[033] & x[035]) | (x[041] & x[042] & ~x[043] & x[033] & ~x[035] & ~x[037]))))) | (~x[033] & ((~x[036] & (x[035] ? (x[041] & (x[037] ? (~x[039] & ~x[042]) : (x[039] & x[042]))) : (~x[041] & ~x[042] & (x[037] ? (x[039] & ~x[043]) : (~x[039] & x[043]))))) | (~x[035] & x[036] & x[037] & (x[039] ? (~x[042] & ~x[043]) : (x[041] ? x[042] : x[043]))))) | (x[033] & ((~x[035] & ((x[036] & x[042] & ((~x[041] & x[043] & x[037] & ~x[039]) | (x[041] & ~x[043] & ~x[037] & x[039]))) | (~x[037] & ((~x[036] & ~x[042] & ~x[043] & (~x[039] ^ x[041])) | (x[039] & x[041] & x[043]))))) | (~x[037] & ((~x[041] & ~x[042] & x[043] & x[036] & ~x[039]) | (x[041] & x[042] & ~x[043] & x[035] & ~x[036] & x[039]))))))) | (x[043] & ((~x[039] & ((x[037] & ((~x[035] & ((~x[033] & ~x[042] & (x[036] ? x[041] : (x[038] & ~x[041]))) | (x[033] & x[036] & x[038] & x[041] & x[042]))) | (x[033] & ~x[038] & ((x[035] & x[041] & (x[042] | (x[036] & ~x[042]))) | (~x[036] & ~x[041] & x[042]))))) | (x[033] & ~x[036] & ((x[035] & ~x[038] & x[041] & (~x[042] | (~x[037] & x[042]))) | (x[038] & ~x[042] & ~x[035] & ~x[037]))))) | (x[039] & ((~x[033] & ((x[042] & ((~x[036] & (x[035] ? (x[037] & (~x[038] | (x[038] & x[041]))) : (~x[037] & x[038]))) | (~x[038] & ~x[041] & x[036] & ~x[037]))) | (~x[038] & ~x[041] & ~x[042] & ~x[035] & x[036] & ~x[037]))) | (x[035] & ((x[036] & x[038] & x[042] & (~x[037] ^ x[041])) | (x[033] & ~x[036] & ~x[037] & ~x[038] & x[041] & ~x[042]))))) | (~x[038] & ~x[041] & ~x[042] & x[035] & ~x[036] & x[037]))) | (~x[043] & (x[038] ? ((~x[033] & ~x[041] & x[042] & ((x[035] & ~x[036] & x[039]) | (~x[035] & x[036] & x[037] & ~x[039]))) | (x[039] & x[041] & ~x[042] & x[033] & ~x[036] & x[037])) : ((~x[041] & (x[035] ? ((~x[036] & ((x[033] & x[037] & (~x[042] | (x[039] & x[042]))) | (x[039] & ~x[042] & ~x[033] & ~x[037]))) | (x[036] & x[037] & ~x[039] & x[042])) : (~x[042] & ((~x[036] & ~x[037] & x[039]) | (~x[033] & x[036] & x[037] & ~x[039]))))) | (x[033] & ~x[035] & x[036] & ~x[037] & ~x[039] & x[042])))) | (~x[036] & ~x[037] & ~x[033] & x[035] & ~x[041] & x[042] & ~x[038] & x[039]))) | (~x[042] & ((x[035] & ((~x[043] & ((x[039] & (((x[040] ^ x[041]) & ((~x[033] & x[036] & x[037] & x[038]) | (x[033] & ~x[036] & ~x[037] & ~x[038]))) | (~x[038] & ~x[040] & ~x[041] & x[036] & x[037]))) | (~x[039] & ((~x[041] & ((x[033] & ~x[040] & (x[036] ? ~x[037] : (x[037] & x[038]))) | (x[038] & x[040] & ~x[033] & x[036]))) | (~x[033] & x[040] & x[041] & (x[036] ? (x[037] & x[038]) : (~x[037] & ~x[038]))))) | (x[033] & ~x[036] & ~x[037] & x[038] & ~x[040] & x[041]))) | (x[043] & (x[036] ? ((~x[033] & ((x[040] & ~x[041] & (x[037] ? (x[038] ^ x[039]) : (x[038] & x[039]))) | (~x[037] & ~x[038] & x[039] & x[041]))) | (~x[037] & x[038] & ~x[039] & x[041] & (x[040] | (x[033] & ~x[040])))) : (x[038] & ((~x[037] & ((x[033] & ~x[041] & (x[039] ^ x[040])) | (x[041] & ((x[039] & x[040]) | (~x[033] & ~x[039] & ~x[040]))))) | (~x[039] & x[040] & x[033] & x[037]))))) | (x[033] & ~x[036] & ~x[037] & ~x[040] & ~x[041] & x[038] & ~x[039]))) | (~x[035] & ((~x[040] & (x[033] ? (x[038] & (((~x[036] ^ x[043]) & (x[037] ? (~x[039] & x[041]) : (x[039] & ~x[041]))) | (~x[041] & ((~x[036] & x[037] & x[039] & x[043]) | (x[036] & ~x[037] & ~x[039] & ~x[043]))))) : ((~x[036] & ~x[039] & ~x[041] & ~x[043] & (~x[038] | (x[037] & x[038]))) | (x[039] & x[041] & x[043] & x[036] & x[037] & ~x[038])))) | (~x[039] & x[040] & (x[037] ? ((x[041] & ((x[033] & (x[036] ? (~x[038] & ~x[043]) : (x[038] & x[043]))) | (~x[038] & ~x[043] & ~x[033] & ~x[036]))) | (~x[033] & x[036] & x[038] & ~x[041])) : ((x[041] & ~x[043] & x[036] & x[038]) | (~x[033] & (x[036] ? (~x[038] & ~x[041]) : ~x[043]))))))) | (~x[037] & ~x[040] & ((x[033] & ((x[041] & ~x[043] & x[036] & x[038]) | (~x[036] & ~x[038] & ~x[039] & ~x[041] & x[043]))) | (~x[039] & x[041] & ~x[043] & ~x[033] & ~x[036] & ~x[038]))))) | (x[042] & (x[037] ? (x[039] ? (x[041] ? ((~x[038] & ((x[033] & x[035] & x[043] & (~x[036] ^ ~x[040])) | (~x[033] & ~x[035] & ~x[036] & x[040] & ~x[043]))) | (~x[033] & ~x[035] & x[038] & ~x[040] & ~x[043])) : ((x[038] & (x[033] ? (~x[036] & (x[040] ? (x[035] ^ x[043]) : ~x[043])) : ((~x[035] & ~x[036] & x[040]) | (x[035] & x[036] & ~x[040] & x[043])))) | (~x[038] & x[040] & ~x[043] & ~x[033] & x[035] & x[036]))) : (x[038] ? ((~x[033] & ((x[036] & (x[035] ? (~x[040] & ~x[043]) : (x[040] & x[041]))) | (x[035] & ~x[036] & ~x[043] & (x[041] | (x[040] & ~x[041]))))) | (x[033] & x[035] & x[036] & ~x[041] & ~x[043])) : ((x[035] & ((x[040] & ((~x[033] & x[043] & (~x[036] ^ x[041])) | (~x[041] & ~x[043] & x[033] & ~x[036]))) | (~x[041] & ~x[043] & ~x[036] & ~x[040]))) | (x[033] & ~x[035] & ~x[040] & x[041] & (~x[036] | (x[036] & x[043])))))) : (x[035] ? (x[036] & (((x[039] ? (x[040] & ~x[041]) : (~x[040] & x[041])) & (x[033] ? (~x[038] & x[043]) : (x[038] & ~x[043]))) | (x[043] & ((~x[033] & x[039] & x[041] & (x[038] ^ x[040])) | (x[040] & ~x[041] & x[038] & ~x[039]))) | (x[033] & ~x[038] & ~x[039] & ~x[040] & ~x[041]))) : ((~x[040] & ((x[033] & ((~x[036] & x[038] & ~x[039] & x[043]) | (~x[041] & ~x[043] & ~x[038] & x[039]))) | (~x[036] & ~x[039] & ((x[038] & ~x[041] & ~x[043]) | (~x[033] & ~x[038] & x[043]))))) | (~x[033] & ~x[039] & ((~x[036] & ~x[043] & (x[038] ? (x[040] & x[041]) : ~x[041])) | (x[040] & x[043] & ((x[038] & x[041]) | (x[036] & ~x[038] & ~x[041]))))))))) | (x[037] & x[039] & ~x[043] & ((x[035] & x[041] & ((~x[033] & ~x[040] & (~x[036] ^ ~x[038])) | (~x[038] & x[040] & x[033] & ~x[036]))) | (x[033] & ~x[035] & ~x[036] & ~x[041] & (~x[038] ^ x[040])))))) | (x[034] & ((~x[032] & ((~x[037] & ((x[035] & ((x[043] & ((~x[033] & (x[038] ? ((~x[040] & ~x[041] & x[042]) | (x[040] & x[041] & ~x[042] & x[036] & ~x[039])) : (x[039] ? ((~x[040] & (x[041] ? ~x[042] : x[036])) | (~x[036] & ~x[041] & ~x[042])) : ((x[036] & (x[040] ? x[042] : x[041])) | (~x[040] & ~x[041] & x[042]) | (~x[036] & ~x[042] & (x[041] | (x[040] & ~x[041]))))))) | (x[039] & ((~x[041] & ((~x[038] & x[040] & x[042]) | (x[033] & ~x[036] & ~x[040]))) | (~x[042] & ((x[033] & ((x[036] & (x[038] ^ x[040])) | (~x[040] & x[041] & ~x[036] & ~x[038]))) | (x[040] & x[041] & ~x[036] & x[038]))) | (x[033] & x[041] & x[042] & (x[038] ? (~x[036] | (x[036] & ~x[040])) : ~x[040])))) | (x[033] & ((~x[039] & (x[036] ? (x[042] & (x[040] ^ x[041])) : (~x[042] & (x[040] ? ~x[041] : ~x[038])))) | (x[036] & ((~x[038] & (x[040] ? (x[041] & x[042]) : ~x[042])) | (~x[041] & ((~x[040] & x[042]) | (x[038] & x[040] & ~x[042]))))))) | (~x[038] & ~x[039] & x[040] & x[041] & (x[036] ^ x[042])))) | (~x[039] & ((x[041] & (x[033] ? (x[036] ? (x[038] ? (x[040] ? (x[042] & ~x[043]) : ~x[042]) : (x[040] & ~x[043])) : (x[038] ? x[040] : (~x[040] & x[042]))) : ((x[038] & (x[036] ? (~x[040] & x[042]) : (x[040] & ~x[042]))) | (~x[036] & x[040] & ~x[043] & (x[042] | (~x[038] & ~x[042])))))) | (~x[041] & ((~x[036] & (x[033] ? ((x[038] & x[042]) | (~x[040] & ~x[042] & ~x[043])) : ((~x[040] & ~x[042]) | (~x[043] & (x[040] ? (x[038] | (~x[038] & x[042])) : x[042]))))) | (~x[043] & ((~x[038] & x[040] & ~x[042]) | (x[036] & (x[038] ? (x[040] & x[042]) : (~x[040] & ~x[042]))))))) | (x[036] & ~x[043] & ((~x[033] & (x[038] ? ~x[042] : (~x[040] & x[042]))) | (~x[040] & x[042] & x[033] & x[038]))))) | (~x[043] & ((x[039] & ((x[033] & ((~x[041] & ((x[042] & (x[036] ? (~x[040] | (x[038] & x[040])) : (~x[038] & ~x[040]))) | (~x[040] & (x[038] ? ~x[036] : ~x[042])))) | (x[036] & x[040] & (~x[042] | (~x[038] & x[041] & x[042]))) | (~x[036] & x[041] & x[042]))) | (x[040] & ((~x[033] & (x[036] ? (x[038] & x[041]) : ~x[038])) | (~x[041] & x[042] & x[036] & ~x[038]))) | (~x[033] & ~x[040] & ((~x[038] & x[041] & x[042]) | (~x[036] & (x[042] ? x[038] : ~x[041])))))) | (x[036] & ~x[038] & x[041] & ((~x[040] & (~x[042] | (x[033] & x[042]))) | (~x[033] & x[040] & ~x[042]))))) | (~x[036] & x[039] & x[040] & ~x[042] & (x[033] ? (~x[038] & x[041]) : (x[038] & ~x[041]))))) | (~x[035] & ((~x[033] & ((x[036] & ((x[042] & ((~x[038] & (x[039] ? ~x[043] : (~x[040] & x[041]))) | (~x[039] & ((x[040] & ~x[041] & x[043]) | (x[038] & ~x[043] & (x[040] ^ x[041])))) | (~x[040] & ~x[041] & x[038] & x[039]))) | (~x[043] & ((x[039] & ((x[038] & x[041]) | (~x[040] & ~x[041] & ~x[042]))) | (~x[039] & ~x[040] & ~x[041]) | (x[038] & x[040] & (x[041] ? ~x[039] : ~x[042])))) | (x[041] & ~x[042] & x[043] & x[038] & x[039]))) | (~x[038] & x[040] & x[041] & x[042] & x[043]) | (~x[036] & ((x[039] & ((x[038] & (x[040] ? (x[042] & ~x[043]) : x[041])) | (~x[040] & ~x[041] & ~x[042] & x[043]) | (x[041] & ~x[043] & (x[042] ? ~x[038] : x[040])))) | (~x[042] & ((~x[038] & x[040] & ~x[041]) | (~x[039] & ((x[038] & (~x[043] | (~x[041] & x[043]))) | (~x[038] & (x[043] ? ~x[040] : x[041])) | (x[040] & x[041] & x[043]))))) | (~x[039] & x[042] & (x[038] | (~x[038] & ~x[040] & ~x[041]))))))) | (x[033] & ((x[038] & ((~x[042] & (x[036] ? (x[039] ? x[040] : (x[041] & ~x[043])) : ((x[040] & x[043]) | (x[039] & ~x[041] & (~x[043] | (~x[040] & x[043])))))) | (~x[036] & ((~x[043] & (x[039] ? (x[040] ? (~x[041] & x[042]) : x[041]) : (x[041] ? x[042] : ~x[040]))) | (x[042] & x[043] & (x[041] ? x[040] : ~x[039])))) | (x[039] & ((x[040] & x[041] & x[042] & ~x[043]) | (~x[040] & (x[041] ? x[043] : (x[042] & ~x[043]))))))) | (~x[040] & ((x[042] & ((x[036] & (x[039] ? (~x[041] & x[043]) : (x[041] & ~x[043]))) | (x[041] & ((~x[036] & ~x[039] & x[043]) | (~x[038] & x[039] & ~x[043]))))) | (~x[036] & ((~x[041] & ((~x[038] & (x[039] ? x[043] : (~x[042] & ~x[043]))) | (~x[039] & ~x[042] & x[043]))) | (x[041] & ~x[042] & ~x[038] & ~x[039]))) | (~x[042] & ~x[043] & x[036] & ~x[038]))) | (~x[039] & ((~x[038] & (x[036] ? (x[043] & (~x[041] | (x[040] & x[041] & ~x[042]))) : (x[040] & (x[041] ? (x[042] & ~x[043]) : ~x[042])))) | (x[040] & x[041] & (x[036] ? x[042] : (~x[042] & ~x[043]))))) | (x[040] & ~x[041] & ~x[038] & x[039]))) | (x[036] & ((~x[042] & (x[038] ? (x[043] & (x[039] ? (~x[040] & ~x[041]) : (x[040] & x[041]))) : (x[040] & ~x[043] & (~x[039] ^ x[041])))) | (x[038] & ~x[039] & ~x[040] & x[041] & x[043]))) | (~x[036] & ~x[040] & ((~x[038] & ((x[039] & (x[041] ? (~x[042] & x[043]) : (x[042] & ~x[043]))) | (x[042] & ~x[043] & ~x[039] & x[041]))) | (~x[041] & x[042] & x[043] & x[038] & x[039]))))) | (~x[039] & ((~x[041] & (x[033] ? (x[036] ? (x[038] ? (~x[040] & ~x[042]) : (x[042] & ~x[043])) : ((~x[038] & x[042]) | (x[038] & x[040] & ~x[042] & ~x[043]))) : (x[036] & ((~x[038] & ((~x[042] & x[043]) | (x[040] & x[042] & ~x[043]))) | (x[038] & ~x[040] & ~x[042] & x[043]))))) | (~x[036] & ~x[040] & x[041] & (x[033] ? (x[038] & ~x[042]) : (x[043] & (~x[038] ^ ~x[042])))))) | (x[039] & ((x[038] & ((x[033] & ((~x[043] & ((x[036] & ~x[040] & (~x[042] | (x[041] & x[042]))) | (x[041] & ~x[042] & ~x[036] & x[040]))) | (x[040] & ~x[041] & x[042] & x[043]))) | (x[040] & ~x[041] & x[042] & ~x[033] & x[036]))) | (~x[033] & x[041] & x[043] & ((~x[038] & x[040] & ~x[042]) | (x[036] & ~x[040] & x[042]))))) | (~x[033] & x[036] & x[038] & x[040] & ~x[041] & ~x[042] & x[043]))) | (x[037] & ((~x[040] & ((x[035] & ((~x[038] & ((x[039] & ((x[033] & ((x[041] & x[042]) | (x[036] & ~x[041] & ~x[043]))) | (x[036] & (x[041] ? (~x[042] & ~x[043]) : (x[042] & x[043]))))) | (~x[033] & ((~x[036] & ((x[041] & x[042] & x[043]) | (~x[039] & ~x[042]))) | (~x[039] & ((x[041] & x[042] & ~x[043]) | (x[036] & ~x[041] & x[043]))) | (x[036] & ~x[042] & (x[041] ^ ~x[043])))))) | (~x[043] & ((x[038] & ((~x[036] & ((x[033] & ~x[041] & (x[039] ^ ~x[042])) | (x[039] & x[041] & x[042]))) | (~x[033] & ((x[036] & x[042]) | (~x[039] & x[041] & ~x[042]))))) | (x[033] & ((x[036] & ~x[039] & (~x[041] | (x[041] & ~x[042]))) | (~x[041] & ~x[042] & ~x[036] & x[039]))))) | (x[043] & ((~x[033] & (x[036] ? ((x[038] & x[041] & x[042]) | (x[039] & ~x[041] & ~x[042])) : ((x[039] & x[041] & ~x[042]) | (x[038] & ~x[039] & ~x[041])))) | (x[038] & ((~x[039] & (x[036] ? (~x[041] & x[042]) : (x[041] & ~x[042]))) | (~x[036] & x[042] & (x[041] ? x[033] : x[039])))))))) | (~x[035] & ((x[036] & (x[033] ? ((x[042] & (x[038] ? (x[039] ? ~x[041] : x[043]) : (x[039] ? (~x[041] & x[043]) : (x[041] & ~x[043])))) | (~x[043] & (x[038] ? (x[039] ? ~x[042] : x[041]) : (x[041] ? ~x[042] : (~x[039] | (x[039] & ~x[042])))))) : ((x[042] & (x[038] ? x[041] : (x[039] & ~x[041]))) | (x[038] & ~x[041] & (x[043] ? ~x[039] : ~x[042]))))) | (~x[036] & ((x[042] & ((~x[033] & x[038] & ~x[039] & x[041]) | (x[039] & ~x[041] & x[033] & ~x[038]))) | (~x[042] & (x[033] ? ((x[039] & x[041]) | (~x[038] & ((~x[041] & x[043]) | (~x[039] & x[041] & ~x[043])))) : (x[038] ? (~x[039] | (x[039] & ~x[041] & x[043])) : (x[039] & x[043])))) | (x[039] & ~x[041] & ~x[043] & x[033] & x[038]))) | (x[041] & ((~x[038] & ((x[039] & x[042]) | (~x[033] & ~x[039] & ~x[043]))) | (x[033] & x[038] & x[039] & x[042] & ~x[043]))))) | (x[043] & ((x[036] & ((~x[033] & x[038] & (x[039] ? (~x[041] & x[042]) : (x[041] & ~x[042]))) | (~x[039] & ((~x[038] & x[041] & x[042]) | (x[033] & ~x[041] & ~x[042]))))) | (x[033] & ~x[036] & ((~x[038] & ~x[039] & x[041]) | (~x[041] & ~x[042] & x[038] & x[039]))))) | (~x[039] & x[042] & ((x[033] & ~x[036] & (~x[041] | (~x[038] & x[041] & ~x[043]))) | (~x[033] & x[036] & ~x[038] & ~x[041] & ~x[043]))))) | (x[040] & ((x[035] & ((~x[033] & ((x[041] & (x[036] ? (x[038] ? (~x[042] & (~x[039] | (x[039] & x[043]))) : (~x[039] & x[042])) : ((~x[042] & ~x[043]) | (x[038] & x[039] & x[043])))) | (~x[041] & ((x[036] & ((x[038] & x[039] & x[043]) | (~x[039] & x[042] & ~x[043]))) | (~x[038] & x[039] & x[042]) | (~x[042] & x[043] & x[038] & ~x[039]))) | (x[036] & ~x[038] & ~x[042] & (x[039] | (~x[039] & ~x[043]))) | (x[042] & ~x[043] & x[038] & x[039]))) | (x[033] & ((~x[038] & ((x[036] & (x[039] ? ~x[043] : ~x[042])) | (x[039] & (x[041] ? ~x[036] : (x[042] & x[043]))))) | (~x[036] & ((x[038] & (x[039] ? (x[041] ? ~x[043] : (x[042] & x[043])) : (~x[042] | (x[041] & x[042])))) | (x[042] & x[043] & ~x[039] & ~x[041]))) | (x[038] & ~x[039] & ~x[041] & x[042] & ~x[043]))) | (x[036] & x[038] & ~x[039] & ~x[041] & ~x[042] & ~x[043]))) | (~x[035] & ((x[039] & ((x[036] & (x[033] ? ((x[038] & (x[043] ? x[042] : x[041])) | (~x[043] & ((~x[041] & x[042]) | (~x[038] & x[041] & ~x[042])))) : ((~x[041] & (x[042] | (~x[042] & ~x[043]))) | (x[042] & x[043] & ~x[038] & x[041])))) | (x[033] & ((x[041] & ((x[038] & ~x[042] & x[043]) | (~x[036] & ~x[038] & x[042]))) | (~x[041] & ~x[042] & ~x[043]) | (~x[036] & x[038] & (x[043] ? ~x[041] : x[042])))) | (~x[038] & ~x[041] & x[043] & (~x[042] | (~x[036] & x[042]))))) | (~x[039] & ((x[033] & ((x[036] & (x[038] ? (x[041] & x[042]) : (~x[041] & ~x[042]))) | (~x[036] & ~x[038] & (~x[041] ^ ~x[043])) | (x[038] & ~x[041] & x[042] & x[043]))) | (x[036] & ((~x[033] & (x[038] ? (~x[041] & ~x[042]) : (x[041] & x[043]))) | (x[038] & x[041] & ~x[042] & ~x[043]))) | (~x[033] & ~x[038] & x[041] & ~x[042] & ~x[043]))) | (x[041] & x[042] & ~x[043] & x[033] & x[036] & ~x[038]))) | (~x[038] & (x[033] ? ((x[036] & (x[039] ? (x[041] & x[043]) : (~x[041] & x[042]))) | (~x[039] & x[042] & ((x[041] & x[043]) | (~x[036] & ~x[041] & ~x[043])))) : (~x[036] & (x[039] ? (x[041] & (x[042] | (~x[042] & x[043]))) : (~x[042] & x[043]))))))) | (~x[042] & (x[038] ? ((x[036] & ((x[039] & ((~x[033] & x[041] & (~x[035] | (x[035] & ~x[043]))) | (~x[035] & ~x[041] & x[043]))) | (x[033] & ~x[035] & ~x[039] & x[041] & x[043]))) | (x[033] & ~x[036] & ((~x[035] & ~x[039]) | (x[041] & x[043] & x[035] & x[039])))) : (~x[041] & (x[035] ? (x[033] ? (x[036] ? (x[039] & x[043]) : ~x[039]) : (~x[036] & x[039])) : (~x[043] & ((~x[036] & ~x[039]) | (~x[033] & (x[036] ^ x[039])))))))) | (x[042] & ((x[041] & ((~x[038] & ((~x[033] & ((x[035] & x[036] & x[039]) | (~x[035] & ~x[036] & ~x[039] & x[043]))) | (x[033] & x[035] & x[036] & ~x[039] & ~x[043]))) | (x[033] & x[038] & (x[035] ? (x[036] & ~x[039]) : (~x[036] & (~x[039] | (x[039] & x[043]))))))) | (~x[033] & ~x[036] & x[038] & ~x[041] & ~x[043] & (~x[035] | (x[035] & ~x[039]))))))) | (~x[036] & ((x[035] & ((x[041] & ((~x[033] & ((x[040] & x[042] & x[043] & x[038] & ~x[039]) | (~x[038] & x[039] & ~x[040] & ~x[042] & ~x[043]))) | (~x[043] & ((x[033] & ~x[038] & ((~x[040] & ~x[042]) | (~x[039] & x[040] & x[042]))) | (x[038] & ~x[040] & (x[039] ^ x[042])))) | (x[033] & ~x[038] & ~x[039] & x[040] & ~x[042]))) | (x[033] & ~x[041] & ((~x[042] & (x[038] ? (x[039] ? (x[040] & ~x[043]) : (~x[040] & x[043])) : (x[039] & x[040]))) | (x[042] & ~x[043] & x[039] & x[040]))))) | (~x[038] & ((x[033] & ~x[035] & ~x[042] & ((x[040] & x[041] & x[043]) | (~x[041] & ~x[043] & x[039] & ~x[040]))) | (~x[041] & x[042] & x[043] & ~x[033] & x[039] & ~x[040]))) | (x[040] & ~x[041] & x[042] & ~x[043] & x[033] & ~x[035] & x[038] & ~x[039]))) | (x[036] & ((~x[042] & ((x[038] & ((~x[039] & ((x[033] & x[040] & (~x[035] ^ x[041])) | (~x[033] & ~x[035] & ~x[040] & x[041] & ~x[043]))) | (~x[033] & x[035] & x[039] & x[040] & ~x[041] & ~x[043]))) | (~x[035] & ~x[038] & ((~x[040] & x[043] & (x[033] ? (x[039] | (~x[039] & x[041])) : (x[039] & x[041]))) | (x[040] & x[041] & ~x[043] & x[033] & ~x[039]))))) | (~x[035] & x[042] & ((~x[041] & ((x[033] & ~x[043] & (x[038] ? ~x[039] : (x[039] & ~x[040]))) | (~x[033] & ~x[038] & ~x[039] & ~x[040] & x[043]))) | (~x[033] & x[038] & x[040] & x[041] & x[043]))))) | (~x[033] & ~x[035] & ~x[038] & x[041] & ~x[043] & (x[039] ? (~x[040] & ~x[042]) : (x[040] & x[042]))))) | (~x[033] & ((~x[039] & ((x[032] & ((x[035] & (((~x[040] ^ x[041]) & ((x[042] & x[043] & ~x[036] & ~x[037]) | (~x[042] & ~x[043] & x[036] & x[038]))) | (x[043] & ((~x[037] & ((x[041] & ~x[042] & ~x[036] & x[038]) | (~x[041] & ((x[036] & (x[040] ? ~x[042] : ~x[038])) | (x[038] & ~x[040] & ~x[042]) | (~x[036] & x[040]))))) | (x[036] & ((x[037] & (x[038] ? (x[040] ^ x[042]) : (~x[040] & x[041]))) | (x[041] & x[042] & ~x[038] & x[040]))) | (~x[036] & ((x[037] & (x[038] ? (x[041] & x[042]) : (~x[041] & ~x[042]))) | (x[041] & x[042] & ~x[038] & ~x[040]))))) | (x[037] & ((~x[043] & ((~x[040] & ((x[038] & (x[041] ? ~x[036] : x[042])) | (x[041] & x[042] & x[036] & ~x[038]))) | (x[040] & (x[036] ? (x[041] ? ~x[038] : ~x[042]) : (x[038] & ~x[041]))) | (x[041] & ~x[042] & ~x[036] & ~x[038]))) | (x[036] & ~x[038] & ~x[041] & (~x[040] | (x[040] & x[042]))))) | (~x[037] & ~x[043] & ((~x[036] & (x[038] ? (x[040] & x[041]) : ~x[041])) | (x[038] & (x[040] ^ x[041])) | (x[036] & ~x[038] & x[040] & ~x[042]))))) | (~x[042] & ((~x[037] & ((x[040] & ((x[036] & ((~x[035] & ~x[038] & ~x[041]) | (x[038] & x[041] & x[043]))) | (~x[035] & ((~x[038] & x[041] & x[043]) | (~x[041] & (x[043] ? x[038] : ~x[036])))))) | (~x[036] & ((~x[040] & ((x[038] & ~x[041] & ~x[043]) | (~x[035] & x[043] & (x[038] | (~x[038] & x[041]))))) | (~x[035] & ((x[041] & ~x[043]) | (~x[038] & ~x[041] & x[043]))))))) | (x[037] & ((~x[035] & ((x[040] & (x[036] ? (~x[038] & ~x[043]) : (x[038] ? x[043] : x[041]))) | (~x[043] & ((~x[036] & x[038] & ~x[041]) | (~x[040] & (x[036] ? (~x[041] | (x[038] & x[041])) : x[041])))) | (x[036] & x[038] & ~x[041] & x[043]))) | (~x[036] & (x[038] ? (~x[040] & x[043]) : ((~x[041] & ~x[043]) | (~x[040] & x[041] & x[043])))))) | (x[036] & x[038] & ~x[040] & x[041] & x[043]))) | (~x[035] & ((x[042] & ((~x[038] & ((x[036] & ~x[037] & x[041]) | (~x[036] & ~x[040] & ~x[041] & x[043]))) | (x[036] & ((~x[041] & ((x[037] & (x[040] | (~x[040] & x[043]))) | (~x[040] & ~x[043] & ~x[037] & x[038]))) | (~x[037] & x[038] & x[043] & (~x[040] | (x[040] & x[041]))))) | (~x[036] & ((~x[037] & ~x[043] & ((~x[040] & ~x[041]) | (x[038] & x[040] & x[041]))) | (x[041] & x[043]) | (~x[040] & ~x[041] & x[037] & x[038]))))) | (x[036] & x[038] & ((~x[037] & ~x[043] & (x[040] | (~x[040] & x[041]))) | (x[041] & x[043] & x[037] & x[040]))))) | (x[036] & x[042] & ((x[040] & ~x[041] & ~x[037] & ~x[038]) | (~x[040] & x[041] & ~x[043] & x[037] & x[038]))))) | (x[035] & (x[042] ? ((~x[043] & (x[036] ? (~x[037] & (x[038] ? (~x[040] & ~x[041]) : (x[040] & x[041]))) : (x[037] & (x[038] ? (x[040] & x[041]) : (x[040] | (~x[040] & ~x[041])))))) | (x[040] & (x[036] ? (x[038] & (x[041] | (~x[041] & x[043]))) : (x[037] & x[043] & (~x[041] | (~x[038] & x[041])))))) : ((x[037] & ((~x[040] & ((x[036] & (x[038] ? (~x[041] & x[043]) : (x[041] & ~x[043]))) | (~x[041] & ~x[043] & ~x[036] & x[038]))) | (~x[036] & x[038] & x[040] & x[041] & x[043]))) | (~x[040] & x[041] & ~x[043] & ~x[036] & ~x[037] & ~x[038])))) | (~x[035] & ((x[037] & ((~x[038] & ~x[040] & ~x[041] & ~x[042] & x[043]) | (x[041] & x[042] & ~x[043] & x[036] & x[038] & x[040]))) | (~x[038] & ((x[036] & x[041] & ~x[042] & (x[043] ? ~x[040] : ~x[037])) | (~x[036] & x[040] & ~x[041] & x[042] & ~x[043]))))) | (x[036] & x[037] & ~x[038] & x[040] & ~x[041] & ~x[042] & x[043]))) | (x[032] & ((~x[035] & ((x[041] & ((~x[036] & ((~x[037] & ~x[038] & x[039] & ~x[042]) | (~x[040] & x[042] & ~x[043]))) | (x[039] & (x[037] ? (x[038] ? ((~x[040] & ~x[042]) | (x[036] & (x[042] ? ~x[043] : x[040]))) : ((x[040] & x[042] & ~x[043]) | (x[036] & ~x[040] & x[043]))) : ((x[036] & (x[040] ? (~x[042] & x[043]) : (x[043] ? x[038] : x[042]))) | (x[040] & ((x[042] & ~x[043]) | (x[038] & (x[042] ^ ~x[043]))))))) | (x[036] & x[037] & ((~x[038] & (x[040] ? (~x[042] & x[043]) : ~x[043])) | (x[038] & ~x[040] & x[042] & x[043]))))) | (~x[041] & ((x[036] & ((~x[040] & ((~x[038] & x[042] & ~x[043]) | (x[037] & x[038] & x[039] & ~x[042] & x[043]))) | (x[039] & ((x[040] & ((~x[043] & ((~x[037] & (~x[038] ^ ~x[042])) | (~x[038] & ~x[042]) | (x[037] & x[038] & x[042]))) | (x[037] & ~x[038] & (x[042] | (~x[042] & x[043]))))) | (~x[037] & x[038] & x[042]))) | (x[037] & x[038] & x[040] & ~x[042] & ~x[043]))) | (x[039] & ((~x[036] & ((x[042] & (x[037] ? (~x[038] & ~x[040]) : (~x[043] & (~x[038] | (x[038] & x[040]))))) | (~x[037] & ~x[040] & x[043]) | (x[037] & x[038] & (x[040] ? (~x[043] | (~x[042] & x[043])) : x[043])))) | (~x[042] & ((x[040] & x[043] & ~x[037] & ~x[038]) | (~x[040] & ~x[043] & x[037] & x[038]))))) | (~x[036] & x[040] & x[043] & (x[037] ? ~x[038] : (x[038] & x[042]))))) | (x[039] & ((~x[037] & ((~x[038] & ((x[036] & (x[042] ? x[043] : ~x[040])) | (x[042] & x[043] & ~x[036] & x[040]))) | (~x[036] & x[038] & ~x[040] & ~x[042] & ~x[043]))) | (~x[036] & x[037] & ((~x[038] & ~x[040] & ~x[042] & ~x[043]) | (x[038] & x[040] & x[042] & x[043]))))))) | (x[035] & ((x[039] & ((~x[043] & ((~x[036] & ((x[038] & (~x[040] | (x[041] & ~x[042] & ~x[037] & x[040]))) | (~x[041] & (x[037] ? (x[040] | (~x[038] & ~x[040] & ~x[042])) : (x[040] ? x[042] : ~x[038]))) | (x[040] & x[041] & x[042] & x[037] & ~x[038]))) | (x[036] & ((~x[038] & x[041] & x[042]) | (~x[041] & ((~x[037] & (~x[038] ^ x[042])) | (x[037] & ~x[040] & ~x[042]) | (~x[038] & x[040] & x[042]))))) | (x[037] & x[041] & (x[038] ? (x[040] & x[042]) : (~x[040] & ~x[042]))))) | (x[038] & ((~x[041] & (x[036] ? ((x[042] & x[043]) | (x[037] & x[040] & ~x[042])) : (~x[040] & x[043] & (x[037] ^ x[042])))) | (x[041] & ((~x[036] & (x[037] ? (~x[040] & x[043]) : (x[040] & x[042]))) | (x[036] & ~x[040] & x[042] & x[043]))) | (~x[042] & x[043] & ~x[037] & x[040]))) | (~x[038] & ((x[043] & ((~x[036] & ((~x[037] & ~x[040] & x[042]) | (~x[041] & ~x[042] & x[037] & x[040]))) | (x[037] & ((~x[040] & ~x[041] & x[042]) | (x[036] & x[040] & ~x[042]))) | (x[040] & ~x[041] & x[042]) | (x[036] & ~x[040] & (~x[042] | (~x[037] & x[041] & x[042]))))) | (x[036] & ~x[037] & ~x[040] & ~x[041] & x[042]))) | (x[041] & x[042] & x[043] & x[036] & ~x[037] & x[040]))) | (x[037] & ((x[038] & ((x[036] & ~x[043] & (x[040] ? (~x[041] & x[042]) : (x[041] & ~x[042]))) | (~x[036] & ~x[040] & ~x[041] & x[042] & x[043]))) | (x[041] & x[042] & ~x[043] & ~x[036] & ~x[038] & ~x[040]))) | (~x[037] & ~x[038] & ((x[041] & ((~x[036] & (x[042] ? ~x[043] : x[040])) | (x[036] & x[040] & ~x[042] & x[043]))) | (~x[036] & ~x[040] & ~x[042] & x[043]))))) | (x[039] & ((~x[042] & ((~x[043] & ((~x[037] & ((x[036] & (x[038] ? ~x[040] : (x[040] & x[041]))) | (x[040] & ~x[041] & ~x[036] & ~x[038]))) | (x[040] & x[041] & x[037] & ~x[038]))) | (~x[036] & x[037] & ((x[038] & x[040] & x[041]) | (~x[038] & ~x[040] & ~x[041] & x[043]))))) | (~x[036] & x[041] & x[043] & (x[037] ? ~x[038] : (x[038] & ~x[040]))))))) | (x[039] & (x[037] ? ((~x[041] & (x[035] ? ((x[040] & x[043] & ~x[036] & x[038]) | (x[036] & ~x[038] & ~x[040] & x[042] & ~x[043])) : (~x[038] & ((x[036] & ~x[040] & ~x[042]) | (x[042] & ~x[043] & ~x[036] & x[040]))))) | (x[035] & x[036] & x[038] & x[041] & x[043] & (x[040] ^ ~x[042]))) : ((~x[036] & ((x[040] & ((x[043] & ((x[035] & x[042] & (~x[038] ^ ~x[041])) | (x[041] & ~x[042] & ~x[035] & x[038]))) | (~x[041] & ~x[042] & ~x[035] & x[038]))) | (~x[035] & ~x[040] & x[042] & (x[038] ? (~x[041] & ~x[043]) : (x[041] & x[043]))))) | (x[035] & x[036] & x[038] & ~x[040] & x[041] & x[042] & ~x[043])))) | (~x[035] & ~x[040] & ~x[041] & ~x[043] & ((x[038] & x[042] & x[036] & x[037]) | (~x[038] & ~x[042] & ~x[036] & ~x[037]))))))) | (~x[032] & ((x[036] & ((x[040] & (x[037] ? ((~x[035] & ((~x[038] & ((x[033] & x[043] & (x[039] ? (~x[041] & x[042]) : (x[041] & ~x[042]))) | (~x[041] & x[042] & ~x[043] & ~x[033] & ~x[039]))) | (~x[033] & x[038] & ((~x[039] & (x[041] ? (~x[042] & x[043]) : x[042])) | (x[042] & ~x[043] & x[039] & x[041]))))) | (~x[039] & ~x[041] & x[043] & (x[033] ? (x[035] & x[038]) : (~x[038] & x[042])))) : (x[033] ? ((x[038] & ((x[039] & ((~x[042] & x[043] & x[035] & x[041]) | (~x[035] & x[042] & (x[041] ^ ~x[043])))) | (x[035] & ~x[039] & (x[041] ? (x[042] & x[043]) : (~x[042] & ~x[043]))))) | (~x[041] & ~x[042] & x[043] & x[035] & ~x[038] & ~x[039])) : ((x[039] & ((x[035] & x[041] & (x[038] ? x[043] : (x[042] & ~x[043]))) | (~x[038] & ~x[041] & (~x[042] | (~x[035] & x[042] & x[043]))))) | (x[041] & ~x[042] & x[043] & ~x[035] & ~x[038] & ~x[039]))))) | (~x[040] & ((x[043] & ((~x[035] & (x[033] ? (x[041] & ((x[037] & x[038] & x[039]) | (~x[037] & ~x[038] & ~x[039] & x[042]))) : (~x[037] & ~x[041] & (x[038] ? (~x[039] & x[042]) : x[039])))) | (x[035] & x[041] & ~x[042] & ((x[033] & x[037] & (~x[038] | (x[038] & ~x[039]))) | (x[038] & ~x[039] & ~x[033] & ~x[037]))) | (~x[039] & ~x[041] & x[042] & x[033] & x[037] & ~x[038]))) | (x[038] & ((~x[041] & ~x[043] & ((~x[033] & x[035] & (x[037] ? ~x[042] : (x[039] & x[042]))) | (x[033] & ~x[035] & x[037] & ~x[039] & ~x[042]))) | (~x[033] & x[035] & ~x[037] & x[039] & ~x[042]))) | (~x[037] & ~x[038] & ~x[033] & x[035] & ~x[042] & ~x[043] & x[039] & ~x[041]))) | (x[042] & x[043] & ~x[039] & ~x[041] & ~x[037] & x[038] & x[033] & ~x[035]))) | (~x[036] & (x[035] ? ((x[039] & ((x[043] & ((~x[037] & x[041] & ((~x[033] & ~x[040] & (~x[038] ^ ~x[042])) | (x[040] & x[042] & x[033] & ~x[038]))) | (x[033] & ~x[042] & ((x[037] & ~x[038] & ~x[040]) | (x[038] & x[040] & ~x[041]))))) | (x[037] & ((~x[033] & ~x[043] & ((x[041] & x[042] & ~x[038] & ~x[040]) | (x[038] & ~x[041] & (~x[042] | (~x[040] & x[042]))))) | (x[033] & ~x[038] & ~x[040] & ~x[041] & x[042]))) | (x[040] & ~x[041] & x[042] & ~x[043] & ~x[033] & ~x[037] & x[038]))) | (~x[039] & ((~x[040] & x[041] & ((x[038] & ((x[033] & (x[037] ? (~x[042] & ~x[043]) : (x[042] & x[043]))) | (~x[042] & ~x[043] & ~x[033] & ~x[037]))) | (~x[038] & x[042] & ~x[043] & ~x[033] & ~x[037]))) | (~x[033] & x[040] & ~x[041] & ((x[037] & ~x[042] & ~x[043]) | (x[042] & x[043] & ~x[037] & ~x[038]))))) | (x[041] & x[042] & x[043] & ~x[033] & x[038] & ~x[040])) : ((~x[038] & (x[037] ? ((~x[043] & ((x[039] & x[040] & ((x[041] & ~x[042]) | (x[033] & ~x[041] & x[042]))) | (~x[041] & x[042] & ~x[033] & ~x[040]))) | (~x[033] & ~x[039] & x[043] & ((~x[041] & x[042]) | (~x[040] & x[041] & ~x[042])))) : ((x[040] & ((x[033] & x[041] & (x[043] ? x[042] : x[039])) | (~x[041] & x[042] & ~x[043] & ~x[033] & x[039]))) | (x[041] & ~x[042] & ~x[043] & x[033] & x[039] & ~x[040])))) | (x[039] & ((x[038] & ((x[033] & x[037] & ((~x[040] & ~x[041] & x[042] & x[043]) | (x[040] & x[041] & ~x[042] & ~x[043]))) | (~x[041] & ~x[042] & ~x[043] & ~x[033] & ~x[037] & ~x[040]))) | (~x[041] & x[042] & x[043] & ~x[033] & ~x[037] & x[040])))))) | (~x[037] & ~x[038] & x[039] & ~x[040] & x[042] & ((x[041] & x[043] & x[033] & ~x[035]) | (~x[041] & ~x[043] & ~x[033] & x[035]))))) | (~x[033] & ((~x[041] & ((x[032] & ((~x[035] & (x[036] ? ((x[043] & ((x[042] & (~x[038] ^ x[040]) & (x[037] ^ ~x[039])) | (~x[037] & x[038] & x[039] & x[040] & ~x[042]))) | (~x[040] & ~x[042] & ~x[037] & ~x[039])) : ((x[037] & ((x[042] & ((x[038] & (x[039] ? (~x[040] & ~x[043]) : (x[040] & x[043]))) | (~x[040] & ~x[043] & ~x[038] & ~x[039]))) | (x[040] & ~x[042] & ~x[043] & ~x[038] & x[039]))) | (x[038] & ~x[039] & x[042] & ((x[040] & ~x[043]) | (~x[037] & ~x[040] & x[043])))))) | (x[035] & (x[038] ? (x[040] ? (~x[042] & ((~x[036] & x[037] & ~x[039] & x[043]) | (~x[037] & x[039] & ~x[043]))) : ((x[036] & x[043] & (x[037] ? (x[039] & ~x[042]) : (~x[039] & x[042]))) | (~x[036] & ~x[037] & ~x[039] & x[042] & ~x[043]))) : ((x[036] & ~x[043] & ((~x[037] & ~x[039] & ~x[040]) | (x[040] & ~x[042] & x[037] & x[039]))) | (~x[037] & x[039] & x[040] & ~x[042] & x[043])))) | (x[036] & ~x[037] & x[038] & ~x[042] & x[043] & x[039] & ~x[040]))) | (~x[036] & ((x[035] & ~x[040] & ((x[037] & ~x[038] & x[042] & (x[039] ^ x[043])) | (~x[037] & x[038] & x[039] & ~x[042] & x[043]))) | (~x[035] & ~x[037] & ~x[038] & x[042] & x[043] & ~x[039] & x[040]))))) | (x[032] & ((x[041] & (x[037] ? (x[035] ? ((x[036] & x[039] & (x[038] ? (x[040] & ~x[042]) : (x[042] & x[043]))) | (~x[039] & x[040] & ~x[042] & ((~x[038] & x[043]) | (~x[036] & x[038] & ~x[043])))) : ((x[042] & ((~x[036] & ((x[038] & x[039] & (~x[040] ^ ~x[043])) | (~x[039] & x[040] & ~x[043]))) | (x[036] & ~x[038] & ~x[039] & x[040]))) | (x[040] & ~x[042] & ~x[043] & x[038] & ~x[039]))) : ((~x[042] & ((~x[036] & ((~x[035] & x[038] & ~x[039] & x[040] & x[043]) | (x[039] & ~x[040] & ~x[043] & x[035] & ~x[038]))) | (x[035] & x[036] & ~x[040] & (x[038] ? (x[039] & x[043]) : (~x[043] | (~x[039] & x[043])))))) | (x[035] & ((x[036] & ((~x[040] & x[042] & ~x[038] & ~x[039]) | (x[040] & ~x[043] & x[038] & x[039]))) | (x[038] & ~x[039] & ~x[040] & x[042] & x[043])))))) | (x[035] & x[036] & x[037] & x[038] & x[042] & ~x[043] & x[039] & ~x[040])))))) & ((~x[003] & ~x[007] & ((x[000] & ~x[006] & ~x[009] & ((~x[001] & x[002] & x[004] & x[005] & ~x[008] & ~x[010] & x[011]) | (x[001] & ~x[002] & ~x[004] & ~x[005] & x[008] & x[010] & ~x[011] & x[012] & ~x[013] & ~x[014] & ~x[015]))) | (~x[000] & ~x[001] & ~x[002] & x[004] & ~x[005] & x[006]))) | (~x[112] & ~x[113] & ~x[114] & ~x[116] & ((~x[069] & ((~x[076] & ((~x[071] & ((~x[067] & ((x[065] & ~x[075] & x[078] & ((x[064] & ~x[066] & ~x[068] & ~x[070] & x[072] & x[073] & ~x[074] & x[077] & ~x[079] & x[115] & ~x[117] & ~x[118] & x[119]) | (~x[064] & x[066] & x[068] & x[070] & ~x[072] & ~x[073] & x[074] & ~x[077] & x[079] & ~x[115] & x[117] & x[118] & ~x[119]))) | (~x[064] & ~x[065] & ~x[066] & ~x[068] & ~x[070] & ~x[072] & x[075] & ((~x[078] & ((x[115] & ~x[117] & ~x[118] & x[119] & (x[073] ? (~x[077] & (~x[074] | (x[074] & x[079]))) : (x[077] & x[079]))) | (~x[115] & x[117] & x[118] & ~x[119] & x[077] & x[079] & ~x[073] & x[074]))) | (x[115] & ~x[117] & ~x[118] & x[119] & x[077] & ~x[079] & ~x[073] & ~x[074]))))) | (~x[064] & ~x[065] & ~x[066] & x[067] & ~x[068] & x[070] & ~x[072] & ~x[073] & x[074] & x[075] & x[077] & x[115] & ~x[117] & ~x[118] & x[119] & (x[078] ^ x[079])))) | (~x[064] & ~x[065] & ~x[066] & x[067] & ~x[068] & x[070] & x[071] & x[072] & x[073] & ~x[074] & ~x[075] & x[077] & ~x[078] & ~x[079] & ~x[096] & ~x[097] & ~x[098] & ~x[099] & x[100] & ~x[101] & ~x[102] & ~x[103] & ~x[104] & ~x[105] & ~x[106] & ~x[107] & ~x[108] & ~x[109] & ~x[110] & ~x[111] & ((x[115] & ~x[117] & ~x[118] & x[119]) | (~x[115] & x[117] & x[118] & ~x[119]))))) | (~x[064] & ~x[065] & ~x[066] & ~x[068] & x[075] & x[076] & ~x[077] & ((x[067] & x[070] & ~x[078] & ~x[115] & x[117] & x[118] & ~x[119] & ((~x[071] & ~x[072] & ~x[073] & x[074] & x[079]) | (x[071] & x[072] & x[073] & ~x[074] & ~x[079] & ~x[096] & ~x[097] & ~x[098] & ~x[099] & x[100] & ~x[101] & ~x[102] & ~x[103] & ~x[104] & ~x[105] & ~x[106] & ~x[107] & ~x[108] & ~x[109] & ~x[110] & ~x[111]))) | (~x[067] & ~x[070] & x[071] & x[072] & ~x[073] & x[074] & x[078] & x[079] & x[115] & ~x[117] & ~x[118] & x[119]))))) | (~x[085] & ((~x[092] & ((~x[087] & ((~x[083] & ((x[081] & ~x[091] & x[094] & ((x[080] & ~x[082] & ~x[084] & ~x[086] & x[088] & x[089] & x[115] & ~x[117] & ~x[118] & x[119] & ~x[090] & x[093] & ~x[095]) | (~x[080] & x[082] & x[084] & x[086] & ~x[088] & ~x[089] & ~x[115] & x[117] & x[118] & ~x[119] & x[090] & ~x[093] & x[095]))) | (~x[080] & ~x[081] & ~x[082] & ~x[084] & ~x[086] & ~x[088] & x[091] & ((~x[094] & ((x[115] & ~x[117] & ~x[118] & x[119] & (x[089] ? (~x[093] & (~x[090] | (x[090] & x[095]))) : (x[093] & x[095]))) | (~x[115] & x[117] & x[118] & ~x[119] & x[093] & x[095] & ~x[089] & x[090]))) | (x[115] & ~x[117] & ~x[118] & x[119] & x[093] & ~x[095] & ~x[089] & ~x[090]))))) | (~x[080] & ~x[081] & ~x[082] & x[083] & ~x[084] & x[086] & ~x[088] & ~x[089] & x[090] & x[091] & x[093] & x[115] & ~x[117] & ~x[118] & x[119] & (x[094] ^ x[095])))) | (~x[080] & ~x[081] & ~x[082] & x[083] & ~x[084] & x[086] & x[087] & x[088] & x[089] & ~x[090] & ~x[091] & x[093] & ~x[094] & ~x[095] & ~x[096] & ~x[097] & ~x[098] & ~x[099] & x[100] & ~x[101] & ~x[102] & ~x[103] & ~x[104] & ~x[105] & ~x[106] & ~x[107] & ~x[108] & ~x[109] & ~x[110] & ~x[111] & ((x[115] & ~x[117] & ~x[118] & x[119]) | (~x[115] & x[117] & x[118] & ~x[119]))))) | (~x[080] & ~x[081] & ~x[082] & ~x[084] & x[091] & x[092] & ~x[093] & ((x[083] & x[086] & ~x[094] & ~x[115] & x[117] & x[118] & ~x[119] & ((~x[087] & ~x[088] & ~x[089] & x[090] & x[095]) | (~x[101] & ~x[102] & ~x[103] & ~x[104] & ~x[105] & ~x[106] & ~x[107] & ~x[108] & ~x[109] & ~x[110] & ~x[111] & ~x[096] & ~x[097] & ~x[098] & ~x[099] & x[100] & x[087] & x[088] & x[089] & ~x[090] & ~x[095]))) | (~x[083] & ~x[086] & x[087] & x[088] & ~x[089] & x[090] & ~x[117] & ~x[118] & x[119] & x[094] & x[095] & x[115]))))))));
  
  assign xin_ready = (z0_ready || ~z0_valid);
  
  initial begin
	z0_valid = 0;
	x_valid <= 0;
  end
endmodule


