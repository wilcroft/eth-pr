// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:12 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cR7thPlkvhWvwBXIRcNrJ3/wtsUGMAZh9DxDZYvlkAHlr2d36GAGeiUGoDIQg/88
BfNZXiLHtVQcjtVDgF1yoSJyV8J8vb3V9OJZVh0lMtlzEfBhuNf8o3us3pJolXDl
dW3l7RoxJVRlsPB+guI6PheC7HdmZU4UYgE6VU337MQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27776)
o3e7zNbM3wJFmHlydSLT6asMoU1kcBDMB0RlvhcwvP0q59tGekIObu3AX//FG+/U
ecscGOzEJB+Wv/sfXvOx/sYDlKYVGl1o8bggaFvACCaIPIaix36myX9Q9smfzB3d
WXJgKHEiN/7ZyHACMv9Tk7AR1CyffFkIc0MEBpl2NlyGfbLnsY4hrDlomdnwF9Vw
mhPs/Wk8Sc1nvfN5O7EXOH3O45X4KLopSZsLcR5PAtXI3lmIOvw5W/ryL93P1voN
nuQP8gjiSn9mNGtm73szutsEXxX2EbOzUMngAIyzWAFYvJHzzH8bmKrWCioH2Aap
aQdk1zeTIxn7WWE9OgwEvGDZfOatAnfYeCzwoCQyDGiIutzfNcdk88J+Nb9l5Vf3
00oYS6mq54cBMw5V6tfAjKqFZdJWtmuMYlKRPvxXjKaCdGOfTMMcvebhKJ9O4Ica
OBQT+TncuvNXMHL/WN5Q/TipraHUBIg8vmjR6krA9mEnk5hCw0ZDzLViiF0MSwHz
52IzDLU5txacB1y+Q+eM/gsfV/OPr/O4um4qJFzeGGoDl5ipS1S3SkJ7a1HKvgh4
gJDEH5pt+KCnGtyGRSJxOQP+XMJMDJnS0ofcM9372kcMwgXpOxZ4KQu8CW8h7THd
HkzpyTxEbwmM8ArVAu9z+vUdf9VMVs/WTrxsRIjjqHom8CD+8QEkn8Ian21OwtJz
cbXIGtKX71fnxnBwNnFkSlWjAn1Gui0O0utW9E1ZPDw0LQI8pfXoANS4z5J46AD6
lfmIYF+dISkGptDthUV6HzBz7F0SZkNa2VNd4o7jgkyR8nRaP3+GmcmVH3QK8DMF
n9+BrHEv3RjM9Xmvs1pLAswAkuS14fQ7w7wFn2zAGkEN6/4ZYRZ0DBuoQtGfAMIS
665qfPuFvJXdt5AqE6ilcXsO9x2GMVFLfeyBFr77Jx8mihu1IBZFWlOn6M/39tS1
vxRQ4TDal/MPDGoqkHHEOQc0M/uiblFBZrb7A1ETZUJlx1VFMwH0jsEJDT6xDlVO
c59TrulBSDFaD+kpcRwfaPyDEfib7Jw16sAVovr+K8A2ZzY2paQw74WRUhDUR0vn
YR6GsyK9Dp8kYGutKnTlAjbIUSWR8iB6t3dIPyqoUaaGgPJauEIbU4SbfvWR5xl3
bVb12aogXxx1A5OVWCLDB9xPeGGGksI8vlR7XMCNwSdFZ4scZAReo2x7OGnw5T+K
RvTC83CprPRemOYRcSQSToARj3P8q1TXTyxlCx256ZFiKphyOQzIaWKpQzN63UPF
+Gz57sslVrt4UA5I3MR/wmxYfm6crDyb6FPHupqz2yAreFzqZzEytXgDmuiGFlvq
b/b/ljVUX7NCH/MAg1O0OcgBZq6zPOTUNYFTDV1sxKejlL5wEnWBzIy7w6abRgwP
PHdURvM/zuS9271Ao63U6+c4R3BB6SNOa/xh5VGo9TGCtgmi4OVcG3FVqEqwpkGQ
5r1Vlf13plvOSFUoLOI7d3d4rTjGflmsyZYvdKHLXIfDoiYGmzqf8fDYAnOZ2cnz
+yeLK8A4EcJnWY5bR5Zpz7bsYfDa/kTKHUUc2UiD9lUBZWrArOsyZus2EcL5ZufJ
F87FArj2H8mfaILpgbsb4O0nP2qQD3YfXMA9p7lD8skG/koVM1D/kwZDv653L8bG
+SsSsoBy27KSdiEKDNFpLT/M67qACMTyHWq2lsXCCVLOQAvd670YPfXj3+zzl1aE
wRtA/mDH3/94MyKo76XLf53VOs0x1UwOTb6a/jhOXuoB5z4DvyrJtBxDdYFeFc4c
VfW/HemR6kbws/WuAvILCfw0nYXs3kVQJEZJKFjWipyFY3TgHa74LvY5z6jIPLVO
CSSW8djW//paWKKNFeoHtaWfwgene+w8eZ+hj/Ql33GpiJAQYThtlphE7UVLHRZY
gVhcdSlxVzbGrInuIsvJ2GSD3yOBjMWzJo4yHRD1Sj7bPQd+zE3WIhb5MQnOjBS+
T9fJs/N/NdxBs4Qmu97NNigvyVpgGMfVahHc9T2b940WZGHZmuFJTp5rfRHdTIBX
plv/1VgKZFvB7n9zW262I+Q0aY914YH10Vd66MibeeNoC78IS5vbTV41UF+/a7l/
Vid1HEpbpVUhCJyV0tpknc5rp4dnfOn0nxtHcj1tAP3F+qb3YErAuSGX0sgNYIWR
tFzKAA9R3aBEfs5vqboBycJmEGhRA3MdPgMHzoJn1sJ1iUhsnyhle+t/trugKoZf
RbPaQ22Aa9Gx5U6GcDrntkk4wqCSH3+ecUW54CE+4ImnamaIPYj121qffb8IlIzf
f1ySPlaeQ8qyz6rbodLKRL6blfvXSRfvXVuGuxJ4b/flXAnRW2P6SOL8H7kbBsNo
7tmuVPCUquUdptU3lXmpbhWSb445aJCu3MDsD2xPzA12W+YNw+Gxt3cI7w8LeAkC
PFGhMCoAsJidUJIpubdSB0pEhazBQM8k6H41d5s55eNq1vfK58tA1HGZidxfJ4bF
71thcWte34WZ0r98rtZ8nqb6xDzWzsU8yxQrf7tTaH4BBABQuoq+JTVAQoMwQrPL
Z5pk3nmKt+HTykVwun14V0PHWDeKokEFc5TrpjJ1iYkyWsnS4Ki/A7eyDKjb+Y+5
AWGRtzm2jLGSLaURQlNSCb3hcV1rxdc7bCV0v1ddtAkX53dzvYj14c898FG4U8+L
mVokbuIaaxvs9vYxuUh346RlNc3w2SATT5+pyPSiF4NqTCuFw9+wYOidXBpUuGT8
w5YEIqDo61siLzaT5uY4Qcibc5lZBEV+95YE0JM7loiRG6wR/s6E8msSmoARrorC
MpR93ysMX3jzTn8VkHVrSj9swxyN1KveUHX9gnsZ82gtS3IJTgatvHLp0wcTJqSw
kan98Benku0svSJhK0fAAx4O4HqAnVZRVIpBgoV/eSStHp4MZuyyOk+hMhwSLjMW
ZJV7QqjG40Vf76nM9evtMwymTmmB/Bsy0zI64dpJqqVunShmUA4/Iq+rLexoYcay
5gOPFtBW4u84X1rpd5t03iKQHW9WXntPgPta+XvTfPJ8wvIQnBQiP38cnBeqK3vh
ItHQkmJK+/Zmu6BqZv9USFEzlKkawht0VTpv8dhb65zm4c7JG8HXwlwty5JXj7Vp
CdECpzJDdjxkOQZ7oFbaG3KnanR3FYrQBj8aMNCKh6fUggSAWFtqIMSyGEAqlIbL
c/z0cUS7fWQAAIa8xogQCweLIbANKSFpupKzqi0u03bwBbP/6lJ7LgN2O5W852GH
xSqUI6heYfBLJl983F8OkdIu+IlpHvNaf3EAVkyiTRYGIFMaGjEg6TQRoCnwFw46
ePM1D3pV2abFC/gbMvaOa5fqpIOJMnFcQ1q9EbZw8g6eseAjyZn5fvJdSBPgZyLx
UcH4hMXmKI05DnH6tyyDqpXjCOo4TpWj+OWZrUkEIdi7359DzN9Aneya1fkwNVFY
3jt7cFJQ7b9fkuN6hYrp3tkuEsnIbrGAJzo6H6V5Zzwzx/vm/UvVxPJOAoSKpP5U
9TxN1qrg8nfbPYKzRFGLBr7IaBSo1/AULNiZAD0HFTBJTRC8oi5LDZy5KScR2cbt
8CnSsAVcYftQUPoD9V6q+G82B7qLc3rFoqzi55mAUT1JWYh1DB72eB+ZObeLCxgO
YHSq0nMZlf1tATU3IB3MVJdy/CFyoeS5v4aUw48sPPtJ8EfE8kKqpjofA1nbqzSC
LUjiwAVAhvuX6SPmTUARBHBCQ/BRYz66RvWOW2OGgxeJXI/lqxfNfD8N5KLHUt+G
TrolFnZdi8JWiP9yAaoEYcS0mVwtQ3Y0I+TWbLjGVmG6TjQGhSaeKXHjUVY2hXnN
2gwAVQ0eUVVCZ6AWc+Z+UitObWVFpobhzvEmqnG7MNwVOWSXOxu31E40zMpNbQEu
HjcRrT2cNKPaQdzwLuBdvJ0EGHnCHvuqe+ykow63Yn9FBpBcQobMQgqyN61ZGtDB
DtbzDEL9sAVvYkXiHyn3QBprFG63BeWCiKZyhTBLqDq4g4bNp8Q2GVEy2bB0aWkm
KIyImTfeHh5Sa4Obvu/a6GAQzzuALZywsILSvvqVwS9X8bgWhq252EGNfeiBjjoV
Kuoedgdca3ubp2Z4ZEqKuLHkB8lCzTPx4xJ9qhh8uIphlNqlX7UcrKJQu9p1Ejui
uTNpMv+2bCPRaF0g+3aJdmRMqAnY/rf4TQq7R14Vpmfl80ZPXEUPHOWe1HLiWpR+
oRHNq/zwa8iFt4fJIwhEjKNLCCugbawxuz+Dl9hSvwLlX1c5GOXXyWEN93yAFNn8
MOuCuZig/wqrMpPB3Nosl0rKOlf96Pc3jFhE2fe0THIUfTEUZVwJeOn4U98pYorJ
VLScL/KOJ2DVynRp1HsBhQTi9VveSdhjE0+VzxkVWkyPCYLwmgXpcvk9UyoIrnmO
iI2XtdIa0VIMNPndKwV+dm0UbwErS3bI7AIMbZ4p6WvqVyVfPm3xtv7pk0asOyD4
TfGdNNyqAZQ7m946yM2rJxZoiadb3WJFZLsivVgIxyfuwP1m25tLdGcK1d4Z48qB
1o4oPhqL9l88fgDMxD6ldOx2N2o5/d+Nx+iPyWMSNHzhZdEPI1twqkMO25NZEbzm
dnIq1w0mhyE7XhJJrJ3NVR8BqRS8gl8VWeQrtxSCYCZS6xcvdZJgGLuzoj+lxH/D
gdBQoajngIgj7y0KQe+9dh76yJfyJ7oYd8fFZVVI2YS9snNI3i5347eJKkeOmfIB
dEremgmleIRxD2CNoTLPGsgRqsTHWrhD8qy5IVzrcalywk6N2jp4hIrGgesCXML/
amSdb/F471l2Eq8HQDHD6ELZ62GIv0Nhy0At1YY1BSYmIP+qv3rMhWy1wdNOAcWm
ATgn07dSqE67ohEjjzk6IoZrPzfsnCUjheq1B3WVHHcw5bkbo9zrnt2HJLPILkkX
MiOxHHeRwImHtkU9tDFk2TL0Q0opmDCXaCCxR1Sld74Z9hc11AHf5zwdqrhgBhLX
c4GSILc2WOPFXp4MckG1hxqrUTWOgilQ7Z3l+Yak9RCWAogWkvB5bi+g9bZkNLLc
KhlbfCnnf1xolP+i/euFDdgcWSmU1+wf7QITNuzdEuLLT3B7r//CqKE5aiSOv7B/
SEQzC2Vfw9WAUh1VDrPZpv42/kyW4oAaFISBMfolcs170FPt01XjxPkXWHrHol5n
/QCku47+cGjDJWOPl9gFgUK54nK8XtRX4R1qmmhd3QsKMGDSDty3q9quVkwhsxFe
1x7ENcqplAYOUpHPISj79FhKkXeX0xzAVD55k4iXmi6iRvqmz/utUg5+jZwey0zX
3CwKwQJnbL1oaP6+lnDJLFtcsEggYSjSoDTleQkrrp/G8qWozcyUrl742M4FwgnH
hjZ1pUUSrqE+lUsO4Va5inNtBXMfeQ0olpaRoSwlPnHmhH+UdXvWMMUQUeQR2Fyx
jMaT34vGTpbLwBltJz1SBousFwoEh2o6IDETJdiinpBW5VqtijHJ8Sfu5RCmpMmJ
knpdok0t1e9Bx/0/IVZ2eBBMLAWA70kujHOea0Ot2JkbmiRd0i3is79WS0Mc7SXG
yz5TC/3vsHiaZRI88MniQRFxB4b7q2mO1e0iQ4uuDR3cbgXg5h/OhWmv7zwNCafH
ArXahsyaXN5Vfrxv+iNUmPAzozhJ9+uQoR1+OSD0Egx6VMioesBygZsOHvjBPpqt
24l2gY15uW1RTPRrsa72jhv2XwgwE+IqhKlMK7T/GbRo1BKzothhvHZxDRyDMSJ+
7cvoj8/GPrsfnhI8V1Ep+zx0VFvLQfm5SD+nvaMAnTLxgDLxjZ5LjZB7k966XqwP
QKxl9yBYhKp9eMRLxqt61RIIyep6FUcQtbJCsWAA9qjMjYySCu7El7No4h5k644e
AIPVRUptW/srTl6oKiULYYTy79XMwubNEyaMw72twddCnxh1vT6xHhuqKEPXu3yN
wgW9Bhh1MHa5lpHT8V5ddF7k7oJ/puXyHKbFNIg+lRoyRbinuuvqD0sw2gcwlH4H
PSqlltRgBV6YFQIwxmPccDIhF94wqAjJDowy1IylxsUq26UARkFp+4mE4lyD3tN3
eg7VLLf/+UfHP3j8t7Z3A+IBfOG+mgrAFxvi/y39kXpvNr5J8ZNZLognxRALOYIf
H1QNODdqI/x7oK/pINTXOV+l8N5lpM0vsoOmt9GnVPypyDmVYVXLiRCEm0EaPbcI
/EpoaWBAL7fZUo1sP/5eYsgmQQ1UveDReUI/06lS1Td5WVQ75aJlqtCYJSbRFHOV
L71HB6/zLPgDhOdGj6rfdg7YdElEODMMqyTs5v0sUf4QPhOI6eNsBlTzEGJD5w2d
drU1ehnWq+cXvfcbQzuc24/soAKjUuVMmv2Fd6I6o+GQOllUrqpSZvk0uZZeSBdn
mmYsIsE0PEHIlYKjENAKgJC28+G0X7iYxuvbPY/kfROs+XAXFWiKh+BxMncdbnJK
e50XmhA5lKOmgHZ0yLqrajmRCG9l67Pch727g9Bm0Yn9Z6j5AsJwdyItl3NFrSQS
D3Bws0/wvgA9A7xDiGTtih23/EBbtniDLPxHCvHLTU/0FqH6DKJurDXdM2AX5Zho
z366QiLQMXtJBZbEAmO/bDE6kLvKEtGCUZdUz3CCfzWuNCqCsTfPkJ27bifD76XF
sFNs/RLdGN6Ne5zYHp+eWnLsOgxonJVyEHsfZXRNOVFJS7l6pZM7dBG6zeMFdAg3
LyjRQEGlR6mz/h2Oo4rnFfV4O3qzbC5k57K0aNmu9353Z8a5jvX+dLMYh/CJHyAR
XNTTZFc5GB5zob/WVc9vv/tDIOvNIbO+IciTfKaQYbRQIAwgjPF63Wus2pjFOdie
sEVkBvXVaTX7ZL4VtuW+Qsqy7bPJ7oY/+ngvkMqgJ+8OlLm2Ez6uH2d547X9A4eL
vPHrfOqcJlyKDWZbMk1mYAR21ep7NhxtpgHG3+oqB2oC08bx7F/95gJNRVqzOQ4m
2+NWOpKATLTjU9bZXn8NMM42oKp2LhueuefAFrb+YkfHIbwl4CCxR+TkwQKk29Cr
stFXW0jHVic0h9t0TfXvDIuBWZ1dqv91SaWlunbrqIBY1UDoRxxMQoIEl+ED6f8h
7TNVcyKvLpKZNw631ON5nQS0/+90RymG3lfjpzeCXdEmgr+ztAl7YmuSgYV0cJGB
Nb4lEpgbJtyrGaLH91cp7r/2lt/CRj+ggn9gqX0RgLBSl/+a4DLVbTvW84KWzeEU
CtYJ7b1PFnIxtT+oiqH9YZLRi3gnomXDzoz6PaQgvuaGRORF1kUdEBrh1qvTe7H7
EJ8zUeu4ehIYwXRFG+E+SPGsnPGAv9VanLQ6LRtdQYVgE6WhqIMdT97J6t+IViaZ
YwpGvIdTOSClfshbsuIIg2m865gQ5UbumsCO8agIzMC7qF3EjgBzZQRhbOeVBQqB
uYDgjE0RM4w+iDlfVLRHGY5tlnbDqBReWDPUN1DhBhE3RHDBfxUDkx01XgPiUpFH
lXXLctv6v35NTORjrK9PujQsu0CP+5XjLmDHgzXAzDBikt0yM2kgDqzlo8ykSiSG
IykJggNhT0gvt9OPT31dJvV0PvYJc3HoPYxa7HWw/fE7E85lIFYJG7PZYH7ZVP0o
XCn1N0nEosNxX3gKK0GazxVNYhsqvgiINO75EChWSJx6VXPIKUm3fb1UP4i5aUTe
k1bLMsMYA7rwm4k9U91EY/botw72rfdSaiLW+gw8IGdZT9SZKUtQv70++midZcx7
25o566ri+nxO/qk1Kx8TsYQ6xDQQrhjyvxSzVtPGLfgF2hdWg1YCS2vVwN+dTkyT
Sp2jPkq8rJzpRP3GmRdpVKHzrTYVQth/30S6KJbK901LzqdAhI09qzSUoQ9NChut
47HIwYUbSmTwo3/Kz8pyVIJK96OATq8HpNjtC4boIvToZwjVM3izWZvPNr8/FpKI
gQtfiVY629U4AEDHSjvsr231ShYnHDTLPw50QIqRU33zxt5UuZ84xKqROjfxuN6g
+kZ7uEQwOby1jGQrI+Dr4abM18yGTrKn00WE+dmw6NSYb3ffyAGjpoOXYHexOg2Q
+GvokxQlIA5P29J9tRQL7Je6A6NXbybrRApUuI4dCzs3ZiSEZozj8GyV+kB2hKJ0
UdIjjcwY0ZSqHzji0OHEwfRahQwzfl16YbjO/V36tor3QbgQNHc/fqPi4UWUT3/k
dML891Lwz0qTHuxRj5xjOYN3SJQ7zPWZgNpsC6Cca/t62/Sy/56Es69FxvrQHhZ5
/6o0JpJ0srAnDKkzCfOeY8pwHURbvyM7I0XFwJAvryqBOWcjn4XQMfDNjJW7c1AM
PhqZF5fWR/n5kA8ZLcqhNc1/YKXrfgbGY1HNTuxLEB1L3eqA0iXySmKbpjDjywKc
N9BG+S+KSHbxDoDl/bJD0NKblyTMcxwG1nXOR03gxhCc/Yk++YXqCswQ85fIkwHq
m5Qd6wB5LeaGckR5ed1Te8bB6ebhXYJxcbzNGtEcSKGTNH3y1A7e7yUq9tW8Rssp
dpZRfWCGOwmjLZdtfBYy8/KLGYj5UVoC7Rau3niXZZeP5lQnRMQ/HxjJpIwBVRzk
WPn3Iu5hvdjTRPogWUXON2OcNGlDCvmpqizrn3PhrkO0V+hrtRg2/2SYe3655ASB
mdsyzamZXs6W2h+J2lS2SYoK/HfkwMJFg4GYH5Id/ChKh0lrcZzeIaRnfsivPAa8
ZeJoYe82TWUl5wGioJEF9GPmHB9X8q66mYfYyTAvqdms6qqHJHIz42RSSiVJ1lFJ
Ey/5n/zW50LdIlFvIWcq9wIiHVwwJaITCPNKoAZTF9KqhtwpEGnBWq86UnbGIkrw
5WdK2LARkYFk6CipHj8tIKFDYIap3gGzDq0A+mntghFwg8ihXLhCD9KjPdNX+VHE
GB+v4GM0ojtRRJxFEN3lY5qx4/N6iyyN6l84/QHoJQkjqB+2KTtFnJmTwu8Oq/jQ
Kq6egxDZMqMAhwkIh9loddv7s1dcBeKrIrq1HvRBBHH4s7Ky97aarhrE/ymPnTGb
VJqKJhGq0hz+R6E7hVpNPkQGsoNpXsr5awxmwuu2Ghr/w22qISVmxJyYuwdIUkzv
nvZ2X/hRomA74T0mDjipAt2Lun1Ci50yNKfSC09Z5h0fJNMrJmcOUY8/jv3a3Uk5
mpqMg1mKoNbNBVSAnT0cK3NNaddxvtRTncE1/VoTNsRskSvFf7rBUtX8w0g6NhO6
G8Nhdhg5NViBc2uqZVAvbdx6oS48pYUxHcl3dBQR6WzX7VuLxmNHxd+vfwsIMqT+
0oUWaXIQ41S/gQ8V1lgtyEmT0SgsXx15KWpoCRjUYfxisBVluFtfcnqGAjiEyT29
Qd2Vleu3ldkmVuWNqul383pptQUnJvl01N+AwEGattaZR3bCMoA3pdRCSrrkV0sg
BkryJ9Ia8daeo1u14RhGVAaw7Nvo/DlCHCRKXZirOFodl0/2kczvzTzJSciDOA3b
zy78rRHWcMnfTC+WIM8FfX94b7BIvmSsA7Je2DjOlQWPm9HTonD3drkoA2vNUFYt
b4TwX7Z7mg9QQYDXBIyXxoc9f5jBroZt76AJdUukXJMGnIirVyyOEG5ms2vfukTs
m1rEWowshpMB7u5Gjft+5S/1009lwvJoswlmIJpc8bDfIOuEMxRHnx41xk1dfFtI
gBa3GCjSD+IxcyChLIWIQGpwoPc6KODYP2byno8rimK3ui1HMNfOZcjqZDk4Fw67
gDIKlzjiQn5vVQvX2nfEq8h26akxXVncJimO/t13VkVbYFH+rlI1f9mydcde18zY
RGTaEoqwlbFJ2EcoUG/7zRMUoWYk9am7xipShGDPhVGtI+zb8Sszn9WjlCFGJiDq
u3EXt7QnlZ3p7uBv9KEtNbn3Tf2cRZxM9nzNp9gNwmQo3/Ow21kFfhLJPROBuNXd
kEHon4YZQ3+UUnlS+EawmDgqTa+5/eHzXCScsNpTYudm2eb1oVPvn/vMUAMz3oLr
kd15H7voOhe4E8UtE6zfB0AYdxfIKZc6kg2JUQ6AiWxdnEU0GqhP7Dep09D24JZb
ssYGfPhWx1uq+KEQW2rYLbRLWs3d/hXh5GylYwh2FTUOATdfu0p3wkBWElq5DuJH
iXi1lJ1EmnKCGQr2/NR7rvpE1ajlT+H3i/NGy1WOGVjyAjZ34oU2kdz9o06n3VZZ
VhCiY4Pjn1afVixth32vlVA+T+3uSkyZZzpYUz7G5/FoifrfEbQtnPfPquUcfWw9
DfQqdD1GasR+QYFgpBPiRitZZSvePZbWwHePkN7YQ5iM/+V/ZPS6pi/1ceiMTMWl
5EULHriZyTxkjbVJJu13NiKgDR7/4ypyYEtGTRWMlvmpGBrek7A9c+zGirZB4ySP
CWl4GBxDXAiMVzy5E3pIBbSm6UJ0AScOfTb/mU301ighPl5c/uRG8PTtgeK3j1pI
bexCBC+TM97+pcIds5ze23I+eLam71WeGRiqO9a+EcPEzU0edAtJJDchswi+Io96
oibdoCGbiJQMzvVIV5ojDHJxnI9VlEyPGPdQ4yx2f1QiU7LP1KZmqnPQh/nxNJOv
pEZpfc5AagwqzdadctOZfB88Bh/TA3c0wN3iMS1mu4iQ4V/bjGuNG3FzuTzUldwX
5aW4W8NvXFaARdbUhsR1xyzpZaCN3sINw2XghhKom2BRee6Nm/F/XcPKcOFjkRsn
9Rl7k7pSaqGHJWiDwxdpPt4X0gBfrzJjbr/+K7vDeNjmt+huDkx2ckHYkYNti8vH
WCxYlWWDrnG2qGMbz4ojsSkZz7TbbphuZNmTwoduGSdKsDpwlcbCujsBecKBPXc1
dZXtGm7qfSb43tIl2LtCkx7BwhNBEoWTS8q0r1dYRWaohNfSg1DFAF/hxpp4TWdG
hgC5muvOpdCz+jkJkUX8MqJbsFtAdOZqqVBnhZvy7709pPdknPrt3VyZ9tjVHbnG
q98BRD5CkUdhsy61+sEOBtsCGhwVPtUB0I/PdETEhYXI6Ls6Tc/RCTUodFrNjMYe
GX4wvKcYEpyfRVOtdsdIAM7SEuTg9YeRL6MblTFnjOV9jANUu+9ldSkYsR8gZLOv
zY4wzehGEvZq+jFkWdl3E0Uxs5vjcaaJiZtff07KOi+oxDFzAW6OgWmk7gsCU8V2
zeVOmW3qZrGDUIPKtYNcrVTkeBmCHVInSGPrhNRAZcSZCHvgYCulGfpjuQj6K66+
hxxbism6/XSQEETSdeCxz5b9z+IgnfvxDpdyaj2NSm+w88UKmsym1zKwteugYs5g
A7TraBCCaouv9CPNgwBUXfEnbwpgNmmugNe//LQzZeAdroQFQzqZwEJIll6LlgEZ
JX2cK06t1Tamb9449SXXHwO9sQCKJMsB3uuDAE4rkfshhj0kBs0XEWYI/FovHBMK
Q4hWAqyiLfPbXGQNto/dJ07qVjxCmBTlNfsolVuwrh9OyS0AW9/hVsxv2jh3sW66
m2q0xoqR6A9n4Wu6yXXhnYgaCexwJZs81I6kgBx9cryjP+WvH0VCNt5IBzPPwdfI
ZKV7sgjkwvDR9u2asNCs+t7Tcx37zpeJ1i5BBkg/+rbXy8an5Fg70WBTfErAMZ0v
TLIDn13aUaodPr72P2bXUhPAu4R5xl5eIHcinEOm5PdqdJH4AaMwRarqH9pXBrDH
eqHDQZaB3BVRMkIkeUF4c122LZD9/gkSZQQUgQgTUCTZG2fcWOjsV+zVFtCJBJK5
NP6U585zEjFDEDq9eIPshzhtjwzVKutv0CFOLZMhX7KRFEAImMmyZNk9b05vjPcH
FEc2zHQiT2OUPBaviGSRzR6Q2k3AN4O7BEsyA54JeJoQ9d0Z5tN218YYKS2tstOO
XxxJBFcWh6YUwSWOoPNv3EREVzllFoq9MM55nEI14RB6UR+7owSVcy7oVRXdhpA0
YcvguRTnaT108hJaSz5Pd1irfGAyKbV6jy4MinrIUny0CaLrFzD3NGl+70AEk8KH
RYjbLKWfDmP/dGMGIPQ57G8LRevVHAcqxT/KtLGZrbhG7oXsyx0cKFCP62iDksZD
/vgVlz6qtib61y/azUqXw/Vn4PXJR92aR/TCwnwSxZPh19+FbW470aNyRLS6KOQe
bFXbGL2LJaY7cDT+ukRivPsJfRxlBhNlZRsoXgdQfCkHJwid6WEdaAzZTYc92zY/
pSktiP9g53EH2DNdZM2U8w1FX8naS1vRcgo1ZDMi8eHwyPowUnipf127JRPiLJVw
KuPZ5iFYk+t4niisHGtzz1WkRr7qAFSmG7QJZ/o7DjEKrwn0ts3Tkk5MpbzbUBD1
gZ5+kVCbvciknFYR9Olx92iFQNGjCUKH4jciazgxkaG7/HBjFHYsCuybtdtKMGW7
Y7PK65mG/o4mHJLOPEfgrEeipHOXal0lFZkXi2YzwyZC3lSsjEH8kvzIkLYBuGxP
ikC0QCL4jZWVvOzUikJmqCaWgz/txFRRQDa1zGP/W+gFcD+Gq7eI974qZVK9U0uI
bQwPoIHHuXkAP7ZemkkcYEUwUI7y7LcQ42y8Xg16EwZvWllXABs2J/lbxglQMTQ+
Bvoi7YxaePm9Xkrye6zQQEvr7DWtM9zzPoJ9Ur9MmznD4PkDw3LfW7z1RKY3N37t
hdHdCF+pJ2wBwN9TZ9il6XsfzuwhB8xGMONR0gArkj1xS2VGTTKe00k+oZ66pd43
uvh9bSr2ZxRU2+jKX4NsPSt06/5qZCUi68VXJLyobtTW0m8BkGC4RauUagqAhXFU
RSK50OJRbCga0o2si5WExeu3DNLmKJzYBWww0fdkCNsNrIHwWYVnl7K6Y8YzFz57
Daq3kif6ya2jxSCFqkvZ77mx34JYuBmCMPjJk9fzkhj4YPc+rcHzS7a4O/mbLIdF
DajUgOIHD1HE6cDaEfoPn++2wjuEOiilSQ5mliRS1SMnGoG53p/UxY/ZUSEacm37
U5gP1xWNOB1mWHwWKvgQmYJDQdF0qB1sYNXY/NZHE5fyjPXPzOdfNvVYfHfGpSCW
yuS+wTcyplMFnZgurvAuL/DMNcNl4Q/cd0twcizgo1TrUUyZlLtm9OREmITTGKCG
BGwmXKM1FNtHj6/ABzeZ+loGMpLp6OGhtcMiYrDzUf3AAsAviwTrQ/nQHKpH+ZCz
UdihwHA4iEe+UIitiTDypDVyNyvwisXLmiHUT3ur9L17e9uVQ0nTQKqxfBUN7qpR
tUbFmA4Jx89y1TDbLdbe3XvJtT5VX6m/XdPfgCk6VBpnf/U5rI0CBFZeARZyaIny
bMgJbniCc1nVMrbw5wDw45OW5dcqghvq4yeizQeZxBMJKNpUJhOb1DuCsEnZy1Pb
Tpn2G0iZOQrcofFWuJQ20wBhtsZ72lSGTnnXgPFtWJTPvqkKepflo8f5zTlZAIjC
DQCTp0ieGtq9jmFzyfU9+azjSjAqfk9PPpZu92XGFDzJCWehrPKXTI6dAgc94lvI
ATUMObtMZ5F0b1zmLy5b08CsUDMN9jL37TEBSdv+ads2ZsgnUz1y3k/9KNrIpB4O
/Atn+3PBG04gnJ0vcmEdN4targm4e5nYIw5d0lw0YcQRSwg8Ve22FBQO87fwB6b0
r83vTruTPmxwga5+hzv3k0A45eKdV/9EfPbxtNCjJRQMWWWQqeGAdse4mdoY7gYe
IgQsGXebhR/L55NW8H1SDPAPsmf98SwQWRhXODptDcgthHRv9T9G8kCdmZzhNV1y
Mm7jdxvfbI+l7laCzQY4z5d8+j9RWyDem3/qC6PEJgO/yMhgF9XmPs83C3ZGZRPS
1RA8DVZPDM7+Wcyf7JZuCvMJL3sKM8puBXq+T6YnH/ikBMQa7qoC43JDeNtARXSm
SXjVorx5qz+d+AcceYwepS5aPL7gp9zwwLPfuLyE2bIg7w8cC/OYhaeoo6sUu6VB
jzEfScBo79GiAVOGtsl75Q+sJRR3+CCPz4pQR6pa/LzaNzvtkMUc8wAXdGaR+1HG
I8Dg77/JCvoUys8LmR7TzIgAJE8N9l0pqTgmYZGZTW7lyBhwiuVNyaVC2QL8+0o7
ym5u9pFU0SRcvBeBMvSyw+0uUYtqDBZKHRjhgh1JkRuyG5LrF1FUNdnlNy45fJFO
BHi9A3nXWiWo2w1mUb0g0bEfHtZxnl58BZQ6duj7VRMPWbJ8nHbDMa4xD44N1LGY
1e16TFFPmPL8zjb5dAxNzrlIzB4DulnP/wdkPO8K3rE7Q4d7qJ8S8MgxMVgfYmAr
98NfqxWfUJ7NZSKlRNFLWlk5suvvxa2RB7N/gyfCjq0dS26q7jImRy7NcqA/Z9dE
iCH6tPUGxWdIABN8eIeHvZhugo4WBZTIFxlb2ACCjDvRS0xds23vFuFmn+dCCl3Q
jkX/RgWlQvBYycUQxdtw6+B0IwIoGRmgqocz8Rntp6AdJgb3PdRshrgbui9luDnj
dDJpqqZlqxOrmj9z1xLiOesntHLDrWz/6+jAhaBCxg96UCGybGPWx8tjDTpDHMJc
uBnNaYAPK9Qm2sx8P6EqFuz1OvYKiHC5NJDi421v668rjyNCZwDg1QWszQqLbTbB
A/ZviV/ID2VaAvq8/hiA9rBFHo2jswhnXTYNNAGYXTbyqR4B1eYXltN8vnorCcMm
gM1AdsanI8hcTSDMnSwZsU9EqMM+Qox0RzJQASYOCrY/xBvZXHloiuQYW2+Qzx2Z
H6d3bzcbQPXrMgCCwWJgHxkcApTlA7jbHXaZkJtl/DfSsh6v6uBoeHW2/QNZl91h
c1VCUDBg1tPouzzOE3PK3UI9FuvB3DaizbBQKouy8IReO21olZwctGmvKmqcAKSD
HX41XtTyTx3JEh5xuIuLE5HS6QWakcfpgSZbbRTurmHTVy152NpYsHMaDrTU8VtD
x1kJTgeztlZpC4eDYPIbcPfff0OimkYq47YtIglvL+5TFQBzUNkEHpvl3wAqNwuf
taR/8CXbDtgP5GKIkbNh7gGPcpSQiPOk4w8Q0VNkEIBr6XdCCuedfHuF61NrjLHg
nb0ceZjMGphTxro0zYvzYiMBD7QabfDI6cG0aJAk8Cb2LRCfizjZE5mbE3ilHdoR
/NW70Pk2Edgx4kiqeTaptgD91kWj23lJqBO4TFZVE1Ot8s1WyGAzezWYxrTYwKMR
UOQRxiWxng8J4JK5qhAyCjWzbq4pYJRX1R808TFiRlOQiiIcxVVNnhQYhoq2g6Uu
H18psGoK1EXyFy5RVtMyWBkXELzhAckE6YYqD/cOmW+ILkFlO8gR1ViIGgnn4qXS
3zq571pjONwec8TfLIQ/wvlazm59HgVdq4LtqTUql+9mLT9axf9p1N2rIDegK/ki
gTCJ90gmMR6D4syni+AvV8WRJVRhZ7qEq29dEaaSSkyGo2R3iaG6aZEEPZpRm3N7
XDgOlSjlx0vD8tUu2kKUWtpBfvavXHMLoQenae2yoJv4dUc2b7JA5Wt6Kx5iL9PB
MFjagqXVts21cMitf8KDsrlgJfTq9Dno79DAKACfanxDBoIDPM+haaFUpd0W5RkS
7izxMDqABzuhe+skLbQEKiMFtVvwQ0asK/rDM2tMVga+62NBNVku806+VRfYsufc
QT0YSQixTBk0QedQqYj5puhRgp9PwZXBCYpAZPjVOQA7HHALKjUVJRGci2uHz/yM
KcUUGb2jewmpH0jGzS5TZILmKvmLUgvvAgyah06tLnQ+GFyFDwqslIzFPBSnVuDW
LSKT9j6G1gGGF5YxbtMFBfe3QaDacadHgZP6G12Yo1X9bZOwdl4dNlVj774eDibo
Mv6RMH9LvxcNexYiGrm6PBQWbR+k9WbCPiTyjNOpIpCVYidCurdwfs9a9TbfpTI8
EGwlJhEB9pvwXNlYS2bSFEmNPlSZx/kdUc60vYR3i4DXz3VNijFQrz3avfO8xhdh
LI3Hc3KOXRrWRGpExLzZoIDkBEdrpkaN79n9UsFPfs2YVUAdS+Q3awHlsxkuNmSR
30tCBx74VqXHpca/iSUKNmG7/EPTWXlxVndAlS6NbTdi2i9bruX3yftV5NCg/qBi
MDV+yH/dSGnIjPbE9vsK7UawHSLoZrLSCBs4mIC1AQWqR6S0+/Kkn7VOdp7ZSyYk
FUF5d8rrbixyEhR6+hKNVk6Q85wNxFo+6kYCOEnZjzAlsWoi2UIzkuGVrgflq+J9
+g6dJNMovPeH37w4gcWw+IYuTxdG3UdCpcpS881ksAbwQimMoCEwWeXkwF3/GXA2
k8uBeJhYnet1nPZBJA2zCVasdiyG16YDgAkVbhZTLR66jwnbOF/oI4VwyZn9aNAf
BYbscH/4PI3h9ybQWpOks4GqEUqbIoNZD3r8FTEcvLEa8Xnimv9OS4y6V22g7pYU
Z57dgIJaQlJQFC1hgum+ZuYveaz1uXYtNOCbZJhK8LkYr1H7n0qLY//9WIk/WPk7
1HhR1l+F5Dsh5rl9hVD2EP8zzef9O6UIaHurP1ST5COMlEOlsi0mxZNOR8RzbH3r
25v2BOAOnWw01W1r297QuLVq6VBIAn9aE/Q7eHi0HYxLS8Im9B0J6M9UDlDl/v3v
pw0EkcUgmC4rjNYysZXfoBw7+JWS1s6IHmC65N2r4CU7jZzhGWaN48VsfKeztUyV
W02Fr1dPqSTuufG7N2M/Mqu0DGLohfXFze4vZLqXbBRZuSb6vFjKSVUz4Y7x+P4Z
MF4znYaoZP92gPSN/8uJvomTIYt6ImlfLXKvPKuZcrhBd1DuE62UiEA2evwSTdwJ
tFJWgIzWcDXK98bBQeS+VW2HqZt8ha3pUglKTPoq5LmwnhA+c8k9gh/aVcvVDJmQ
GgNASCwTaIvF+68uhsdKg5qW4vLEtgdORz155fVFvkyOZadUiJ/HXT+gcDBqYR6m
sdofnBcq3gFbJfGpmkxzMyHyc3AsUSef4x6vJ4ZBsmaONUCFIGf7YhJ0dehLMAkV
vNI8tS4E/mVV973FS4qrQbNSHJjuM/enslc7f2k978/2cyRcwk/A8104BC3VmrWh
1EZGuhh1VZdkwKdTGYYrnvMdbnSAC2MFU+m1WUQsDapPqT+OgZsTVr+H9E9XbHMf
BkLgHVlCy3Mc2/RsH1MTChzQvTD2d5M9Q8pym+hZ7+hKGQsXjJz1s6mZUocpP+v9
ns73RsATELsG71OJlcJ6aHO9ZwV/rmZXjKYbraKwx1XqfDAp3HIhH+xsxxTw7yIx
v4QBtRhPVe4hCjBCVU26fDlpxuSz2cmzqoJ4Wi8HFtrey3PJ9o6omrO8BedlAtza
ljuytRtCEA/0A9ofwv9vj4aRQFQWgonmVO8eyxHUFv+jBi8DUO0fIwRWysXu9o3L
TspXlJHUKUfEimBlAoyOIgn1flgXlIuAU/aUpbAa0pyQsP7BcLTs50ZElGJ2vreg
4fOfGtmYSUVSg6epumYAfLIZUySw5eIOUulZuklUSalYHnMdL36bh/u7a2qvzJwp
dAOfuCpOZxjJLYBHwnR1a2ga1fR+gNLPk2mzYYRYtIoz1JajtrV3oEbb/BKGAzvC
RyqWsPjPxrMXM3tY6oZDnAKPdUwFSVL13nRonZdn2Nu/Oq9ol3r+SXxW8Ung/bWC
rP4A0gg0U1KsSMwg5hJDPsC7Hagve0qKiUd2mySFyUcRii04IDn+wARItUvgh+qo
/RaugNB3SwJRfhrpGXHv30GNXcsbwO7Jf5HM7e8fb3QkhCdIc/YiopDkqmfNuwOb
Bb7x/OBMUgfEBjiul54bEesXd26t8ru6O2r3lO4RuXROYtwdyb1NYKs9vm2gbJt6
u59QGJXYfTU3Zakz7HCbVMitWoy8gsqrvS6HhLgXhbNQ82Ig51MYa8g+3vPnczSU
CE+ImY5hyUVGs/i/DbeOZ+ap9H/iF/pSDVZRkRb+OuUPVaoKVni0X7DvhvFUboZc
u1MeypBfzUie4vLaHlG7Dn7KZP2FLnY+genhjGbjxzrb0WRAqwJwJUY6EHANSLR2
MX2BB+GF5T+9kT2RknB9z7iqPlDkHK4VumyTXFxwT2jShE4DEXhW1sT7JBjS7stN
MeXfLs3/s/d7qS1f1NQJ0ZrtzjKhpcVn3tPfGgNGo2SZHsQiDjLsVgwPP1M33YBs
IxXcfvVjTE2LmpELCe3OqNIb9cAtmyLeNJGnzrjWyWijBvPOJ6LuI1ueNOT9lIlK
7k4CCLvdTritodPhCftGKrfQxE4CsfHjOmRaKQmWM17h8hr6Jy+j8zLgIdlDO+mh
OfoNhhED02E0/+Y+8PGRg4wWdmxX6Mme5dyBOqVUiCBdcWetEorNpHe/DpkzVMl0
YtWGr7kLWOSlY/Hq4WIuMvpV8Haz3Jvrgeaj+lVlXo/gAgC0xZScQ+H4YH+z6Fa7
ckZ9haxW/WR6k2Awm/Dq1/T6m0n06oEj7WbK/9m4NkUC5JwLlo00bNDEg/h9QcNx
cIeqjJpVYxYTabTOoumzMHTQxwV40kSNKGP/9CkRzLO8NWFXAgBBFt/KmpEHSdGZ
CqMmXZeSWOBfr1QOCgYr/XgOM5Sv2NKloF61pJ1TYNvDvPBD4agUZ9KVO7BynOmF
Qq7iSalp+w4G+g+1wcOXuda9gYwMHPFovgH+T0FcsNFeM9wc4kiHd1nLpe+a9pk0
4/V619daHBf37goSNQYa8JSleFK4LG+Ua6j1dc3mR9pRV63nq9/FD5tiZus6ycKD
xpA8EmC7nWhnIJqADKE5aNYFd/ISHbKw3SVERbbhtEWxqMbKfWMd6FZvgxe1HrQ0
47FZyoqvRW8c5e84ROCafByrW3+lh8OxQmPZL7LOCxPVtqtdfGPolG7PhGhGnfPL
3RTzEDjDuMNENOVYiHtMDVLnPnl0HPrPy8BGL6UkBhUfyBdI1OS6vfV2YjL3VF9w
O0jr0AudODF07orMR/E0LJ3FuyzbrH7Hq3dhbX4SY25l9J/zspx8BBf2rYpEReBi
/GpEKiHr2qPSMeHwobLV+cv+n/g8kZQRHKC4E8l2LB2KZFDp4UYq4iD7HOOiS5ja
SvZCbhnRykoKjkoEU7U85/eGmFp7vFY8TQ5GwLBtXMjwTyoTfLEZbdAFvzYS0Tot
Y1x8xV2J2FdR6NimPEIt0jZQtJp3Aal1RoZl8d6AIbZuWnHJQ7bkj8ixCX4b0qq3
2uM+NgqB0QXR3xKvaba4TL8WweT9DHg4vhhWqb8jm37Z0ekNNN5diCyqc46W03My
X3vndTByD+IUX7XrtU1dwTCIzCeO8wzsUiimKorLh+66Fbr/Hgt8uIKQwvKpbVj4
ETIgykMs6LSD4v6auRNew9DOMusqjY+e3wrLWCtIlLy9B4LyCHovJh0vd4tkDL2V
3a+EAXtLBX0PZikGjNs5iVTUAx/NjbpCyxc+54/3n6b5v/o32PNjlpVoRltJSSts
rMQ0TQ4WYe1on7TZEbZOFE50AZ1nN671tFI42sKtlWbZJaDFZNa09UYArNdw9J6t
00CWu2mjeLtQcTGSG88YluZSSnmvEHPsbz6rn3U6otxvJeudOot40VV3V5eSnLil
p7r/Jy2glQFRlSWIkmGVIBuXtFrZQSm4P/z2hBEKlru3l1eR8hGFBcehSSHf7qPb
WDGmzoFFpM8CxGYLdcJURIGI43bRi+ehvbhcTthXzRoVUTUT62nvyDPcXkNhx+nO
BD3SVCu7Z1HWyKJrMMFp+wAbD25H02EQMRrdXJJK4xXhwTx6AlVBsTFCqZerWuny
/P8g80SVWVkn7iBTpaka81MxFh3EP2AqVaN20toKuCd7I0ASgItkSBfDy4S7wyxr
FZvKNj/FVy360qaqixtaUw00IMDVsXX5b01jbgRqOgfLe6V/ss2o30NXEyv5rEuG
4jb7P5lsEEFahQUe06o5whfBEIkTyeyro0mBTYuEhKakzMx7lLd+ZiumfScwnm5B
qjnEXkQPPMJFn3lEZbcRAI7PGMQiobjJveqenMn+ERU0M0X1k65RSWzCoFlv0CTi
Cj0JehV4jO9peHpgCZydrOYYgEPM5eYuJxdmaRVg6nZTtpttytVTOlGRSNsvVqSK
GIQp8ceARTL7i600q4UxGSoU7j5CNPBf+TmwDCnvMzMepnh8ymau6tN9vl1EYFVl
r7f4MNZpKOqQM0EbIPVvtJqkp5OF6BeSrmt6M08lnYAxspOy8DJ7RevhjaLD4cMf
Ff89jpZZ0bNNRL8pS6BdYgLrqG4UYb3MEcwuMhQ0rtekeK7V8KUnhSh9mBsTFRoL
r4XiDhswOP68aT7wxClvPOV0Kosu+pFP51ZYKYjR8nqPxdrSYlFZtAfr0mxH7zIW
GeI0cbaAQdwlduY0HSZzIHZoUX65+PePVjvQeRUH/neOWt5e3BpJA7MXTZg41iIz
GiiMDKwGJlZ4bZZ7otwXr2l+NVWH7urjMCHlUWuPwfWe5oirIZnIGUVkL0Y/B7pP
5W7LtEnN4iuw3XvyfzTHO1sena46cMLDo06JRRrhal06f/DcxGNZ6EMtcN47ckQt
g4/2NNcyHw0kmmSlRJBje6ZXaPsGEqps1yrDlV/kJJKc/b39FzviNf1QtS41vRk3
WcQlVI571yfjcfWMt0O3PddZN1Q6TdukvG8s5BOcAdQP3iIKSFGTKhE9F2Tv73r8
sXnMQOQI5fbLpDLZ3bGPWoz4kKYDKxIKRPHUThEK+EzKG0agIzADrqbYJdTVLDTv
mH1PRdox7xT2KmLdqdlHbvx5eejtC1ovnYGBC24w6v+q2nrEyhZtrwInU1LBE2lt
j/EG1N2d17i7hVgfa+znO/UJTOqcZj4zpXNoYwC527bemNUOUMrG6JD9L3UwBTsp
yi4Kcg0vta5rGPZgb7u76Tn8ukb43lz+qQ6+2vlKmQvY7dPHLygu8sHO9ERNMY6s
JTVv/9oqY77++MB1VGiKuBygHowl5T0rLfAUyL2bQHgnBE/F2HEa+qHCQNFqxJ+t
dgNaLAWpgfw9rtGlRF1VEX8ZUOqhjfEgVVEl76nu7gIGHqr0EyISlAdheB+KdGxV
86wjLMMZa6OGArQW1smjjxW6dzzL2BliafJtgGDxzxDLvQXdoY5xeAbxsVxYgKeI
FS6+EngVfHLGoQU9P3JCTdlCywfHAu7Ypj2QqfjB2XLi+P3lL8hSp3SIozUQhIbo
QGU0zJVrOcsLBHIUPqeCnk+fcfMnFyHn4gtmRb/Qvt6NuLktEm/DxySzVhMrJFLx
bE5NsRWvyPK0RJrhlTtTrLAOlmWbWrMe6cIc3M83PPCoeie4HlyB/eI3QIIeKk3u
6aiV4sQ1llBd8SljqQEfn/0UxAjC5Uevdf+Xel+7mCAxoXTR+KL+qL9iBG8HUItg
MqQGEbAykx5+YOEAYMw/OYT+5bv9PITGI65JfhzudZj5R/jEiqajDsUhsJDabVRa
wtovz7+DmjfPGpX3DSq3OSBUNczqDwI92KNxCS6nihxyn6f26eePrxU3AYdeM9vO
DyWUXSelJx990dZcgX20nnyZrMjYynzW/o2ERJ+MvseJdE6TlDtJBgkU2ghpg9FD
pO8t4iHELZ3FmVhUJs9wmspMvLPRmwLkeAXnx6T8ZIKrP2c/+RWfJ25f8nSbsu+T
lAgua1l1AEOf/K+5DsNKmthR3JXzh5lC5vFsKJkNX4jVmGdD3F78vN4oBNKwzfzk
3GDDybXVR9RvhaQHBQ3/070UGSjh5jVfK3JFxk12vvTdvWVX/xUM/cXw8u3THDqy
BFhCHq4o3jVFLmAuBulGjajRVlbp1zwh0bO/ECMbEDqS2clP4SagVgGKZzC/anB5
av8x0uixSR9x00jyj2Zn5trvQGcQr/R8oOfLvF16u5nwySuQIcGuIw68Qi37PviE
nEtvqo41LrhzwqpReXkFS8F472z26KXS02HvY7MhHvmvygVi42+/o/2OqmKRNBUl
xL9ydPZtpV2B4YOStg0bFqPVmvMjDD+vfYV+9kaaTVpFLdX0BaxOK0uXCZvv2Nkg
Hlavod0GJaEbRZ9VWq7z4L3E8ZksFMY74kZJlsNZ8+d3Mh/idQs+UiQIizP/yHDQ
wb5UOieE1UPOwbm0isdaRFpUun6D7yp1HJMssEVG0e+LExueuCkkVDBQe8FH5PXd
zON6XJURHeIfzRZ6Qc+jzpJKZLZn4L6xGP6r2U5LjmQgysIrA1IrFcM4pcfYkP5j
f8i4T9m58x+B/c7fCGdx67R9goiwU/wlzJiOSTjl7NlimnL8GHNJZpoAXigtjG8/
aPESo08mxPc4sIJ5ITA3EdwMRHfmG/2kWkPbZoRXvmXV9xiAJlXnsffA6irGYgOY
n/LZuaZYibtfjuhGoHRUUeGl3XOBl5r7vgtg9bUHYniXJBzPA/pS991JjheQqsbQ
y7WgM5ygOG8zffsmhM57kCNtCntUq9IHEuhGr7hAeMHrSRVEkTjPVqp1Yaqz70EQ
N3V2d3S9IvNX8hUeFDyVIexvnrvK5988A4BcJWqqTHtPD/fNNFq0tTj1M3otBKtm
iY4e84qmHSK09cn9xams09pqPAVz5ZIZ2gi8Xt1bJsyeF38kTylFq8rHJ45eEEAh
vMmmhyCQOrHOxi7kaG8U5yqW+3BS63Km4f34UzOvyUx4n7CcBi2+zSSvk4ixig47
ucgg7dWiQkpwpwAiyIFSugAOmsxvgP9Qh0QmybiUt+2XN3EOxjcdph7SPyIaFKlH
Q48QU7VWUFs0h9yVZMVXMui7eVinAIUrV7Jj5QlEv0DOK6P3TtmTUbFSHe4jS7Wm
+eJm7gkcCIvMMv8ZM2BXQXUtu0pdxhE/kU6KgkhwO7XwhRhQEKPxKRZuFH18dmuU
Hlw8246CwGMHepwNKiTubz36E9A/wSAwR8Erph8IwcvEb0zWVa5AS0KgPU7aiXjA
pr12sG2r3MSEGfBYYyFS6UF/r1YvVaoTVauf9H8FdpXUWPImANnHl1E+mxBFpe7H
+vSxC403CM9S7xe004Qps8muCaPtVfagbkL8QP7oBDoJo+ammnHgvx8/4Vjb8fEV
3Tyc57Azz/M+MRAflGCX3Y1W2IUPKkl7zFyvOIdxeieiOnSZyoNoqQDm0gJRebSI
Ia9ezkPK1BQszcA4A3PmNdTpq7s3Yex6M6llee8e1Szt41QvYrz570bfZB9aHMzU
tb12WZdK2FbH5KhB+3+m5Zccz7LNgJOMe/7QaMvggBqot5LyPGTgwmumCJ2RjLRB
qHokXJZmzvU0djwoqnpzXIPPyajrrW+x0c7f8HEZDVkIsP1Qk50rBKV+2Os4k1QV
lDYHzp3so68WY7Zc0iMF8jz7gtzC43zu0deUMz6T6sZ7Sya6RSl9WymtRN5LtNJS
Fx/Zyy/noZcR9uYX9ouAUQg5zRYhagp2K7YQ8/3unxS0vL/Gzf4b7ZQwwxOvaR63
roljjBnBwoPdgmbp08XQTkKu5v0T4g/ReA+5KVpQGWDVtaeJj88EBswuOjxNnfQu
JT6RoOY729u6ZS0mnVfNP0plMQNOsor9DCGP4Y/ei+zgF1GFKm5RdrZIOalQG1ZV
T/EgHgcUFEQbScaO/bMyby1XRSlyNlJWnJyyFDE0r2ohuuvGXoQxwETZy+9MnVO/
4GW57DFx+fJZylIazReS8lx33/COt1jaduNKaE+bdRIzLlwL4IT6io1cHCgB20Uo
BR2TWa3sIkIWYBpoRAQVrqF4RR61IPUaS95UH94dCqubCu8TMHIun85qPvKOS00U
W1d/CBOV+150c3RJUEjlhXxGvO1Q5ehB7Y7dbsxWe9OEvlXGwdyKeY2I8vOCaSk+
iZEIUn6SwlBLtflHC8xtKd0qoMhBOLqwrEhbQyVjNUXlUyBRbTDDjKDicpa5aIV0
xRppBykGDZFk53g4pXUP5uuQAk02S1gLNX3NutveInxuRQF499hvSvb0oIwJxpV8
T+iSt28wsffQt0wVaAwpg2eYz+nIA1uRT8DtWo0ymVB4ZwmTr2xfZkGaUaueXu8V
8blwcOcNz9RrtFv+UUEcxVtwm7ManuOr2Zldg5MPPbSguwjWx14Ikd41CYYSXR/0
f7YmNfOz/6fwxs+yuPafAw3bHg+vcOJGPN+UpZwRFRwZ+sC1FEuIveGmd0tCBnnq
urx54JgupFQ9/U2wpi6jLU5Lm7pK3Eh5eBPpVJCVd82XTEvPDKmcJ8lBdplL0NXx
9Gl3s+KiBXeNACKopTEm4EcKQ9Y9Xu2v2+9b7i0WVpjjE8ZIjFUF0No8O6ACvwPS
wDC+Q+tpyqKNtibPNQuLdpgbafK/lLE0E7foXEKPQhk9/kwFH30hSYtrvBLGmGiS
WI+lhrAUVZbg0OE/WCXJilCpt2U0hWyVZaaNcyL5pipBylG06wVheK2SzNg/1d1Z
gErPGzsK0B6SpdR7JcupOmu/eQLInlkR9cqzr1zYCybTghGUSm8i0KJBI2YzT4l4
P/oUECAAJrD8mPBtKE3oQbpzT15XGn7+2HPar16ICchk0IIM0ePc+Ek5m4330kiN
YXGYLR0ahAKRq2j1iCZBeIOYYlP11oZWziN7Janm2jiAXoEMJDTA8kAEm0ytt09i
De7Vu4g9i4lt/VePicjE7PoVoCVd8I9VYc8+l1NjhXoiPPx9Owkgr7Js2PnMdJcX
DysyPc3JZ0P3kfHmkDXhCST9LcTykkux8oEw/8JCmfiL/vVMCbD4UqrzgtlYbYTf
ai9sE/1VClUMp1VT3igp7vHlbgPkAnNkJRha54U7LpBe+ji+MbggkL3wdakWgsUT
vy6N+e7J85gUNuNe7hJaHm42mTxoD07+q/AVmRTzCig8jd0hmv+ouWUTJ0/tMt0m
6rTlMHGLmiKSF5xvKNGg4JnMeOoOuqCn3aq0djnxJuR/u9ptGUK9gqtyXPaqjELj
ReXP5xKSiCGxiqlHo+J2clW39SCQEKgqfEfnbu7sKEV7d8WPJE/fD+55o63yNeva
oy8C/gRlICgD/5YOExHPsnh9NxtlOoDcBwcXRpUx2l/yWfsnz+LjeazrsRk8It/U
Csv9j+ZebfM5ZUJ5oSIvxPJg4pBn4iA+qThb1ZYQwH9hMT/4lut+Rl4q1HimXJSt
KBYnqyjZPqIuQ2SiOexovIH5ROB4J4WElqMzp62rLybtJUxjfUfjP57jBOWqZLkb
s+71GqvJVhcgaQ4HXcD7NNgg6R+6JBOYhfkRvnfIIrt+YhmINMa5jSnJXFvyjkIF
V47Y9K6C/q1YSR2uqaewIBRP5lTawzjg3SjK3NlDY7WpPVH+bSrUlRgM+e/D2R+D
IZwtM/Z/XEiitqG54bkCEYznnT4IxC9U3zLGoo5PQEiStd4/cMKyignrNi5IGCZh
ZGRVXv6wlzKQw3toiiNmKhBc0qFd0vkvkNH9XTM5F1tQy28nZF/VuM+gIpWaUo6M
+0+AGZS3jQMo7sHjOeI/5hZCC1YgigZ/y85KL7/Ok4jw0CxghF5tG5L+EliYM1AE
iSxVuHql5iJs+bcu5WSzRN9yy8aTsqz2Y/Q5agmYLUtQHxqVj/4PuHRlnu2WoMwC
kMOKuaHXd2xAt5WF9EBaMs5Pz/nSi82tx7Kl2OXlnn+P/f1CgpFrPwdHen6GC25E
jlGFM8UBDnhG8/kG8ilgEMuG9TLpvkpd7SCvb8o1F3RqrCqgRv7ixJvYRCGnjfUJ
TIZnMYb33D9DG31eEZhJJl67XYqa3irYv2U0h/aSunDW+BQ6xg5bKX2C9PgoaOnm
iUvMl31TaHvs8RCbYmDdWvct5MhLIFxuRhSrmsP19AYhxqI6BanxMDFGAXR/bIP8
qfXSkK8S0qtSYvtvCGUxOHEL78hlxCQk2MDSUe6WPTaRtLekWPmpgn341oegB4p2
qAIXiHSPaFG0/lEHQKPj/czGNY5nOW5cDgs8n0kTmIWDGyrdtiV67YMZef/A/xNK
l8Xcrt+m6s0Iw0bwqMG2ySvKYEF0qzq7pRuK2zyRTRW4C5vvPudR2fki4TFdLNl2
L/uWKMT7q1xn9Om/0ltCJfu1jH9j8YI9FIWaEQeezGi3MlCgsqUMhV5NclF/nxGE
IHgJVBQUgHmVTx1uPazeo9dR6U99mdY/d646x0tnrFcebR4VJQMd3WlN01f3q3nJ
8hweVkG7NZpmsL4l/7+vuXjardo0eus/23Q8llGFIJVV2nGj7te35LTm3YnIb3CN
6hCebcTEig0ZXya1De1fAAQ1xwyQBKo40/5f/MzYgwaZ+zbk3BOdOfJPrD/AeJxy
06yXUz0TeVKDusOYpn/xsB5wTK2relhlZm8vx5rTpgN51Z4waTQGuk6HEnIy50NQ
MZGlNpBXJMgHoxtAhc74Ufs3kG7PWsN90fE8ljYjygtQgwQpsF5Xp9Lq/KVTo6lJ
JUee6ytJQ8+3OWwCeevOVLVM1GDHWGBDvHNkaPiOernGNLIAjb7JOxL/hJ6Lia+P
s4az0mqnWY1QRp08WAhKhSQzCjvFulR7bMhMoqfnqdWqsEnuYkVWH5byRIHP958B
tkyHIFHSuxw+iNv7JhdqsAd0uv9ekO6+jXr2cv/SFOXf+kxl7gPMfKc0CeycHiic
kXLLyBUJuYCBGfr5lpmX7QC1FVNGkaPj4c4GpAiFmEyYDRkOJjqX30Arcm/VFWgj
ZFFkOe8MuBAMqrvPDDPSekkrpzUI1MIaXX8sR5tNOAyRChfssCo0mhiiDtsDWJ9e
eabkYnc8BfTJh7df/piOygXxjNdPmQPP6E8YPGdTfg2r6WtkSQBKHKJ4t7hd21yu
OaH7dMtRQIk9oFfelMU0VjVCDoH0L3AYdb4XJtqftYmv34CmzjxzFlUax5TwdgCH
rfG2mDbfty3VpaBMEkWwvN+eFxltgit0MRqdZmD+s5kHRtX6RxiyitlSwPMlACgZ
me9hbbX7sBC5kP7s34HgD/pzHdI3gyU2HAW/fgQoVmuz8u5GSiXIXn1QxDkJ3+Od
XviLYd9dqxqcHDzXf5u5SEsxA1/IKu//sKViErlG5Q5MnaoBW/rTcwgFKnCwQ/ug
AVAoEQiWd9QOXVFHRlOepZO8shHdcUc+peMFm88WnJji7QbPp02/qxzDzhajAR+m
ChKHl/vTmSkfN6gtMUwGTl8VYjkd4QNtDizfZeodQJ7hOZbkXflh+T0tKhK0CfAx
6s3uZ7rU7+qRcjZGLdiChNOpJQwLtjQGEN9SmzhSxg21aoYR/1YCdkjUQpSzdJlu
prkdAhrwXT5okICyGNVyVHbjFbl3P90klXjCEEWjaAunW0xV8zNLMXxuhQy/vtjF
Y9FfEb6TgSmHRAu3594vLEJgRofV/mmJ//Um21Js0oQPZy/2z9gsVKeEWv3jWCsU
Zxu4T75pvdHNp5Fi/uirHmTXT1/Lr2IAfZp3w968j0+HzbZ83wAXDBUM/cbUOt68
5MQQZIggUczzWdz25MYb1g1hs68BjyTdg7yvEmnKzxQ3icrxegAjgmju0L25P1SE
dUG8RxIL2LFHc4IN6i6HmFVcg4J35GKtmA9QiGFAeY87qXwsRheuPMDnPTKEIdCI
16MVO/PNvzeg7A+tD04IFbu++luAiAFsuXwcTZxq0tTefy2XcgHSTd4gQIyVh9zu
khRhIdkPXxmz/PJeT7OtGlV9zwKFHIX1Z9KpFWZmkUG4Q1x3GRxPxOeUyiccGPs8
8CNbKA4hwYACRbryRfZQuUfbEsUsCkPXCsPq8QI1RSYR2FXFN68C6sPnrX1iqIrk
PEiVbVM5qG5DIs9EKWTNVwGP49QkkBReBNlXaXl/yVrXhBnAzpfX80APdBVkUQ5m
WKNQpaamb8CQv5aQ3zVQkrJc7cscF00uh7BPGJUoPS4HrmrxYHUS0I6JZfRk6hX9
iH10tvqkA4A3JYEyZMKWAxqheMDf5lHbBazk3p4wNi2QjkE3WT5qtL1wUtx7qE4Z
DTg/SznX8e44atBLaprRO/w3uvRztLdG6EqYH7IuLXSzca+Nj7TOoigjwgPoscYH
BMcsL+bhnjNJmc/yRF4ZyNap0MoRucXoU1Ag2HHjeLvUKuDDLiCjuoj+aPsCnmHl
mKDU3+QLceK3tBP2L3qVFs45bgdf2QsIFdt5jtvwzbR6oynLiAwM8HHULCptEa6t
QFJzlQWslEPXehgalRWAUV4LBW5MchNwSJ+VJmY1QsXnlKDbfzc53I53kWVPjobD
DnmClObuR/iUxdB02nP5HNiSK5CVcLXICfx8xnjwdBUiUyaOj0G1wv2J7vgz6GCq
XMq1Tt5uHcxM/II4fKebGQGRxpoOMUf3NXd+If5r5MlxMqj6vUuTHh98esCwNAk+
J5uFvma8ox5+Q6e64dnFA6xdivm63Ig8hwE5ATIZwc7BXXBY/ERHvyk6MyJBdMkz
5xwUZXUmpNSJwhngkx6ETEVCu7qzJ74jupOEldnZmHovr6ua4iPPp00rIUWS5K3p
ZNvhL1/6Fu5iSgD9R+YJyfH7HHS17x/hv4vvJ/zj8MqVyfMvSgwF+GWbJqZLSz/W
wiJ4bBuSqd15yDm6F3ss3Uyu/oR2gZdiSDAxJUX2NgEpYoq7fbnLCKi62NU2MODL
b+8UeTkeloKBGRLPd8Sih5ZS2SNAZlc0IinyDxrgg7jmPRK+E0eXKj0OzJwhg85d
0rRrz9+2PksVlOSenzilxFOoPyobQ2EjlZTMFLlJYf6Yg46xfA2L8O8MN+k5FUuF
bUiq9OouR2aLIrPHmBbeBB8hlCQih6hpyyJwLCHQyYV8durXBuaEAbJldmyiFA51
fM9HrDRQpzb8ta9+s+G6oqOLNGpS9HpErJujzgT3f5ecIBD0+bdHilKaVd3fFsnL
xzQ9lhC2c6yUgG+oxehVw+Fv0ju1VS0GZOGBltIhuGfVYX7cYm7R6dTYsScFdP0X
z2fiUTE8TxLTo/eY8xqhfD8PLGDCF0eO6zRcaDhS0Ebm4Dl9aG4Z1mwiLNOsz3ob
pFEuxw/l6gH4sA6c8SeZBDvgxdcOraLRF9Jkd/7bqFchbK/PdShgyrfE3IzIOa9Q
DBqWyrMwbFy7JPwfO635x/JsO0BzBHKx3IMs1m6zaJWLJ/N4s6M1ZCSJ6fxFgLSi
nYIEJQxCJB0O8xc8P+i3IA5YMkeEo2Xj1IGt2eJnq9rWCqExVqkFlWH1k6MHsLvH
sas9zj8aDuriopb0DmVa9wvJGvaBr12YyCABcKn2RcaiQw74d8Rm7xGeHF4siaeF
KD2A4H5y1so4Z+sxUsqVa6DZGbQ9pRQerhq051F6TK47OXMf0+pVSoS2byhGB+yV
dzrylvkUkC8MG6P3xLZDhbdG8Bzxcuov2O+avQen3HLayk7C3O5RdVF4xAyHvatd
feBijturUnHTg+CoTcO5DuYkDjsu485nCpitPn3oH9lQP6kOx3T2j5+/HrmSX3MT
AIsPn77Z5JH555vm+L7W6OUVpe27pRtZ6DDxbLgbQHN9iVyI45UQScy3+dYSJqeb
BJwxVqovI/A/mAsxjbIt56qOudQ7xg+KG1mcLmGB+LmkYi3A4RdgtZ8gKHg7mnti
8gnEGSa8sjsg1q03qGGTWfuOai1ms9Dr2RKIajmMh749GJhcV6mmM4ruxbPVOP8D
Cn5KEAn+wgz2uygW8GY1w5NwzN7wGuAeCeRns7C95hMkZL2ZQ7ve1rK6uOp6SaFJ
KN2DQYcz/HwWbUbsBng+ME+hxJile3w7w+3kTWl4W47SHdIbBHpQYb6WtPQAdU6v
OnoXx3B0xJ6bSRfvV7US4XRZ4AFIw5v73+ZjlEo6DBjytIM7RDCBRzXIIuBMS5e9
ntU2Exc12pC4Yazk/EjA/tuOaeTtSID6NNNmBZFXIoPK8tJPS708DRvz+cYFCgPP
8pHRR8jB7agrhrCLnBmIfhA9LQ6FvFbBxuQN8bm4p/1WiI8UdJd4YNDn6XGh4W2L
hK0DaSRn6z5SbwGLr9gthjz6wIpMY0lFsO1ma5+V4SHoPGru4XPNGEmNOqTfHYf7
TCjFGcGIej5tuNJp6Y3PqUentQiaSrb2Pcbe4UmAvX8SKQmL3YS9ezltPTUISZJt
8tRo58fqrdnlCSHPumQXmIGq63RSvcH233uonsUqjaKKTDBlkzHkX5pJnzbyXkfU
Hp4z+wCVS2M5L2AjVJdFTzJY2AdTUvV0vAFmJZDE/MwX+QFQ5Bms+mW9tuKuK2Ap
MFuILA7a7K00Apn4u2QNn5HAhIt3DuzR5NH3ylR1xZmcw6R9N8fSfSjO8pP2RuKq
lB6s4DZHn0NFtDDdqBrCsQeF5fZksm+w7kZv8lGnomzLxd26DNGj8eZoyvvVL/VQ
LcyTbILb5x1BYdRkzqG5EMnSWSU9ftawzEFsb1eHDl6BAA81Gcai9dNvcc4Sl+sB
LrmRRB3fkj4tAKbB+oeTEJCS3s3HmSCcD9aLO1JV3NUDX68M5tmklCDSHbYjUloO
RpcaMLDBX7vDfv/caIS8om52bWU1+7BE9WyP31tGRUASEp8w+xTmSjezJ6442ncz
WfDTUc51b6iqyJERgd3eeOFZrEegsq9VroD/L64DLBSV/1WxLbTp+rWmEsr6LO6a
5l/9WMO458HXc1K6sJQTiG3HJZis1c0YtIMhy363ISLvf9v6fT3yIlEHHvA3gd+i
YpRudS7F0N1DoKHYBk8HqdJjA0OWNRgvDujacNuHvfsdvJhudNzJdyaJ8XoPleUF
D32E0haQ10xbK1KUdn7yf37wIXdEiC40nJl8p0fexKr67n/4X4WsajE2CV4A6bLk
XMOqgvI7Wr7M9tEjna9Yqa7nAiBnGSVMsKSX0sLzM8Ce6rNy4y4ERfYD5+VMjlpN
iq/X2+/gWNkUVIlTAxRnMm7gc+BOuQ2rDGyCHe6FBHKN9Vhr+HNnA3K0mjrz3NMm
Yf8ZKTf7ikEnoa3lt+lFrAbWmGCjDAFHnt47EcjBkLoYFwozo5+fDln0Wvn7cYBE
XU+6VU4mwKzRLbKbB1+Ljr4dCLGZ9ZsM5uZAHAdQi+OPN+KvT1CG/1bmqNSgEKv3
wy8Y518om/O7CMVfUvvQUP/ogrn8xWy7moEB1gduupBUDOCtMtIfEY8XQHaG4SAL
R5vXUXKpcXcx3YKXrnIj03uTBK2/V+O2z4aJ029vwUKpQ9Oct4/k7rb79WWjaMaL
Vgw2vkT364FzCj4AYL9Q5xX83DVDPC9arDalFXzxOXtewUsg61tnavcgMw1cngRj
UPoQ9ZPmbxjiMwdizpfqONxpQoiirACrbjdw75mHbKjYmuaB64/T6kKhD0TEqMxC
WpQZ5Kk3aCYrXomMApx0Cc6oVuUXGfIYwp4M0yEoaZeF6ditV3n6icGO51PJ/GQu
AyJWlCN5aZ7da9AKwqKlrunDGU2i1MBHSfDSuWGZz2QiecC5qoQwSHy57abTIW1P
9w/UVn11uWZX6UF1J69vwzS57DZGXdJhmip/h9LSeR5twnPa/wsdciRJyby9VIlP
Efj7oMpA3ubR6lf3drd6hQOpl+L27wZqdBgpZUEwTGJCQkdBcCIdhtZRATYGRFxG
+bkdWvaFInwHytPAfl7VtL3PT4WCFsP4NVJuby4yP08FnFQpYbpEwe8Pi5EEALpg
IBf5knFQ2bD+Hws9kzx6fUIRh6+9vcMiLZnRQv1r3G6M1hpNL7Vay35BpLoEAHqt
JNYF2K1NkgVoB8SP28you2+zJljuFAkeYt8fpUjNCW7o7VAzj6UZchUWxTvJCqZ6
PTtLdwcAS0au79HNrKVwCnKbYTkKRzVBaaBPBsBBOejRZmAP6ghpaFVnAOdo94cn
wi51aUerl60FIbooo1pnaIXvX9VoAue1F5ABaGcjX0+fy2cTgLBb0W/cM/A8WWLb
b/ya6TU270mHxA2LPpe1ygQVxV4RllDmVPX71KHW3xs+FzcXkhWvYHkX0KwYyw7g
WszJIq7YBwUiaH7a4uxORtbczIEJGXl6QnUCCuemzTbQWpfDYELUNdyRVHX/QcOB
FcRlMwpGXOJFrPzBgegYpdsAyHOR2pzZuoEUW36ymb5pmexnifAVmXxIvbLlSfHc
9+wWGqG4JD1AtCQnohsq6EC0TZCR1npHTg9d4dAt8RJWqIWumJT0fnWYtXfcBJAo
p6KlCvJr/jvoZeAsbbDHj3/29jbSoO0M5LyNX0b3JyPDtbnmMfEZVFEAz4tm6dDy
fK3V6OBY/Kr7gkzkpV/4VzDOzcXuCwpxh+XGznQVOCMgDqIOJRNAgEHBhtAJd8ZZ
MEPUiNCPxfQyKPXaFB6rZ2aPp3/qUMP5oMa9DGiCHZH5ZsAq8TGZaqwplCzNV5xh
QR5K6gnu53ZS+QCMj/36DBBsUFBp2J0QPZNgwGaah6/B0ArcSuK+NrSaXGrO27oj
HC+7VdO/rMMcCM/92z9X1GUMVQFmbmJGDiWd+OdwI+5U5qRAkGu7ujCF0OdgkWZp
I5VIWMuloHO1QhDFomE7+WrF//sBs1uagG5ONHCUA2+g2hJH0vz4SKVk5DkNrtIP
+tR6V1x7qPFMHVn7cy/mPQAqiL2bCyxvp0CTvee1tjqows5Tu8BvUNtVaSMk5D5G
QDLBD2l8z4Y7T1mvYlujgpAbCOrI62w8r6rhyaWBC9ZM19YV0dP3zuinYvg4zlC8
kHoytRRGkaOadj5pNSbaWSVtWwElQ3q8sTpKmPNCpHMzhDArBVPZxDRD6eBdyp3T
SMQfZHnI6ZxAOW4cAyvZGFpoOAu39U+efxBLN7gRQ8qk0QLjPeFYB/tRa+y+FGiQ
/JGL7sylxVJStUWj2oXsYFDf4omiWXAfAkrjh55v5K+ZMbJkulXul4rTywvKfk21
mhCnxacu5vrUKi26WBS6Ua4JjNdcqpupW6zuYOAdqJYAcs0YmNBajWOSB0XJHiwS
eItmo7BxSJ6FxI9nRdLFs/vhsHT00ebC3RlwMYVgQTRQUzGnzA16Bo5FvJXaHreJ
W7GdnF9vFZ7ydCsZnxYJuXxlaY7sRncGS1zVUy4VFHQ319v3A4NHnH7HvA9bntI0
4t4BzOpwhj0oacz4HtBU8R0AWDuM+HmmYmQBw0tTqoOWQOkRqu7zbdDlxpD8mAR5
CEBYlB3jfYcJW3wd9W42/LUIBaJBqM7STfk376fIXUPbQuURXdWm8x5EycR9lexd
JvojL9CF9dLeVmoJaJsUzVul674U7RFejGGicF5QSg8INGDxumTF9pgLv78Nlwq1
Xz0RsoiRFlrPvMEoSC5GJogtdgDfQ5+If5EbHOoKGOGNG57NCvrJ4nqvL+lOnArx
PHI6uWYzT46GIkRuAejXmTkzi0ICBw15B5gSQcVN1n88UHuPQaX4ET/hk/GVBX81
HU0kXKfYL3uZGFoasoD7/7HXtaGnAl0Z5Guw43toM/hNouG8I9R8+HIjm2kPQl9m
yAWG0oxmSM7WWJ54rrnPo7mPKwxIhcgZ+XdV53viD2ZiXhwR14z1mvayMa6pVmC3
MNnco53JGL/pV3Gc6w2bJnjRcv9q1tahxuzrAMfjLokeNfASaVVYoNwaMG+xgCaf
YX4ar1BY8NqVFLhz2uhxD4rmhtuVld9IurqcbJtAYEqUKCrlG1GKvbf19KLgVCHD
/inyDjOQwUJr+Gj3cMzCFK1ek3MUhic7umt0vMZf1jEFY8XSDCEJJJ2ryVUd3+Uj
7P+146X8sMbvCcfGq31eEx733U0rrCC7QcWghqOyiOxuhWxu9p6Hb7lGOcogtq8F
a3wIiyrJrSKo2Q4mQmgZlNpr6mVWH7lDYxGWrHLDCA0F80EquZ+0rtHLhQ+foqZf
9J3R8e9Bm2ZrcM//m6F+fdMN61yeMLdLNtPGNoH5gX21x7vwFZ3/0hL4oaLxO3In
vCR4KbIaMl4HiWk5ePd2mcTbUDPNqWKfRmPPVrHTIsXXUM8ELDisxxBNBalQ0el7
45TPhET8yvy3+Sb3xnCLa7bj14dl0ObLX6TkTN49faswfEi+mTnIQk8W4GSsg+/s
e5qkudgD7Ep4nBuewOiVlk041Qagul808kCqGxmToT6GC+up8dhOwvcIInxbhbI4
hQqLFQKxlSabpWrtYZyEX9F+BMvF9aA/wWLdhMYpNLgalvc8dDXhHdPOjelpSOFg
fnCB1RAlGKPplF1lCc388tEsupTKfnjziy7Xbr+DumYNBxks7X/PkYEdFpAGK4N9
jr+omnjvC7o0RR0GzeRJYbfGjPqZfI5rE0UThDnDu3J2FfTa8bUrCzAY0dWo5Xt9
HnfmqnEUNKq1kxfF8yzR3gaa8zZH/FZNFvyEcaB3PnLjrV8eVeTi+oqYxE8iR1Xy
XhtPT06hz76I1Q1d/Uu1dWC0OmdqWoD+BQ6guEqKIEaJmNRyZvr4y+M1GA56+gxN
Ab6RzjcyTsdTva41fb3q5/07eE+5hfVR8IPJeuNxPrLw5KEshKSYLkRdvgssCypB
YqRrF8kv2ladVw4pgF1bFASUOl2aoRz2leUNIZODfjpIfn6bSIbwv7qH2y7lBck5
reZgsHbjwMCQmwnAKVP8e0ks9BdO4oqDfvqS3qyb93vk2uSZ/Lm99UeeGpeFkUOb
yUjBmU5horJfYDw+99E9JnKKlJS0mzAPWfw78fi+60nEwFKoCV0IkhSZ+kJgPJ9z
x8El/Xy/NeVIln5aVZEgfYD/8o3s9p/jShDIrWTNRT3zC9L4XDrUe0ufMiuDx5O3
v3T7h4PX4cVsTMKWO1IPxjACJy7yC8YyzTon8Ow9KgTQLZCFFYhq38gDLLYzFZil
pOMQyTAqkt/2KbfrBnXaI6usyB8PspdAi0ZnOqMiT1/6KY9Viw2Oqa6TGYAyLuTx
TkV5SoERjGJAyNUkZRqGRm5rgzXCFE90QifXnZBYT72qd8bytTnaQSiACngqRroI
U89+pHSdfLLnkh4k06PNxsmnlE7NDbduNNBeeETXPE0AtlmNdiT+QikDoI4S6avF
ELXJcfpxM5WH97ZlFRKDHvJB7Qtx/9sjGC7D2zqWVFmtkU9YDa3KY3rs1ATebpob
nBeIMWAtZmuXZAWWCqaiVr16ZSne+9pJlgBLmrJ5GX+2ohIMMdTsop27gcjJuehY
hbCET/iW/vi0bvqSlTIPanB+cJ5lGvQDhperSllUjz6p41umPcyChM0i6/MERj9J
5+10SOw/06EcMnnhdNnharVXmkfgL9lPHbkIBAul5mlDWl52t02Yni5aDBIcLwTS
dtxfK3lWnjZXr+HTQFM6RjwcvfJ3VxfV6Atxh2a13ZUkyhZXjkkUtiCZeH9/VAXO
S6QVusJZz+55l732cd1s9gLIqyoHJ2y62Pzv438US0to3Y6fcmEdqxHLooCsSyzX
Xh/k5wSdwQf/DmiB8nBFHSI8oQHxkeBVp4vfnhYvKn+ZD4ujYREx6pKnlPYMT7lJ
lMUE5bxVtQ1IIYzo/tA13I7yBirW2HWxkfE6/eBE016yLbzMTtX/nWvm72b7bxnl
JQqw/cg427HdayHs7utyAgLaLf3RnMcyra3itP8ujWKsW/DMsKhXzt/xKnWoKAF6
CJ0d+yCiK+MwsBMnp81NiD0Qvd0r6DnEPLsTvlYAI74k2jm4HfyQUshJVLUcrRTy
grGTlfiXHYsS5doVhuf6QAS8pxHiwWEQm/wNblIy9FMADcywBLJvNHA3uNeUWmeo
Bf2ZcoKU/sDrC/lnZK2Qh170wP45ZNl1cIFG9aaEO9J/ckRxARyVuYeZwlgXN7sM
jMbLV7XxwTiphNuzVOXPJHS+jcYIUxKkASZqsVmzP2gcDJu0tWcITl4po0IaNW9O
bb+UHrGP8/PsHf1jXWjlavs/hquwc0LJdpLd9s8KrF0GuY7lggLTwTvY23ZmLoj3
dO+L/15htNaeRGiOobh/hDnVeHJIi5CcsvLCoxsJALcClSl6PXTu1gUEUNLajodd
kVRKOm4j0WCm8EsP9dBHpbXIoBatI7k5JcEa26LpIHtOxnzsQR+12Ajcw2GCo2AF
+/iY436ckY0HSr30PQgj0ZS8zgijEKLhY3HmfJT6mvWKvE4H8RmGkhbjLg2AcIPo
lB3i4J92q4onGDl9B7LaL5n6ul1q+Fu062fUONqHKKBtAOxlFqJPbkPBCwT8YwZ9
PamIF99fa7vU1tRLL8FGbiy6KRQEOUSn5GUID7j2VjPv5eq8e6RfyedQNYBlz1Tt
8ifjJlSqDrDAb7sQ6F0tWEYEK9UTW6VOFBTRosZD+Hf1HT7ouq5lIxysmzag7sgj
EGaEiyuEWjBrViv3o0/U1+8wBLFvoslJTWIZmPkoqciYg45YMGPLcOkRpfW2aYAS
K39qpgBKMZgVtc/rb73jnAAbyCqk5KPFUfsFgN/yuQfijSYKF3a+3ocb0iR1uiD/
tPOYqkrICdCpTRcjNgr9G1EnPaSCtKCqjwpl5gTpuGEwwQlOGbxEn9vA1y4Pq5GU
1KdV5p5o5zYbsv4oO/gLS9T8w/3EheP1tC2BfrkLEgIpitr35PKYC42I2mjC6bAh
1fU7IXGPh8OQWjbdXWDbOnOjxwtSWFI6944N0vcLFYXbeH9ROr6dFgVpoE41LZ8i
mgbyR8pvTa6VIObIIMwiwq40SEPFSaKMeHqp/xts+MRoRzRXaIZHFNGGzPAuqH/M
YpDfqn52aEmIsHYjglQho/FnUqCQlaXDMVGmijAIIYTFxxysHIajdU4dIDahA6fR
BD9qucboE32TniJlH692DWHzT5Oa3jblgtHWS4EEdN/A/3SWWV6dUMbxahxQJCfH
r3w4R+O+EeY7hIJmoji958TGOzsoiae7v5HjCQEaMY2yzgZzISoHIv/HjbTF8Ax7
NeHhwrMOF40cKCMX/oB+ot9G2G57KQZHzOdREvPBJGBiJ6qVffR8N4kZVtwKdOrW
G7kNUOz3cgTwIyrxJyviGOu5rZJ4ljQAnFZIThG6DDjw4qgFB8ViT1c1ewzKXMYV
v9pA+vK4g8UUGIetvMbiMgFv7PQKnwLgJYFRIu5oR/dAkm2MDWyT7CXoCT3tWGmF
BuZDQK6/aW0rPx05WtGmhDERgSArsWjnWeANLIEQyPUk0KhFn9GHW3QdTc9aKHCy
3Qqr+RT80+dijWlUvL9y41PQlB2bdURjMDIOgjYMJsLebyVQijfXWzWEnRRVlUai
HYEVZ1l/TP+nP8Bj80Y3SGS0XsEde7Z4oWzCwizrHoGLs4/fp5sOS8ThpHWW1zIP
XvJ8SSwkLNphOH2N9L6VQRxhv5Zz2CI3ZY5E9SiqFKY=
`pragma protect end_protected
