module node_wrapper (
	input clock)