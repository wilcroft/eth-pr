// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:35:01 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GM4QuAO6OtUgdUEM1vXZF3PFjOrAcN4Cyix8N4rb2DyirLDrqmFg9BTQNxh+H9St
dt2yyjY7bIQOU9VhkOrDvujS6lBf6Hz7HElNeiSCIGfpB1hT+tB1Pl4Ahzx05Bac
Wnnmt25czV35kvr3Cofw4e/uGOj7jrHpH4jta+1f4W8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1488)
8/Eblep8r0Zk+2qH7EDvTreCWVjcXVa8kWI76v4L1apxKTB/QngppfT0ENIC+16a
WsQfXqVG6lpkrTgx+EcP6jsR8UlQ/brgW2BAl+iZwTrFbjkjM8DJW7PhvVWwTPjt
JYnB+cej2ZcpGKBzV5vQx+ytn/ZwKx4gv6nFS1A98FdROzjGI0Sb8Ajmd1UvncZD
h1XOQzONvIVquKOEldywnrCBH5ObRwUZsxVNsviaaYYTz+AlpWxGLNDAzMze4+MK
HtK9kFhCdgI13TxVZSywv0aoA/Zb6asnB/219ALwYr8gVs3udbQYRnWt3jqKZL7P
/h0qrH7LNT9uoBblO0/AMroRxiLi9vWuy18qn3tirhcug/QPyAyqvXmZlUgnW4fV
ToMKf6lp05bdmZE/elkYqf83qo6PwHTKq+O4YE0fQNN4PT4bOoK1C+6jusdlJdn4
d21LScQPVshSVnWHZLFNnthX4S2IwFqFT7NLmi7BvmpBctRwI3SrstkxzFVg6AR+
I6XAEw+wEmv0Opv04BEI+1usN/MBnM82jmP1Uynk/Hi/6AXAxWgQkctIujRdNjxB
4BKQ8c9CssgANYmD4M1p2wLD1HD/XrJWdk+GxrpdkWNyP2c5rTSLlgEyZXCWbsCy
MTCQTxL0s0OsYg6rUGBWokqy8RVi/16372Dx6DUiIOrVf+gCb7uaNVPQ90IslIEX
hQrxN4aWM86r+34GbEOp1uqi8ziyuyr8JNKVqDUke8UXDJCM5sZL7vbaf7QqbLIL
SjirNHGgbh6Wr0bWBeF94vnQ2hmXlAJwAn5bVqbMJrUHJNpWtu4iu/I70XWA2Kxl
cI6klPegJ45prfFV/9us49CA6/96E3x/5lnD1gYlAb1DFPuVBl3mcB9/Xt2xGOzz
QU14jrGOL+ujCC8upAYb7cJD1bajkR5BOd1/GKR+yZoFBTFjgAP+sP61q3tVV3lA
syy/eXjjCBlj9W60ogkwcwboD3V2l06vx4aAd+JAWaFCjmzwmpjlS4YSbXsgANri
NxcxmAVLC1pbBTCPgx/7bHvUKOouNHYzL/EwaaXD/p4jySkNGv/KwqUo04i+xY6m
EmW6k0BhOZIO5aYB16PSDi0H7AlAxSWdrkKO2MHVxb6eawEqB/wsqfjeLk8w2BYq
DEBP4D6NcErt6CS17Qp0FdZIiNg82dXaoynrfG86RFg7EpXNEuJeuK54Q0nc0Yqj
zAKKhBC0RgwOLHjOGC0m92SRyrnboD7vuETqOqeqmdUNOGS5Mp47WS5MAC5pwo/i
Vf6llCgFokF1Ws1VcAPPiXy3MgUTaGjYjySZRT0ltQoHKVtqD/N4LDWnwz0+If+R
sdR8LRiUnBMPyzPSnU/KPU/RTnz3BViX9SfgP8iZoWF/WLKPy8/pfVlcm7vcKory
bvi0LQYCBHZewCMQWU6SJsSWsLIZmVcznq+8RRT5XwaTsSt85BSQadYY1+hjt/kq
bJ+LLjlrHIeaPPUVkeCchCq4VUSHF1Sa5fZwBobJBjMt1N2/rV2Qt56+a9WKoJaN
xaSKQXJOmR+lw1v0dcI92lPJJdhhI2X+v4TwejcPiqsoHcrKZYeK1EGBknQ7vx0r
myggNaUa7/KiCwbot//ke0aSu1T1lI6wIVnODcSpqG1/hgcS7aVo42eemBb/3ad9
guvpmaVbJJlJNB37hsGtkBO7/I5KvjTEygu+PJAhKnVnL2HUaADQp5I3F5OV71NS
18vKao1bcOwaXgxZ2FVADhbmehjbKME4yLcZ4glRLW94mbq6rp7x6kUuiQTzreXk
rMVYl8L1inR8rXY/wFfi1zU/lu7odNpw0i23p37l4t2BfvxbUIiR90maF+Jj410T
LZ/jZWKI054tRebMMbruO1uHDxWCq089XVVFJmVMjbJ6+UVa0ncBSIWu2DYOJEHg
RT/xCkADh5mUui/J7LixTRWe5UGtgynkEolUJ8nxuj6pp6PVTf2EBwR8Nq6X/giK
`pragma protect end_protected
