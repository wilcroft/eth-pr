// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:14 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qYY3zujTLVAroBml+IF2Aywjps4sEJ1i3hQI6CvQ4O4MFXEm6dVEDapgAfiokMnv
Lj1yakKBmoRAhEyr+ydSfoWE8wdAc8D17L3Zxz4/CNiierrxVEfxDkXqWKgMsLRD
sFw8fUe7MdMltcBOmpm6J0E1ZIaR0KW0Lf+FFHHFPYc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19504)
edalMF2i6iWgABjHQW5Il3bnpHzfDJglITUbRLayvVZhQ/sZqX/L41B+6je+00qM
UZtWiLPqdM3ym1NbKbZeRqa/onlUkWiZUnAf3Uo/LvkWOIiNBkEjwgYlTGVg+Ucg
9+OZMtu3i7CSAJofP7/J30dsiRTdOx7cyWHE58IjdSOomL3s3TMxne8BA5yiuf/1
IKD7HLWLmKsqTflkxV08Qm9WBTAj7D4aqgs8UwsBn4queLbGSd5krms0mTNGoRBU
/bZFTVhRBOlBeC4Y5Iq4ccwoB7nUNNbP+uVGAvlB+Kb2Lu/LWHPoxTMbpqkKRFPY
51eQNS7rzG2tcgtA6j9+a9wKd6HeiQ1/gLRB1M/pKVyCvrVYEdxv0gO/HWbUGBot
IsGnqtj+raqibkhao7m00X/hhkOkHEzrdli0/v3wiQBK6r4QDSlX4ETfA4kly+Hu
oW2uLvuXYq8qtklYMKxzvDypZQTaJTbFOUh+nYpff1GcmjjrpszkB+OyOCnLuc2i
xGJKv4ToZGUR8hJ80/IqX+OdqxyoivBru5fWGLvAajXpU+wjDlg60ElAqC24LnI7
/2yfJ0tU+BlLLyiv+HnFe/1sab68/VDOzZd2sNGV46/mBhA2QVKwTbcWGv2kErFm
7MLQ5sf+RORexBp2oaF0+WRyJtSlAXVvNcjgF2xCLI2WKZo/7zXwSyOKcnA9tAh4
+wiMLOe67UbufZEOHxrFBtxqiLNbqZPkG7FnzGKM5quetMDGlWGOWKSY4ZqyAQl6
hMkeGpuTKhy2uGeuvmZXOqTYCPtgymvFw4j5HwN4RaCwotejGBKm2I/BkFvVS+PE
C9q0UP6N5ktr23C4xQsxabHerD+UdVB7US0AErH8WH/qtd2MgYkq2s0Rfit73iNS
rxxY1XnGj3y8CeCDUo8XUt5bMx4ODRJBnpx3+6CBjQsdHzVe0hmtQQUJzjMv3oDj
tqOIHr3yixJfVbgVicqeVkaZESd0rsShbrSbg5LJZ4tFhHh6I9zkQLfo8om3Cbjf
mS0nOqzdDS+nJK2Etz2UmJkXxtDgdTNgaDPvCQPY0IZW6Mly6uz6w59L3P6zXME9
28xOzv0Jy997KQWkFfv7COhUEY1Ef4mhSQHGekgwl0tNt2WHiDv7u4qAHqXPnC+n
2rh+iK+aC9nJFxmcY4uP2IkkfK0KkvEPkOdeqdOpIMZN2pRicK4MEETk2KURxAcf
aAU3mH097gPZIfwfM2bA2Bo5VEZVEHtmoVRR8tQmDsd0xFRz4/pxd+UinTEeevYa
dwVIMd2njij8ye37znhYoF2euqq0OHTHawT8UJQ4YH0bmAEJUoEd7T5+NojqKQ+V
B9hBNHlzQtUh40VkyKGRbnzYXVbuSUS5bq8lNJ4qamWUGT5z4g1hCTc4qScDpaqP
JUfMdZlpaX4k65YTHknIQqn41vRgyrYoMAzFb3gi+dtMryMedqDvkPTZVeLue2rp
bvOAL2BPx+xVCA/4Y8Z+st9bduLOqtDdorxuG38om5jeB7P+uAUHdVTCnTU9DyhN
EkPDpJWFP9JuaMhIW+fs1pZDhPK7At2W14IrEoxreZf3Y4NSZMHLLkUYaH3ygtUT
jILxR7l+9REeYFyyoE6XGaavjjQMe7PyseKhdia7xpvgYIJDpUqt0ShfiATfKpvI
yWHMTlTvov3kBfWrdLHnz4uDuz/CHyfOUaL6q0+pRap4Yd0DpHC3oX3meAjYbOGp
6Pz4ZGHsop+4mEo+KL6T2SVIaY47ly4fhK0IEol4yJX8lzTKq9BqZPqiE5Z8XHUu
vYu9VV8lDKEnrlB2reAxCT7FzpkEOhrYYY5kag7H1XLAPoNGwd2q7qgNzY3MBWBY
zuCHTXHFs+sWUT8OZUGM+liQk5uSQrk3WIIOOQ6dRLQkgiKHhmOAqov56PYHVrW3
MywjBoHjR2yUPpEoLK3jhBdSxvV5Rc8bM95pIZBsUFLiMgXPWaEGtefmEoPS7nkm
F8M9Yj589dXlwAOL7n0Faf/2LzKx0FytKznJ8KYkvZtMhFuh0TRXbXE8DYqnEk+L
KSslUql89wyIJPySixWsv/feou+xfOSD5dgHT7fLfZdvkxhMqC7fJy1DFHxOHYrT
f2lGXBLV2hIPbpKFF9EhXit0NRR9lxT+Dgg3Kbe9QyCliswbZmgFXssjhTU17Aai
vwSi8lx0l2VeCgXBTfvxpGyh/fRPamAhCvBZzw00Bt7NOEwkzy07+Mc5CS1oPRi7
6/M6uS/6H13iuNWT5Tac01Rdt/QslQlOq+Jn6ub6EeZ6XBMMEKUm0tx8C7owJy5m
1YiDHvgOM4KRD+2LUrKK2be8tXJVfWz6gGHMmcAK201W/CACPp4bTOLihbhTWrIm
X9+zqaRHIQL+yhPs91kODUZQVGBlfYiM2POu5iaeLfqfzC7GLmZzYP5DzxESwvxB
cLIz2ZOyEV+QczeEkTWQMV6nFE4V0lY7zr4+lwyqMzBV5+mnnbW40dmVvasfOFgM
JMNl5O2zlVGRxYNTojy7kj1wRgCTiDVoPFKjg6L+/kHjIX7EVO/6W8PIWUfBXtkL
vh9/pwKkpCwFnrFqdCvQ29Z04f6KbZfYbFOyD1Jg7npvT3lZUwoHWUVx+zPVXcH7
f+IaOxE1x7NGqXMD1iDVOXPpLve3bdSCRiKBfUQ6fYa1FSGMz+nKEEmZz8ssI3nV
8oYpDTKLJCkSpvHE+tkygYTLO+RfkjNL9/ATcthFSJpxjR01Ti1BRgjYceMw0xnI
ZhpY4anncsyyhpQxHJAKkFl/Bl6BrGS8eL7nJHnXH8zkblVFkCNps1eKxgh2vmL0
ueXmabzZxQzr+hEsZ0IBFfSwqhOnACDKp3FWBhEteeUYEcVWViMLa8oHZTKnRWDj
o+e8h2t+UFncExikebzQTvkf9EaKES1wP+63K0Xe1Y1zK7uSbAKhiQooplY6NFgT
EQn9p+pBxWenn9/6UVL/s86Dk94y69Plx07ycXnacgOy4JEKUfWqZz6NDhiGMwxy
P9IOMK4YuCpgDrrAYNZTdVOrs+0SWGHM7AyNP9KkG8g/cLOHgq7c8PSysW2JBB+O
p2h64kPOKT/4iFKNYfWsOi+DKXgiaCgw4LzrbctN/yo2SvfGt/VofeC1aFNSiU/O
c7zbj74l/aYJ6BIE4Ae5pLZOSh0XvHe4271UL4aypjN+MixHSS11t0aTTm5/VFo4
UYK2xkjS5PSYPv7DtMBafimmXV1QfcrqMQy0VaKgKbpNRNl0CKUv1JTBoyUVQy6a
ogpqu7kOchVrJ0Rd2MjAxwq5ROPoU2Mqmih1TGpoI5WGznS3DrOla42LKv8R1ECq
lYr8R6imPI7QU3DqnwNHNUM1NoIzONLXJVLG9arPtNkpc38FQuGKMM6N3ay1WLAb
rOcPMmcgwVfFrwTeMyjBDTI9vo8iogzC/MB5yHd4dwfI2rsgkyyRXzkS33YJdhP5
x1W3TFnNMskCSphnuGpVkCitIU/yLAgmR/0P/GIdbnlAWqsryMWNNOtQtw5QLGU9
qKmO7+NaWOLhiudM6yegI1PwgsiibPm+hYLt/lczAVV46HhR0aKHyXg3eyNhNtnf
pqQDXxgwc7nABFjAFM5S+x13NPj3NFlcchtQETZvmLTpdHzz68YuoGKPKitqDeRD
LrWAsyZ7RLUv/dgu9+LBpjaGzdZUIup11kQJJyx/uC/mKHG2tWWlfxKMgSz6o8tO
pQIjuDsVivZWG+6L9UvU8EqTINdUHOsTwoy/PtfHm4uQw/4Rt6ewfpuxrs4mKET6
C5VxhIjZ7AHlNRLDumulAvp5bPxEb9fRnsnhtHYju2KbKwTh4TS8El+ahfn2T/Hl
wZtOfRwqtctz0Qi6acv0JN75WcB4zXOVKvZfxKFTRzilCOIzt03PX1/3t/Y0EfnY
EaPHM9LIprWsEXmtIvEYeU6X4V/1LJMoRnQ4dJ0iMc/XZrkncyVR4nQGTknj1DuL
QJ1H2TBF0TQEjBryhVmNfOY2iny+A2F4DvX4TxuIUC96R8cM1qI9YiiwgVyo+NcA
ZFgy//Kg3EoCCj1pI3+CnjLvTxVo5Oy68dRCuhkoWpvrqZgZBJAJ6Tjm/saY/2SS
wX3/C35q8VRzUeOs4t9fBa0PtDvfcZWBl6c0X7nJWybfw3H3wsLsNfgnEYV/tP1D
cT61kE9uuG2qOhw3HyMJZFHPAo4AU7tBHlsQT/RAMsNCps0ub9f0emiMuIQkks19
VS0DpeAbG9+GacoSl9bJ+QgJ3XNkziZyy9LawfPIud0H0Ms0gXzGyxgpQlMfy1Q5
CmAt/QWBqHpH4ildutTjYbcP2X3V6Jzk5G/eE7v4H7+4PawDB6VqHSwSk0Eg8QmT
WPLzPwTFOWaSZqjkDRvTr7hNx8prlMU4bolNaNu17TwZNm8Ow5bfRx3jp34y3cyG
wyC20x33purtDD4e6/ebdXfgKs4+e2noAPn+s0yVT3p7sC1IXKYAXra3Y1BM7iZg
U6wQroTzDPgtpv01Gl2Tg6Sf4UKWj89p2U1PoMu4QgGquFdYnHct/daXawi6OTlS
bqBHIAwnkxmVPnRynKKrwIFn+EVId6oqiYk1u7Y4vM3xI0YKDLc4Z1CfJTGwXVjC
JKPL3SJdru3ZK5avOrtL6keWM/9r6auWiDd6R07PJoCMCOfARNoOwMVDMR/eo9IW
vkERJs9KLBFsun+4yAiusKief9Sp3E2oTlExMnSqY3Pp/xYeJ7+pAciUsK7sUOy5
lYayVJB5fF6Ho58GEGCqmwwGnnsW1SvvZ3SVFcQUmSiGQfIupCx0iiOkvgTOilf6
ejfXMlpgddE8ZeB+3w2wTHusXZP4EovTahg39UkPuKLMqXm7HKyClllX82eJnqkp
AKKEtko/3VsGGKtIvyeR8Vqb7E4qw2r+5TPUvKNNntKB4tmEmUuHCqBwEWnB1sDo
yjB1K8nfTdqzgrUborl8o/rnKihDsc/qoADp6n2qDw6/9NwwbrHgRSQMtI0mmzrq
3luOzDJIR6qjgGmB1MHufXdxTIWUfYbxNfhPW8V1SJqq3HfVg+29v/eM0Waxh9gY
NCXiBxCcVQBY8tJUJZ4tpQIsVce9QNfC5EQTSrtZG501vIFf2b/EFQgl4mvJ5mEd
zGIUmZhxjW9xiS1A+XWb3BWbD0+shdi8SL0Awl2/zwciae3lvbKiVad0InbEaueO
KJRLZPunJP5QaIhJZb6S4rRy0YbjvNV8sqLi6sEyNHdYJJRmExSl3UC0wuMqW9tz
C/U2iWAAXqaf2dCVGNeKBZPwsNbwz/SZox41KTbaMiezSZvY/V7MArSXFJI1DQox
6jLZ0Pz+oNcvq6d3XUAGTdgCdOYNHijY4ak/5X0TFwVHngP7xOMbuSw2c4vrWkKh
WK5TR7VAyYmtnoNNaii31Z/Ww11DngPzQ2YcAfpKEmms6E5rK2zw6PpMgAYLIxcI
T4zeRb4K5o8Wgparq4rJ6VFZNLRQvy7KBuGoHoDLsjVVh1b8wC7d5PZO6M/uT+TE
BErFBwj31QmA4KufZFa+VWk3fzV59/72T8+a+xZAhuP9BCSnLYECPS8JcWZQ1J+p
5dR8heeq1ONfqPFSwpSHnwquwyM/NmKWQHE8UIBB1ihMIRKdxEDsXrl2dP5ebp7C
c8o43Kz86Lqf22ty/YF+pKdRXmJgV35cXIG5osYf/3ctIRVIC4bUfkELPSxHfGl8
EUhI/gTQVp9X6wYAckSyCiBF4dlUD9kSsSwG9Q7vjfuhxL1ToAbTZ3Mp1tK9qcFR
C+TT9QuwfLKzzsZv1Xu44w5FJBVe4QAWC6A6YQosJ/9Dk5Wc7cSaGRUJz6eJrKsz
e2yn+i7FQssjy2//A5pY6QcEgO6OUwnfEv3bdfVtJsw5nwiyf+6PJKNEV0Oc7Ppe
A5TcrE9cvlC8aQOlAW9I4Mcbf/crfNne5fwqkPjVnypDqFw4vi6pSUINNWWkVHGD
UDr1jvm0zZsiw+LfZDyxxBKdtdwZdZdAxBLj4km+EWQiWNpCATR+z9jll5ngNIUY
89/RTeLPOVqrr8t2fTKBZO165f/JYtkX/BxalxlTXBWQd0jxv9umbrqM8PKGTNxv
o72uBFxe2rZU7WQ2EKbKWePc8fohi3giKTcJLBuY8uJOEQAnDGN4v+0o8Mg17TmH
d6qUNeJS3w10ijjvlseTSHmwwSUGf0VfdEFdY4Rx6Vvnw2VPmM53ZffZ2aLIuLpm
pZCjhs6+060cykBSFcfJQNVrJF3RGKbPafAQ3TkyEplI2z91wCnnuaVZsJRJaG4d
Ih6C1wvWqB1VzbYjyagcdHoDHBBLZj/dFR5U+DpM51HQxAIC83GlrnDO3huI+ouJ
HIHx7V1PWi/DJUEXp+6JkLz1CR561JWXN3Mkt+il252dbqO9BG1bdt7sal4AWtcw
rJFzbcJh7DG91kzw86FQ38NBqefCW/7NuJdvO1y7xPJvJgXHqTQg7mvLewBnIf1y
DZmIJOkMLGLU+TooFr9WSfbq6x9KPdD3RcoEbbPkSxSKNgYmB0ymWbu4UdwiWprW
ZPvXrCSl/Tj3remMLncrBt+NzoDaL3iQmPWLi4FB5LwDmjTpRCJw0GuRwtWFbnds
sFdHpwubqbKS4b8EYxMk4fNsExLt+mQMDb4yf39q3/l/meTUiPprLzpK08o8O6VW
jqx7xgyqR3GHD6k8xe7QEGnLnYver2w9DVSdfZjOoTFGkRD+mlb7JNtMMVgJRtQv
4NjcpT+frySZPiV1RT4hkRODf9L2RnIBQ9lEXDQWJTm8sCDC2sQOz2ZMFt2lxnp/
B7vF4gfDG12v1078akklRTk3ADMsAcRSvfGPOACANKWQ7tzSSxR3K9BLeUzB+cT+
AB+Y/mDkIyNBk/EOfODvmtrS5XJHFcL3xEgN51ojeHO/sQxxNvbXuVmHeX1U0uIA
MPg5B2y36cCIg1laD31X7Xnt3nHTuO1gs/LJLn/7sxzFDY3pgX3iBZ0IuzqoPm07
uFW9mx61pIAnsgiiefe5Ednkakzhe9VvIa2pXGk5N5gN0lBa4oRoYU4CAwWFwRDd
kzZ6ex+QkDNj2JbWsM54CmoasC/7InzQ9BdZOisEtpM3+v8Y9bekWaMObGN/lC1/
dcHPVThnIq8JZJ/osDqk3TuJVmABaHPpW49smFUFd2WNGOk9zz/98kXA/J0I2+hA
+oek3qyLNlL9H3V5ad9A3YCLeEPtkujZ43W4vNeiGCibumDWpFLE7CDzBMWLp7pK
ddDhNzi7CbqlKZilD3eNoqFoyDhxfTk6++NMaEcjfXBJ03kQ/LAoro3TkyDuPx8r
ytoejdm3iWZbzoToaD44V5AlvUVxU7fjZWPEgzQLKrO0rzCQjHkX2b9dnkQVloxI
C2sARN5sdefygHePK9m2ALZWp1ysh14N5ZrO2/xUdVdnBl9BYdgDGmWqFjgeAWk9
HeImX+ObXrwcpxCbk0sDdI4V4l153ag1f7JUBr4rYN565i0YkIgpYV8E+T+9Ip6l
nvbDd5WcZ/q5fPokerdKNgCpOTc7fAp0wxIVsCYQXmt44lBp+hBPO0il1ef/Ut2b
tPw5r7YadujWfpnexYVxhxGoe960XasACWat+oaQWxrsWcBf1bH3BwRuxHZM75Wp
p/EcWiUqROGbQE8EYK7FimWdfKfxWoWTJ8kGvDjeT/g8cCD79Qrc0qkQt1jS3AhJ
0dqZLk+fjPH2bKNMbH6IfB+5rwlaAfDr4dyvXaq5X67OrvTjRFohmBdd+qKlUl2j
GUhdSpMUegeDGF6IKL9cux9lHbr5CwiuTEVJS24ukFn7r+ir9fdzExGfHAcs7yQm
Lr4EiGB9pssRAmmsSmXzcmsxeWd8EMdVxsyArJXEw0VSd9Rkr8Kxuo78BS2g2DdT
+OsbSvUUg2AlkKRhb2W+oNQtzCZxw9aUIYpf0ZrY3ZtDFiy0VvfvMvpsY2IS0xCY
kVNs/JtVGnFVjKuxMjhJccbfpgWQXNf3fe46e9YorDtl2HP+gub+0sm3xmrHa+DY
t2t1JNcy+qJdUaIX2waX1YnnB3ewY4i9BtMYQZpLDmA9Nn0vIsc3Q6AFIYnTYfOq
RPO/kSbI8eULQ0+0vA1Z/tbPMuqeWjF6OFmIUPhr25P+gwsi4Y08cm/ptOy++gdk
IQkkf7jIUj8qzOZLLnW/NHsaImNdXz9SZgPqgHV5SjGMZ5WHhuclIHVaZYXGZ8qc
nKg3V6z+SjpG2zOvAgz4KULof+aMx7kgKkZTxlouKjJVpjaNC+0V3Oq7gxd6Jary
IrHUsT/fxGLX2AzYcdwliPwW7LBrBAwPSTSHVY8dqKL3MT8tFld/VBTvwUgPahJy
s6vp5MdJ9Ae6E5s/pUy44rllPnKCzDS9R6E0U/x4hmqOZlXeVZU1lscyPmDlAwcR
wh9StnMmBqlgcJ6ZmV/FFCFoAxGKb78nbt9fXIUHZYHela5qKcj5dgLVmtfUWS8V
jBeiBxBCH9FRp8eiZunEdUGdWii47WBJ16gqN3v8/B6IociZDUpN9oxBW41jd0I0
hBsHzaeghviDssPGlGmRpsyXhG5i697Rymtzqb6GYgKnKV64nPLqQ37RCcs9QzYj
R5M9qOzLhc5Uvl/iN1y6K7vTb9lW6cpTw8ddvMykKFLrLHJu1hM9Ob5zqqK0RwEM
hzE8xqjlDqUvl6QZqAUq5MTjDezIYVrou+E5af9sffeQNB30mJ2hzwtrHbi+hLiv
Z63oclEBQWGal5DYbwb2j039JiwLKkep+lM6e986ZVi98NN0ufdF0nteGIXKgfx7
eN8GS2zaDiMvuRg0hQKwY2h0fnwViRhZYMwLpSSRUwUiGxSKR2L+tdT39LiToY/M
eIbTQT8D2MlWqkrN1D1SB4MIW2UN+y76IGv6oFWoncXQpcvGIBFSAeHkZtbjFHgm
HYQg6s5mqmra+cim6lpNRInYjCsSJaAH2EXY30O419ZojOcVsGTR+TvlyAV/C/dA
x9PWGB85XHt29YKE7c0ahI/5Gz99IDG3p+LT1SQWkGo04U5Eyzb7emvCEhdXapYD
uNhalyU/lonr3BqwDcd60bFLTG6hrcKKMmX8+jZ3Klf3Mh9ZsvNwul2qghsPUsMv
x5OjGGcISlYu5DJ2rbUIrtlkQHb8wI3mjQkje4TT/c7DVPDMO2x5BqUeZjeiGuBa
zNq4DhCYWDOSj5TCS+H38SyRtpEn1e4PGdndAMAMC71a1LaQozN4O5t4Dlew6pNN
sWndV0VlcaHH5vvM5JtcBb5Blb4Pvk8pL1Eod8j3ydB45xuIsjBLM6UaekyqBPoD
q8bnyfCqT6a4txEcrR6mLPBQbVb06d01vbzEuvZ7HqmQgUaVggg6DwckQXU5kLDW
c2Oyc7HbHi+KOkgVMEg1fjLlosWK56FtqbEqUaz3qh3JPSS6JJcVxgGmU3bO2+Lf
jMF60ZvXOOVtSoUqbdxdeyZLQ9d7kRVq+AJRb7G84Uz9cFmuEBbwsV9Ocp/HyNp5
lN7UqG7AnxKbwhocpv2tsEKdWKxii3tBGtSnSIZGzxm1Rq4QHh87OMR2eFYH3Nv2
XYBbXkELZ5960U3OUOww1ALyLX3N9r5WMff7T7BhGfU2xSvbvLYSUggjDWeXmiql
QkheyNQYYAGFuhlyYED6psvA/9eWe/1b11PYAJbW5Tp2Zgj+BFmWrNG4eTrsbtdd
8MQYnRaq2q0eFNUlj5MAWU1eQXiOXPSWngpDx0xmmVRxxmuz6WS79e7rWyP1HQgC
BLEGvddEEuctH0qfZTqlCq+XwX6Ck+CBvmL90suydEF/VEDtgSh6V9TZC3zD8eXK
EAMXNOelMo4wm49AwnWMPZohaXrdnxJuO+pPcakfPwqHysJpOUjRsF1wtgN/l+l8
eKCRkbN4OWFUDH835s1I3BkzCeb0fX+paYWS/sFH+w/3yjfVvQ/SyqXWPK8Emwkj
mot+22bBmQPepZ8/zTVGDhAG6dzT7UN1mIpC4ksZ5r1e9GlpKbSUdB8dC8gDy7iI
cgYsnafaZwFRH0XxyveGRi7LiMBTKps+y0QNN1yKXSptdfj+lU5SqOdIv+eyWB8M
sObTOCZhTfEkKGD9oGeBlSYdZi7kfUtspbIuzjT2D8G8WxFeRBSIs9iM921lQBvU
oG1OIFKya28kZzwVaK0N3tE6jVCTJ0hVwMM1R/gXpAc9VbCQfaYV/jSuuYLTdQCp
VX6BBpC0bRAdF1SQHMkfFIXemV8XrahesjHJ+OeSGPvwcAPesz6cQFDe5SZZKNrV
h563xmF/FFP2qAtaf99ZM0WGBeDHjc5ULZl6U6nFy9u4jzhC0gOpJBsWLDYNSR4R
+/5BUjt/LKZMaKMf7mpct49XkslFRhdBwF3tRUtKMg5Rsm1DIdRgR4b847L8Og67
WcOrY33F/y85a7/gogCv4KrXdEI1FW0Kq6Vjl4Yd7jBT+5dBajDhqzAgZn6Uw7vJ
5j3kKIVI1lwF9SvVfLk72rw8QSQgMtRzDVScYNbgV+HclcdxdyEqs1pyIpsaXQcE
QsZ8wsmi46PVaIcj2pKrJAImP1In2nO6F4B1kys+ZIWyTgQKzNiIt6FWG8sY33TA
aIaoeYpUgu23uQXq2AVBuq8JvNNKsD7IBJyr7O1bzNB0I9eA1P86XMl6pBUIBUWY
Aw2W2roqZY6iY9vvWrYwITXi+UR1yMpZVAFVtSSWSr+c1O8ocF4gAxC9ERsdIMOD
yrt/NhQLZFK/6nKWmGa3LZSVyzr6FW2EdFUKw7KL15zk+rMWclO/OTde3gEXR5IU
sx9a32fdr+3QdmEqnIl++dwtNfBnru7yOAh55V/VE+y2jAh8bQKYtpPpLsO05eWo
Wh65JCXFQklvQUER8LzlLgZLmChhpLHZfdB43VpIRlkQ9Fe13GNo5qbdk85JnEBO
mTuM9RAdwECwtViP1qk6494iYQ16oY5oj27i8lJWpfY0UzOer8r3ugz3p8rjr1Ek
Vx+vluD7c9aOM0v1oMr4AV3mzC+D89sIHsag+/djAvbuhdmtJWjtaRsv9u6WlVTd
LrTJ6lF9oPcMxVx7jNFrNVfoEugBirTznSD7SJOGtV5hyyOSuC7sbBtsGpI0Rtez
gOfD62DJWMRx84jv5tS287wAxoZIhEJaEtnzn8Y7Qj36aFolv5K7+B1+HmHhtGXt
JLfeWxR83MyQM4dF5ehAWk6AKydYkodJPQwHR/IakJkTAUGXUQ9Ix4sm4Uae7Sww
O/kp0K/NLb5vCM3Wq/9mERgXRtvWXBgS53Lh1SuY9P/qmNcPwgtQt/OLZMHyOKf6
jirfEwaOEfRBUFyaGvnQ2IpXiMGEM5zYKzGLAb8JEsHDm1wPjN8/jYjLWu4ZqMs/
yZv8J4yA+4fFYLP+iR2QiU02rF0IuzJ7RIZ6i8O3lRPiwiLAkv+HgPdN7+e/MF27
HAPDfaA4RkvRiC05s8RcGL4ssUQ/29vZU0D6xroCdEhyWlvpvMGhu8+VBreD/dm7
uZkuFS7AzX5VzHZ7PBLHDm5OFloW2mf2KNYqcxX+ROGCjM2F4bSN1dpu9EgplK31
1UsVL0EQtLV4LQQZWnatn00Vma2k2fF2BJGOKe5iPf2AHpsBNQj6ZHaJf6Bbv5hr
896TbYwTWzdyom+AtDp9fmatNpXxv9shp7lllpZOQNtJBIA2hxU+qA7F4eCxmJa2
Ig6dt8XV2Eq/MEaf3rX2mquWhY52uomumnVQjzBr3usHiSQOPXERTuwZHZ+1ssLG
atMXvcUfDhffwILfzpKYZ9Un5AraZhLz+HJE8/sfqmPgDKS3kyRyUu2aOPuol9+g
uA+ycnniHYWCx9uhxokll0JKjIWIGpj8TBQfW60h0VFsggLy8oTy5qpkx3tDSgWs
i9/dc3ohZ5NhuFDEU//CdX4c8rGUL9krqCvDYjgLQgQLxS6KHNItaw/Rkfgmsovb
pZLIy74e3NQHYgVy42vrhOY0vp5enzlJMDuXeKHhhCowoYrZ51I3QwRcAS/YHSAI
warmSSiJdGI9EdXVbOAi2ysdNeXyk/Pom54I3pU3wZcxuy15XxvIMhWysg27vUX7
cVcdcpXPOCq9IL3I/cML4uJsLQPwdk77ZEVOwbOJIMXgBbNEngM/tTXeTXd82GZ0
ciy96LUQKGT0aTgO/CA0cCzz2kzUEfpnKXcqxdTVPMx5f5GCe+GWzVacHIOuLn5D
RU5vRO8qHE0apAucUp9ddDfcsLbny3vCWFWIqwMckdYBJ4MxHfO1Cr1ZLnXSdo2s
6jEdjFhKF2b13BhRHS99JWdAXv6gsRPVIdxRnfHfrchBSCoI6a9Az8V4f0quDl2K
cD6bwUcQ2b6ZN6ajCktS8q4AYxcN4+eKQLByOp86NEnWhqgKB2z+PitwfMkMmzcK
JR3RIgVGl7wfhZ/JgJSK4MafkB3PGAXtwh3iyNDoZmd+AryPwHqmPcclsV2uBpEp
cj26d17/4HLXODERpzFWveenomKnqPb0w9w76KWZM2mCTA+sfEj7qWryTial+Dpy
83i1DJ0HqKpAX1dYGLDacSf1M8jkKjX9ptde3ye0kDg3xy9WmYyGoomjVLfwZAQw
t2ZFSrD/FOraYcneugSJfCIaYL+rw6vAhylwSg3OMt/uRF/ygAinhyjmjE5v+zqy
mZX8IlFF1gpn9dWJYeqeCoP8tFuubg/7v42RgGScyjPBzXGgj9F4HchBEXKAhBEJ
eKh0xDvVRTKkE0f8jJcGtBYmsVbrMJpGIBiOv/qm6qH5+5laWVXdlsmAXgO/Mn2B
0Id3tAmREL1E375gHfxOeBLqPmwcQygs4EuJh5spvb7xHfbISGjD/FzhRvu7EKqf
Pot/FZ3xEVibmNTSqqHyFK/LSPoIJESd7slghWykxrcq8VYd9vErlhN5VCEL5Y9v
o2oI/W6ZQhSK1yzL3RRdncfzeE+hyEsI+nsXkOX+ZZbcFm62w8VK+9lokWDy1V6E
SHC3b5wwWmuPbomsgajD/Fa5QQNFfL0NretKlKL1Xj6DLj01koVJdMtf/YBzXIgw
zqrNudmv3gW8ImTnRseRjR5RladWzWk22yXVlAJiIGNLGOmYpMmzlYOh/N5MzZeK
Z9ziHCwcaBp1oj7XnyImYqctZcqRKLts7CTvqqlEu4xFxLna2ZGeKpc0P+MFA27c
tTWgu7eeZOB8BQgCRyt8XtixKry2dGKudsfvn4uBAL1CAK/BBja7WDOc2rnuFFCB
Ff7cZJspG5vMrqHlCy/I6Id0ke1HrfWEmEIkZTl484AryddvlOTA5XLzrxJ5Rg2q
6MJ/bnQ8I2/q6+MSPPfKwQvc55OwDAeGONgqjwBUsU+m/Nr17bFtZf5Xzho0pTbA
Ak450hPPTpY6r1DfQMOJmR97UhVW1dxANAgE5yht1ZHuHkbCsS/BZncljCMn/BET
3snK8BWxMSnukqQu/vzfOxbY3ZfNxDOR8c0ygex4o2F9JNbFmV5sutb/JILzP2Go
lfU1FT7wC1ebtz6tu3poP44o+k+am2W/bWlVj50dQguRae2fQkL0fRAAr2UtTc2A
OEzNX6aDWIsW/YZU44cWMdJpyRcceWSD15DIv1LsHwP/4qvnQjbszU0U/5vWRjQa
HzNM/4xyTwd9VBMN8Mvp4Kaz0L9NnQNr0LpBPsG4xoBfyAQjT+5VTKxqBsjwVHB7
B5MaW62yWtPAdD3hEzYq3INN/lyL75y8VlxcY/wyJrz1rdd62BmLacIHcmMakTg9
3+gLf7dd+NiStU+FeVdTdPoP7FaUHkPIu47qEnVdAQMv/lV61REv+HcZ5Hqg0+Ru
hKchMZTR6oTNSI2rJKlH4mfrdyrDvbtBU1FG9Q3JvlOtsTxuPeSLqUga+NDYay2o
eoIhz3Pfv1UzFC9cJMF4QhwwkL2awAqn9ypWmtB9sD+qfK1Hde13Fqhql2vKF+Sk
b9dTGY8qtY3w033kCKH0BuKH0hHWXtGNKjpWGdcm7fMvOFQ62eNahEAytXvUjG4o
GTckTScLQHpn5o1i6Cj6aUqLEGPJ1dwfqDm1ymDoL9O9blU+iMO3KGaTWIIYbmT4
LO1TaIO+y+Pa/wNKt6Ed2GGgelxEhsj60Ew5RTBmew+Pv4i7epYsfdv1QIqOpVUL
uIbI2TjvovcjzdsiXtFHrRNYyOrcrcIj/wRfpUdKYqoleJvNvgjGzowqUMIg9rOU
V329ufPxRkTPSpUdkfqBrQOl8HBKXnFNT1XnoBd40DRE8EsXT4iPWDxBaPrIvDJ9
mWhm1NBDOnxdqJUDA5ECwLlyxJLFPKdlIzcuJTF9AdS51utHBfV/R7PmeKRmaFUK
N1AciC5sN1byXqVpv2tvFQS2EQGSRSHoSjzfz3M+Dy2LexpPag7uPnyaNfKuMsAw
chf3UMQoE1oD8wgEzrdSeHm9JYgCahIbxgzRd7qsD4Vn3BIozSfeGkKPVAqSQ8y1
jaygmkGfxXrDvHomzwO85fWYaPWtPndy+7aPFN2VUCkWVhoFLHXmBz6KAUSUqrJo
EwY9uJX6fqtczCWR5pupD9ymJ+592gKwcDS3Lqmwu2zbX2vAdaWA86bBWiBthV97
Z3rLyqg9zTExKAysRdz7XetceOgNlaT1yB5vz8+8yIgzwrZ1OBj7ZYi17RBuOJ9W
44r8OmKTUFZ80o5eTpxOxacbEXMdT/icpcFN2K2mzfqZ96dxZ7hb2qZg7ng3diCP
MRFd15ueQbR8S+k5IjBxNycuyix8+zBsbOE18I/0V9++CltIDQDn5RTVG7icZZhs
11imgzLQmqjNUp5nTYJDQggXUNEe92gRPMrM9xbDR/bjgc5HhVkZDRfzkDhJOZjy
JvXgqlQ8il0MA/225ctdMrAYQYSaBdAL8sHKWivnhBYedUONywaiwHdnK1sDtzql
679u89C0e8eHJCooJv9aaUu/8jwWWhbNJNRorgEN8/AzOIV5QV6CdSYDMSj2lvbh
wH/QZpcjPbvZaZE3vXTdrbcZ2alG8eouyu9i7DAFbeYjN/CHCOC+ENreb4+VnaaH
4HR06pXVQowVtEkBvF3mK3lD1lnD2J+BlMeYAi1CO6//6XJJUZ2ZxFohC6xVX6R0
K/Op+FNnSxTR0aiFNVIuep7aTseqg4H8cWys21LznRepclvIHSnpx6UjHVlBOt8f
hvIoC1oh4+0lS9z2s4Ak/e3IxsmtYAQ+tM6bTEc7JATVmvQIoxHRX77n3ZgOeuPX
XLdDKnODgasKwcPNBacqGfM0DqeEBVexrdcFNjALQIl2dnPnC75E1XaQ7GPOl/08
q1gp7X9Jyo8P+pQOuLY9Y/SU1jQGmG+1VfA2BMKAgACk9X0Rn6A2hMBYkFP445IX
J5uvI/hNC1Y9lsFn8MR2tP9v0aMRsgJxIqJmwvtvNFqEu0CgPWwjwyubS5CMKWp5
o4sw6+j5jtb7ijcsYJman549XxVUgLX+DvI3SyEyU4YN+QK2DJUha5fz6Rm+ejnu
dJNn6v9LpIv/6GLutttrB6nl9VqQxmiodaD1y+9doJsPBw4+9IC9ah5R4LOJ6kvK
1HkhyRcgIyhhrFIIZq2I3ndgAgoNZEPmyPrrBz6pluEfTleSMUiDDChLVlZoOAj5
LBkgSaxa8AegcvidSnksnHYPnpKFJfmvz0fX0q7bHgT19Mx1pvVlf53AYWhjLwUF
x6g8s0QuppLhU4m4HqHa4GWcYQJMjHCakEF4aZmaYNvvwJiKkoOcuYzS+C8hVslY
hoGEPRjsx9usOYgWXA0e7WgJYBxL81pPLiALicC+dYqNIKG9rueWci1LUaTO+w/K
cPHkcHvbw45LEVBr8io8WZVThyCaI8aEUHnBTEbEAceIRzI4ufGIzTM8fCXkLun5
m0p5F8aekaAuNx056gl1dexcTo0hR8gQCEnWlgiiJdBO7bDCSPsHeQS0VDtUzNqj
GaMkn7W7u9/5RGvigueIlnMwuQ8XoqWK3i7jbyDBxHZMl/09+iELezhYc+89+0Ab
gh1ElElYiSrYovIgDovQV3NOuMdjjDlDazmjqDlWHM6WI0MTcmSZefo/G8uaCEPZ
iYmGcyllFAhLIrm9h7qHut8gAGmAcNw8mQXfvcEUqWMYsVOOdI39taDnSnRqnu4a
a+n6qWcNEF8MMnT/CMmBNyUFB/qf0KQlUia1COt00Kaaov50J/ffydV5DuCmzeZb
9kWy7lgzf97UJXvRnCOCj7MZzsyECP2OFK5mKcMJ5HfrLx/QUbBddbxgFNDuhicp
tKTNtryIt6q3rm5nJ2HKjspCumnFbcJ2Wardh8cPTW+s5y3pOqhdyV685kNQt5Rl
ypz2tx4eN5135sT8V4DY2IrmWWfrRR38zau2Uu93lGuAcLu+E/vQeXC9yflG5Qnf
BRioO4sGZEckv3hzeJMZTex3GSjw6vVx1fGd5cI9kPFMDu2SmVTGQSKEAkErbrr+
j12TXK3oY1YGXZ3U6ZsUgnuquENcyzfOM5IS5/qBG+r6pLCJWqjMUy+eLGzKpPJB
OqHnHztA9B5oFftkriL/fGYzJ5qlYi7oigelPlsk5VpIzIeCrVmUCzQQIxOs4MNb
L6x2DfwwlxCKeRffwiAQlWvHexHtxqJlLn2I0aueHpQy5DrKIWX3lS71YCynLo40
fbVRcyjU+vvNhdfNatGp3P1vzRwM23UBEmFfdIfLIbdg5EMm5wzOGzL0cHNF5JIU
+dc7GkWFpUTlGBZLJZ4wi0+PlqlQ5zoqELKMMWw5q36ecXQGmWeEJc0f1aWJ+J63
SGjMffpn5sbmDZPWiZ9K7gmC5FSDDPqWqu7M2i6f+qriUGZaYOLXfKc2mG+PmuLm
G0+GGR4SakNhSbgnbLawa3VCWmMHOmh2b1FYcNmQaiUWOUe+8BQ1M4YX2AcmbJ80
ehGlOaHEYHi9z6uf1vKco09NJ05bRPnirRnJjbRYnKJsBYb4esrpaiy73hvj+G3L
8wmZAFx2C063vYwGNBeX9ftwF+Fz6FiAv1MIolS+ro2suS1F9pJ3RmvYIEn/4cIR
M7s+kiz7dcKN50pfUHnemdVEWZ+9RnSM6iUld2BGCHqmcr8//3TGHG1JimX7Rv3K
yoLkHI6k43EaILxs1trwUmPjNX2zm5ZorvH330YITteNJ37XVx7b1oXU4UUGEoui
bYjhDPXdjNXTRzGgbj9KxpV7SjDSoe3pBS8kYdGXRa+zTAynKhR4rbk/HSqMIVkU
onOA0VN5O7TCKP9ow2FphKWLdlwTE9mNRvDrZG83agIzkv7mEzwuLLquOT8TG+4L
VZ1+Q3BGdRK0Ps/UpA3uTXOL7ZNJ7wim426iHVqJKLmxRkauuphch4c33zQiId0c
449qcGbqGrLXIz06kdnIEoio7/QUshVqSLzoxXO9BhmUtrIjWSXG+NDaG5RYNBQ9
SWZCfcaqsM64tkQ9WlVdjh/7CXVEGBwTnQcBXTovuVZiDQx34hvpdHsiCe2PMUv8
H6oWKbY2qOvCQ8WiMTE57ZUG1BqcOTicaAmv9XZX6IBAsxGowMY2eo+cL1I6I2df
5nOkqOffubgrf4Aiz0+PxAblgU8l42/0jAh/GZ+zoNBQHTpXvOyUD76BKU45+Edw
MPZhYWCvWicVeUWL13C7EQ5LDA03gwyOgGBdjsop8T7uKQgUK7S65vAr/GBxGiLQ
X03W44kTsTanYH0wgLpjQy65skVAuJTb9l7X2yvUzQ7id5oCaVvAQ3ztUtGSTwNh
MGhHlwKbcAJ7VjB5neYvQ3I1YhRDlpsRzWRc7N1x6gBW4Teaoz8SHFPcT0VcIdPE
mmq25hhnW1Ns3m7ZTLF7HpUvwi0zmRDDIRmqICrJuv32XOrJWFfqdv45QtubNYky
tLuYzd8vBohXQoUh/YUaYlhBcKk0zK8+qm6/YqNB8CCPoN9WDS6jRFlCLkgVDBbq
Q6cnXSQ8Zqr9E8JZw3I+Vy3QvV2iqDs4qVwfQYh1/0mAFOD2pC0rCjPYsG4kPBD3
7UtOY8DyXEXlDYdlLp4TN0slBwtiCgUnMoapipxoGA4gmBax/AJRwKYi6lAq3pNG
4AuF6AeKLnXyzXXwdytTZMMZWRa14GaB/WywpXNjIXDFQR8FeXvOHrN704MSrx8T
TM/nqd0LdcydeUhNwUHqYyd3wPGSg7sfZXlTcMauLMvE9VMYp/Bbkk63FW05kbXR
6CenSaeARSqr/MjA8VlBS3c+/QHlehxkXb+nQclF++wxBkOgGMdjZ37zgFjdX6xs
qxqePgNLOW/QP6CELxvnH5+6QLxVlVQiBvjWeA4TCB1qzQI7+nLeDBdNsUt1AJnk
+xX/L+FEB/YmvS7VU9PnXvmCzYfcUINoDtOks6yzTVxZr5rGMqbFTj/RWbhWXK1M
1ci/+sohwdfRc5sbaln7NL4Kwenx4Q6e+St57iYWw00cGW4y/n18jG+TOw8cywCz
dXyjyxNVUlCt6QyDCl8otnM69vh0JaOW8/tzTZB21waQ91H6FM+VzRdQf7VC9WOO
blUirbShCb7Xfn+hSJgIU7WDjt1zq1C7YxosR2LAXQkYwisy6/NF3ZVszfD8Nbkf
TWm9q1Td/LGr2ejNdKAQliXVS+LDbElTCJgTM5HClP0A5JbePMYFXpBFNuw31PVL
9mcRWOzgb4JXTQM+uDQrFloB0VP5+/mRkLG9J9GCQ1nS17aqiHLMo4xz+fH9KCij
1ZRKrzleepbKS5EvwgoB8Ur186gvHFMjZhOXXg2r0Ki6PP5khg/le1BIVIrqkNYf
6IVgMSnwe4BqDxvcgDzyaL8ArIf3v+rdX4emTGiagAJQn7GU3cO37mrSZruX2oev
T8wtOKBEiQHmCSchZbkK8Vdp/0z54FWHocRXb+NoKFCBOVKDHICL4RruTZCH53ED
JAWEgXbkmCHUqqqNEZSAiJhFAWvYXDPezINUT1aag8hy57dLPiVfA9m0KxHvU81K
9NFhUkjj+OejSHFqqh4hvqvaDVlWbFD3wTQSFtIF9Th8m3vsrLEHQZGQrzHIffzs
kVJs9hFu3+0sbQSUW+Y49kgjNWqDj9QmdrJkYVnunNbyWMDX4g77mWXWorRVpvaO
oxl2GVhJ76jWDICSOu3WoR2yewYYlUO3iPjhTpILKGU/oIseMwOGx6yKsAl1inLF
fBM+dZ71sB7bhAtssPQYcKDXza8v99qvFEV+OBNb776655aQDPyX7VoADIlMKPxB
rHialwtvrsGSW74NtswV1fFAOMARVX/tixiCnV1AFPH/vKbrht6+9dZyR5BT8nlO
p6bIhgsNB2W9jqzugq+o+NRm+SwROnSsbNA/6Cl19P1D3T3uRJbRGEAnN4frhV9h
MceOSRVU/JB6rjSjR3bx6v0IVoA9ZPEJ2AkhrlRFQoSXzW0h6WkxKY0z2lY2Ucab
JPRmXbjld0gKKAXox3pv2m+gP2GWi4o/wIehg54eWH4s8EKQ9y8d1ADqLBio9DCl
1ymsjkNrNyHye1fvkwLgi4Ww0EIlW3yGLnEqhz+Qn/t6GJCw7Qy3QGiB/mtwoYsM
poWhd/08DLLmQM7Uw9DaBwAevMVGCBZ7SsuoLADgPXGaTQl+Q+6ForzdN2fhG7JN
Vmq/kmRBzqYIyd9uu8So528rW+an2LfjUie4OAOP3mN9tDAr1aAK+05xxllaJ8K1
lSlk0BhmyH7zEGwN8lRPSNTGvE7aZJhymstB3n7jQIA3+YnjcUqq8wjRgADzfXju
NN4QyTqtpmXuiX5WJjug2Ld4ypFYaUqSAwFl7F5YmxH7W+/h9l+ET73xlcwitiq5
/5visC2v0UavWCrTPsKGtcotClyV4TQ3y0IYgrgQffVIqhiR78syag4i4SE+yn5n
6HTVA2w9M1x6CzQKhQdDes9ITaAPjHSTy378g4xcC26JgECdBSvjf5HGd7v2HNq/
OA2j1MQm/ZYKC+rVwzZnC69YhZQf2bQeY2qg5X480c8zJisCPK2sk4i5FZGCpKTo
8VgvAEzFR/E1iXEVit5F6JEFx2s7936pOgi8+hkIPicif4pcM7XwKMQNw94eUyPW
PHYCnRu8ftsldsjehykCeos7OTQDP/8wxqiWFbLVXaTi3+jeYqwEQsjQGJhtj2U6
ChRwCYhB3fSadH0oRw7dVkAC8AIAUc4wMypU2zwzulV37YnvxhH75ZSUDDhfXaQM
wmls4jq9hPtvRTGCoQZqPUSbj8RAXDJUeidFurZPBXZcMHjB1qtC8+s62fZ/s4VF
Lf5UW5KT5nbZ5HFx08Mp3EUzouS4pRu2UScJuILoNY0TsIooUAlatjjYJwEsWQIP
zXCzGQ7RDEyScq55a8iykzrspb92I9MczyJ4KrZpPcAoVtdRQuRy1LIi6bhffGCI
kFaZQrgMtZh3pHIBJiP77QW35rUK8XZ0SmFopEN+XEqhVXr8O1so8Hu25ZKZe++7
EwY1plwF9ElIqJx1VYjX2m+TfFNl5U4+X325rPI0pcqZ/1YoJqLBCSKCuUKA+PjT
KsCKnKilaWjVrMnsXy516xLK7zce9omreMcYWhjisVJz7T3msU1rN7rXrpG0HRJT
ClCRT85QqnE6k7p0eXSRgxziHs8eqSaMiimb2svmnkoj5pOja5+hLuevNzxVA+m0
P/87T3G1YgR45jjY07tZ7c6p1dsSeNkWd7+Dl5oFTOfXFzoBlihI6LieDckCKCLk
4rjIwEu0CQ/z4sdTM8rH5wG/nhrwkv1vz3dUkdHJrktGTkw9Gbn0bION3r+fWanD
pnp3/AH5SW7hmZp0Yi/hI9jxawaKcozZmerUNAp4n8/cgMfKQwcG63WLcOvymr8r
f+EDCuFCx4vzlrKK3CTG2yXrmmYIn/OhvrEdb28KENe7X8lAfOU0Z8lkx7uDB4Fa
5mdf242rketVVvHDniYI2dvu/XMBfCg44bVNxZ4texJDTOIrP+m5znbkiELxqmyJ
jnUmL6dhDXJKtQGamtiETrjCom8+C4woj0VKLd3jMCU7YDYVFsyU5v/R/T6Igu77
p/GsFieSXDYjWc09wniaX3GgDSMnzoEEVhSUFTMw7yGHQLKzep5b2G/J1RPrvgcU
pOq7NbIPMINm47QiHKybAm1ha2jF7gB7bhDLIeaEuW/KXcXokP30UfKJ48fxutmV
JaWOwL7qDvqFBiW8r7tWWgJ6EURQfteON9SbXDSjEPafn3O1uCJLn7NIbIDkBdGI
DRKrsk885C7C39V8lVlMk42/gco/gAPbrb15L1RvG1WW/0oG9880YzrRyJnzNYHN
53lxL8FSrC108O1IRvuygCTxf+e9R57rrc+UPW4gyy44feTHj5GXwxaGnz4AM1Ue
AmI0ZZTvQRBTAbfnkyfmzbvqZvYdtAQR4/xWogfkQsC5e8Hds7wMZjS9DFgo5ePQ
szRQG5QpbPv1EVsurXOfC0doTCMPrqyLMDAAJ/YIXwxB1KwddkOx25nyYfWN/TH1
nM0+qZcZ46gNQPT2OX8hetJGJ53rm1lKTj2SkGM2JYk25WQ5BeyGOEZcWw7D8vxH
x6NXTeOJrzoyhmohom9+bzSFL8U/Lr2HM3VXgSwQ1JMX6kXnye6uzRrRmNm/zn6Y
ioMwcf2lFz+5xWJ4AvywXxTpvRxeZAFTRoNeLqyQ7Cmv4gX/wGEbKxDHMWIat11h
cDThIZ3RhPv+DOcNXuLMnIYhpfwdGMeKCYiEnGJr8xrmX2rd0CmwyjyID6mEPq+2
eTKB/tZDo3KBMtFDygBsSy0pt9xwNx7S+x0RNDY9DSpy0CHLOBGrX77bi0uAociL
X163sMjWxlYJW3Smbzzc35GBhnBG9Uh7UHFTT+huCebHMhw7avzM/e6p4gzghbk7
QKGD13Ucn+FFTZOglBj0lzEGQq9TNNEfnkHuuA3y+/lAH0QxJiPuq8C9QMl5HJ0i
aUYn5K3yCg+Lwa6A2nY7FXcgbAJgWoBNIYt2yC9zQV6V6dZ/RtMgUF7dkGlHU0TD
iOnLt7/OU4N2xLrvval+sjPNJvSmbFNVuW83ejgc2nPcYu8KE7hwFEJMep17yW8E
juTd90KdQ61pXcVt8VoRJTt0GxB56vNB6RhhsrhrSnHWer487Mcm3gXlzrusu1pt
Kv9Idc5FWJ+u8BosevvC+d3yH8kmXwnPjldPWE2gYfUKvfWalTqLUZU0ayroE8Yy
KbGKqX1Sn7KnL6FWlLxbamTwRGK+xzwYAwAqoI6qlP2UUiz3dC1x8ZkzcNesch14
Hf3Fb/BKaqdjHms5rL8vugbxofJ2WQatP94V4+yhAsOXPsjclxlCsA2GA9MWl+No
EKZpF0KJirN1PyfEQYcvBXoQd2i+qDIqN6db2CpXbmuohGezoTNOkHFJtvhGkXMj
5NJTParDsKjc5tS+pqCXk/lSIRlD6gD2H39Qyuy0WMVFwOFbELopIi3HFyqIvx6i
dlfvjiArZeywp1m8Si5K5BAYtwHgXO8mBifIkfi57Xwu+d1ImL1rFvLAEKSEnU8X
DRMndbn6OYEY13Rs5S015TijZL7ms3ODKqmYVn7eV7wciZIbIWcYQZUTPhNnOGnp
zkGAWRlVtBR1UYf3ecrQdtzKuOAUC6QByVAMPUOcSaoQCRpggHBf2btwv69wGic/
/e5/ukn0053tYizo/LLWd+AcOIjBMr79eaVmxFCA9jBSTc9LxiI3WvbAeW8MXzzO
0PwDEv2vEiCKA+1BWyUV2u5NBYE6+oehvbeB3laHIAtXn6z6/v3o19jzZcViLtSL
Jr40PFSke+fdzsIaNGjuUMvjtfbsHfPrU71fx8DCgAIHEF7X+u5blG00eN+cGy5O
8RE+4tdfgtNV5Fe4/Fpmfbvevawa+/ihIfLwt+WDUIpBDKp3IcCeM/Z4PqWk2AEB
y485Ay1l4XpoCFwHP9dSjT/2CCO4BCBg9VN28Yhs0ek56o1rJe+yg72j6xCePGHg
VbMr+mLBm+gUT9BTcneVE11UFlWAsGGlUUNr0f+qbPurIoqzPc20iXWsgD9CIwDw
ZX+Szbd2NCDIGy414TNVvHy3awCtPvix9dJ7ZGAzrav5DSDSFvvytVuM/WUK7z/M
ybEWN+iD/6o5qiwIZrWIMIjUhITLCwUX0HDU1+SHGIAYvSaWfqk5nfTGhGWE9jKf
cNQuQJEIMi/M7WKQIS2JcOUMeJU+wHjq6L3rXzvgLIKKsNLLEnYXazb6s+PW9XrW
OJ0YFQO71tztdG4wye47n9un3BQliR9BmAPEtcJjmSRXzdmKOmkHWcRrSEep8rG0
M71KzljupcSjvSe4DwRbXweaQfBaFBTm5a2KB2fI11R5XVangIkwrzG1aEnoeTJM
iILXhe6rLhEn3m1J+cw+0g+aP9EHgQRImcvLMJeIfBLsFvEUxWeFPnDOB30ziqbt
ds3/me4Z07bpm94tInqmvUVymcB3VZ1TgIVCe2hxVWo5ZeJfs4oQh8qaaJ1iNmc9
djUmOBQycL3gLlXZrOxca9ecvBH5szrBAV4fm5VXJLUT9jDqttMv+tyzLj3AayPN
UNJbaepGB6uApDbwNJDXebxL6PBAPkuwX3J1MS/MTFoPL3osAnflIN40tROGeEtm
JP2GcKPHNS0dMJGxsd+iU3r43u5I2BaeSNFFLfgfvU1LTbTVWD/l/KzGd+NUL1Jz
2lhpBZ9za6tWqR/22n+LkXXsZLEwlADqSVfTRCkGucnMzKR18lPU9NLfK7b75G5I
y3ssYrfpbLkpJmThytd4mMd8BYcKnmONsgnWiUucTmGdND682eAbPK3kLmQW8Q3S
+ADId2iHcQAfisUaiagkF5IxQ3Jr/o6kPzTO+r0NyqGm8x1f55oXUME89nHlsyMd
NmNysawNUc8ymnQXy0YeNRHw43ornQuhX1H0MuXVY+4alox4CDm19tgqz4IDKswD
JPT1m5XXQK83Ca1dZPzZwo6ol9Zu+a2WYId5E/5MhwJZIiHi06x6HpDgI3nxshYh
5irb3GzJOFRy16HI7rbP1KTqORwiquMJD4sflN9QiDexxGfhjzRhOjc1v2XFkCI7
EqifG6C/lU8YJHhAcuchdTMYsA0kE7AqILBea9AQFqBUGXOoZqFZDwK5w0ZbPt+W
ljPc07/NlWG1CJQAyrrmuUF3gFTMexmfBqdFaHkfwyn8QHwkg6Ym45fEyPTOzBFq
b7Bs4Soq6lAUmSxHCft+C5Goq2TJ+O2Bv8G1TyjZR7FksXcZTc1mpbCMryOVAY42
beUSOPd8y4GK+6ZlHRweFFWxW5CvIufPk3tloG+YjXpUfwon2Q+mOK3UbondWQbQ
DxIqG3NjsBBRXQ1B3J+5YAbQjwoCx4PaL8oHjLm6eO5jhSuyP6/JC5fXlD7XK+at
lsXNDig6w3Kixa0cI7eDNfNq5/d+/bZlpiieRcTwjigxm8UrHtvYtnShxLQR/JSB
0oMJzZghquT+9ekVOC9BZK3aua6V91FAL9pLsdjSHXu7/vrE1y0kaq6OQmSIS2Rx
7zTa5ok5ORstDtl+pobL2q5bZKegIs7ae/ILMJsMe6HuYIaBbzMkomNPM+naDme8
8Bzo2Ozs+LXrEQQg4CyHQXspgvBfW2zOZ6XZTjRrxnZlRx4yg4VOraNKYoINn0VV
IRnaVAR5Qf6YfaqwWMzmS8DAZcOV0EWT3dcQ+IWNCFwXDDvPcz+9bvmiS+JxdyQq
CgWWjL2xJ24rq1pBKUz9U7xifFGw7Xt74CXg6Ub2YlyIpbHEBA8Ynneovq3sSIGh
np7Z8BDuoo6JsRwVsjSfD8aITRF4EiPiHCww4Yuq0NyhP9CaEPStu9Pm3/jQnV46
6oiuV+zwt3nue9p80Jb19eTc8izMm0Q40l9Ji0/0lujVXS32dBdYKtXu8aUE54HT
GckE05C5e47ND/m+VS0AJ3CHgeKahv4p8B/SAo23ol6Oe/SrpB9oXmsYA+a3swAY
XmASrRMVeYY0Y+lRhXkd/KTJU7chrvsSWEW31ZLwckZ5tZu3NcIQn6OWGpHZd8lK
ZRXvggV87VwuimmcYEodJqC2H6Fm4/IMbfJhgeKdJVOWNz+AFZGD252IpjyOcN7W
BRsPNqY0756yG8jHE4E2SpaqnFivNfBfp6DIsFpfjlD87trva0Z7gD9iKOzveaNt
dnAZvwSvaN8OuPj2/ne/kSXIdGV9itNfuq12sI7+VWJH7FPwK4SYfThA3HMIcVZU
nqr2lIRThV7AsPlbAG8e8oJuo88bVX71JQHGQmd50/GX6G8GU8PCJVAdtMd39MpX
mTXOJ1mwQsQODKw5bhHagbnD9QPR6hsREsmRHPyN8icgi2gUaVxR2ocHHj5ro1sk
v0FRV7N/4x1kDzFIaEa2Bnb3xheXgoNw+f2y0hNXg1MMZ+8K/yfVcAKJlUOrPwJa
5Ixha7qX1hSN5z6HlwpjEXWbIBzA+dX5RjrIyDX2yDuCtHn6lYuX0znFSWlDAIGi
x4wS9+2erU0rJLNHJlCS/E8j23FSHpXJ9/BuZMsFZY+EBmRE4lycRRCxpApV4nty
IuCYDFRwgzHF0oy4gWdy9VSVlbiuLILT5UMtIeNi+wxI89gnRmS8a9fM2B1P3wUe
ytXa7jKhonzJnkGhN3tjJkqMjQlfxsFcQ7YqiB20zGMFLbARQc4Kd+v63xO9yLit
5uzsBRrjFRAOeuvJah89qkmeEG9Plmv+E9f0EaJd09kXjWE7JFrph09d/yiY9szT
S2Jt7AkhKkUUn7ZikhXJ7DpcBPxfCZoUTISyet5M7agnmlIClrM6oYbDKFj2F4sH
LLFyGjDW05nUYWrM8EipIsQ7CNvo1SOr0r1CdRuAxw6yK8Kd7qqdSCrH85rN7Wis
V5NIc+tHcXd4rIGAmI9ryZK4x3/H9CT0s0Zr+8ujMLXICuwXqRZrBf+HQ4wJ392T
vhtMXVwNc9SqM9xrNN0uAU2WVlmQq++mhlOdopzsJksOHE/XbGe7rTR1NGDuWkeX
EV36WZ4jz6eRxKsIgS2k+c+P/sY4lZpPpbKOXLMngbz5iYtXVkmz1dL9svP66dmR
81xsKYffvM3dZ/Kzfy2h4hxXlX/1JTIw1mhN4zxch3V1dG/Dh1LvLvRXQtj2pnE/
ibFYcVogo2MppxBVfJAnRg==
`pragma protect end_protected
