// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:40:21 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LKWjoldiLNrheZUBbiPUY0WCifbr7z2gEpgyW7dw9LiZi467rPy8fZEIcu40HYk+
HTuGRV3a4AGGliB3Rc/lqsLKCKn+9M94UrlUudW2yWOwg1FX8Q0a+miEt1HB/FQk
a4E2JcGhoT5kklNZhvZsHr7kj+E9ymQm74oSDrljHyM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5792)
AOm5JgVysFdvARBTLi5HjiUcTtcigEqabFUtjCMtoEGEopcVYhpLkeMJVP/7uQsw
979RvDjCNsWmjJHl4Tjo6YfNVpiWtc0swX6aOKrNttpP240O+c1yp41MuWZ/xAy1
VH256/x6tg2EQWyL4j3Hzt7T/j0S1vcWryLkMue67M3WdbLocGIDY5UA8XiHPOkh
ccmWPnue9BpSSwdzC4PsRCaKZJQvunaB4LpHrCiO+MiRLXtNc3A2S2Mn8DCqxsxZ
Sasf/JOllwUUFiZ+Qzd+qlmAGDDPYP80g/vX2jgT/LLuE3zMhXKxN4OEbDhxC577
7AsQE1nHr9l7/gSzmE7FgIJ4PDOvoOagqkAOetYsBa7ScPOXHap3kg6sEo5V721t
eOe2tzuv3K11NSl59kpYvRnS3Y3UbZIfqvqD0cwsN74t/rXeXTuOu1pFS6R2uEEV
JazCoCJbeqfkKt9qGMlCWqzMGHgro9usM+PhIU88Hx6t+dF8YhAgcfDN6cBxy88x
Fi7gCBRX2HNk5VSN86agQ1oORv1m3p1qDtB1OrAQn/CYg9KqLAb1eL4WkrT/2U7t
5AWo8DmOQUGRcxyvQF6jW+0Nsdxz3Sgu5oGlMbmlPnJkfm1Fje/dMtJdTUr+7Vp/
FDHUyHg18iD171A6iRT4HU886borTSd0h0J6x+C3FLQFBWFeYDD0gdVeD8xi0SM1
B5fR9lbARQnqulB7X1GeNq+c6aHAjaHUuG/jKyrfPZJ6+km8IOh44TyrEsElkQnQ
Q4ynhrDr4cq30RcrcJ+tGlzGW+h4oWLh94hnqXGPLtxOYtmWv4BP+/aU65+UiZC7
KEkVtKlrZNAi6sct48RZEm2cih67yEKZ8l5fuBY3zlGwZjsvzro5bWQOljm5pg/F
znoYufMAzf1T1rMFb2B1ti5o2WW3PM3u49h4R+yDgMbnR6wVM5YIXq4eWM+fStaF
IMMqE2kOrz4FT7hpSj/BPipZl/Hk/sOUTdJearkOpQfacul98IWzmbA74tXY/ALj
7Uy1XXrHapmRfZloZ0aIS7QCr1JZxCmrQAHYVnJm4BJQKwYhoSrYBbejZr1/gCfe
C6KQUFjiCp5sGDjzrHNlaGvXiYE42HxPLlHxqUM9zF4aLpWhBEOUeQazCmnczEjN
zaMcRI+coluylgBpqdn97l1PCu8rc+gjTCEZHLfjLJuBagaDwp19E9JxUKw3tZmM
q3jRw36UJpYLh3OZwAiD19Ze0RMe+GoyV9MUw4IGSh1Hrb28lSAl3DrrEeHjMHoq
0qqM5nadrle0fGmAtFeYKAL0ATY+IuG9XkgF83kjz9QsaMxwFyNgk6IjV2TlPaCA
gbLe8HBx8VQME9IbOYrsLJb06tCZEiQ+rDj1L44GSs0fkS6rE0JuFQI+Ifvqvsqa
0tuJIkCGMdqECMbZrr9qqr+3W39ZtFjimxisf1nUYIOS2Fvf1MFeE9VkheaedsuB
Po7MtxLzUq6HLKdNnhJakL7Nwt5I5n5sWDTXjPq4dRRzEmQlSoNff8+bIF9z1RKI
sX1j3yLhvc85bFky2kY1AV8gi27C//ozkudxPsgrMnl0eaumMlojn1JMqGPUy3W6
uy5TnpunhX3zgiife+DNud4xgIPGmjuF8ENdKTGKGK4H6Bhwv08x9UlAlOGv+oke
KTaotG2swRj/Uo8NZePdFX3oNPSgkEodjzzocn1IceAYj7dv4Ko1NPGiyOU4Ua5D
LOxHDzq0Qgl3KGC4n5ac2PxvJlf/kR8d6tjZuY5T3FimuyclW+prmDdqN4BSWjgv
LM5R/uwMDHkp6jIBv0do26VRBqIlVhcuS9BsKtfUCGHThU2XZDSeMY3ZDgZKx4y5
Cn9tmvXo8bI2ZaNE5/1uecHPwdL1qtCiWlLcxDVPlMCR0oJWnrmNglP0+rOkNfft
DwLWnAnigHaoEWD8zGQ3IngenW1DwKWEPxLKMnbqbF7SMIGLqYOmaCsB/08aejAA
1/QrYcR49saUf5BaHZ3atHdfD7im5uOKojMpgXJOLiNfMd17aIct+F9eMC/xL/Z7
HWXYSG343WLWBVGAQmMlXptyyBocORLGMA6+jZfdpcb9RHkwpdqbErtj53GdoH7v
7xvLzGB5MLnhK4vm40AryDwlngUghQeUSD+kshW+mdJ2bSPIj1O89UquCiZJ64X/
Ukaezq/gjbOgohVl4WUUEDgM4b2EhfkHYwUla2wcdH9m2PSHhKMshKqwhBNjw3kx
YP4NX6q5MJgTVkWsOpJOe1/EhXPqaJ5N+JrO7N4bR7ttjwY6ddd/iAw2g4aeMBHa
ZSRBAn1Jo7rv1FTeS5KJyFxOunS1sz0gIKwcvxY6C8nL8Q15D71CONsrE53uFQDU
xWz+9REVKjlZl3R8VLck/rojM3LXVU5BGpCX266OAY+H2hZl3650mFqFJwZhekFk
u/MZzPhC22LV7l0ss5CV7WuRzpv8Vk5bLT6Blu9ZMfadNRCdF8zestjVDlTrOIU2
QqYl+qf4mlAsdHRwfK5i5v0e4u5LFQ/AFvaEoOB++vUOsahzzOYu1I6jmx2mX+T9
TxDxPhhBva+ciYrkZyOigENMqJR1OVH0/+0MMW43R2JsutA68tNZvqINb35bq6sp
vhgnsiYuPdz+uin9DKRsEHQpWobDok1CMvNWXtyVrpUrNHYjqLM+FMVbFXzQ/+0b
p6Wj/Sy1UVlWpV8CIuKPk2nArp7O4lt9Rpn/ql8nkjN/idrvtbuU+iiM3SWRSbZf
pYLtXnRTwdX/JLvImJlP7FMgv7EhqxfAtJY2H97eypD4Toi5ibHFQ0X2HQgN0HII
KJN3ZkrdNS0foTGlfqY6oTs9jgbW+0BmrzKKkd3iMzp9N1uibkz4COzI1bKA83Zj
/hPltP0l9gAMibHTRc0zjQL/SVzJhhGf+CyfIHHwXqsACCIMwT71EbqUI4Xgek8f
mFbhJQUw0FCmKN11dumQiyyn1MFu9nppSFXkqd7cs/IZ3PvPgJuDV7/Y0b6TOcK6
Mld/K0Xr0631cmNlGruLypw9AQpWmJRC+QSMyTWN5REVinBx1l0tDycCUkFhOn0g
cWFihR848OuItQd5xWRDowhbPsWMaNQSohkOCAtprRl5WZeO4AazMHy754pS+uac
7X99z+ALbDbhhfClkLeFnzak/9mzaO0Ec0gX3DIfi2/GcjIHqsdImE3kJK9PJEVE
0phEvvHZvjV9meo3BBe6GJGGFCvBHYVp+0Jkx6oHKJwudFQn8VhY2mILH5afbhSO
FGAdTNYkvnmt+iu2gD34wAFXsiCR+oWqOaw56ab4Vib7FrbVFZ1cikQ5LD6hPQlg
YSM+I/c2tf860RRlaj+8zMlDGypRHChboXYrymy/5x62Hj93OFUbx90COOltiZRS
34yarUzA99lM+BmoqJGfpmTgaGFQJRELxoJASOIIQ/gqm727lCk2YsLiub/I1HjT
fSuTnYbxErv5sxmTnuyMQzu/s4KeGsVTaCocfS/0mWTE/7LDUogZs2mBt+wMwIXf
RnakdrHVxbLdqH1vzDYrS/M0fRxA3oz4Ht79+ogk4KSXYZQrKjxrg3C2S2rShIGf
+8h4U9i83Mp42EVaD7U+FH1vcGULJXi+rQaqb99mLrqrF1zq/wfhvL0qZvtTYzxG
DU8Z2lTxXEC4EurvxNXq0O4jHApipO3PfGFREYt2pPyTdeRjSROl8y0xzflcMJnU
iF/6+Kar+24jBiu08j7cMaty86kcb7yv61onRvRk7GRZ4akxWodZQNWVSdPpN4bF
8pjFmbn7TGPOb/UhffUhXHDVPzEm6bAUaHOo2yxxTbj8gaNJmCr2GK3aoqIFMiGx
Fixop3JFok3fUhOI7Bi0WePb/dae30HlMuFONzV/WskHvEmRsvzoH1o24OE3LsiD
yRUXLB8wOXzsJj7BbSfYJjNupZwhsOq9v1Q/3yznpHaaxBYrUSQ/1+sCaPWbx/RB
T7FC5RjKX6aWxCpJTqhaZ3Ef5J0LmsRSr/fMS6p77E6001TEtt1+vmuAgwxC40DK
jfZcyQBvkIgLWKIfSsbMbKhOmB3bYXFC4kHRdqGC//wRRCcYrVNOGlvQnHyqpmTz
jZ4/4OQ3fzzGq/pYcw48/AxIsQI+7+eIlg2Qf/rINJJLxEb+k6zXdyTfoYp73clR
fB5FUqvV0jVKQiiKrooDkhNxOQNyDMq6I5ytDdgUfmoHkE2ZeiVTNEOsx7ulwDhp
rUHhL++IEuMh+9oi6GxWL3pepiojWP1p4PHRgTtCqvFeFFToSgWPAY5v3WrQAVSa
dPxJqAUBktsQXU0ParJVRsGvMds7bZLYGDWSjUwC8YFDcGiSfcQhJNJitzw5HcQb
O9EP3uHMZpPz9JSufqlWOro6tZO9JqaOAXh46J445rjVvihhPl8TFT8HnxOew1BP
DpSPSgPSvpSx7WPuwcFFUdOVoAtMzTyKN1AOh5VoZdUBMXNEPbn5gtny5AVmR5I8
yZ58rBUOZ2+4swTyDSuK9Dbj88K/Ud0xdtn6v2TnF08XuxqVWItYBvAjArMFOXvJ
Job32h1q7UB1v9DUCVSFAQmacLKNXGlCal37+jv+z0JCW0nem5M/zlEfKDn5Ky90
5C5fgZn/Asj3hTeozk//nx8kJDIiL+WeQ4TB1l4ArE2GN8CfwO6F/wi1KWHum2jt
rkATcXTTk71e172UM+wEW6I/MQw8HCpn3+DJ85Y05zGE/sL6GQ/tt2oVbuC2cJSt
/G1si/igq9jcz1jyDuDuN4v7RuiSRSkPIXBo5/RHk93B22NzdyYLCOtdAcrdAiaa
HUzXD08depFc+A8CeKsuFTK5PZh3ClR1mK98L8UsjyMpiYYAXQ4foPmrer6yboFE
HuShaVyy71NXYcZU1oL3XifkglfIbHVyBv8qk0A4Olx4qWRSK8tTPW9CwsRTs2hs
+CAvnS4umPIFvARdGxIluN7nXJexI/H/1ekEKUFbYQUfZVuNeykrTCWH8KeTtYsk
RbMqKA9136kNCSicnq+XlAaKAvLbkplkCtpK9BbJCgb32XpljRUfU2LfFebCpY1N
NXn8VL6KkruWRJaKntnf1fJla9A6R7UP3UKnwA636yQejwBjCCmkYFf3qIAwqu6i
YS7gJt+xLtfqtZ/c9WHzFn22hjXkxqg+cOGGc3tP/31tVUQFqY7wDhD/1exZi5hR
QkRCRlFnbfj5bGe2WhdgjDHxR0IFF/tLXwQprUHShu53nlBxAG1DXZPRdgO5u53u
ft36HyroGP6uDLRKOrJhHS5S2HlPabgZ6OX/UoND3lw1Ps8eNry8kzZt6cWBVMto
2Y7VSZl5KLKRJMP1Vdb1ilOZdYPjVrsPP/c3YWqhaNzJFiOfeyU39rtknpnA6G+3
6jkAJ7O/kQiyS2aigAK+vqkDrF/caNjE//918SKU2bKHhC+qjhWwGhs9xByKTyYm
DCMeN2UYGGkyRiY5IR0ZJ9amofW6CXaKM14SOaNTeYbzRH9tR1frKVWFrA7Xl/IW
/UkupUcEbKfW8Mm6Uw96idPZPKGWIqOW4DNVnMbQsxs0cc3neTUYiFVSwmob6bEg
Wb/NdASnoNQ9IwxnjH6kDpxhO5izdK0x6JNOarkw4tQzAmBWZANilzfl052awB7i
6Us+tAhLcSMFRedVSHR3EEBBQOH1BR9cji6nk3x2auxM8iORKb/Huh/lduGeJVrP
ctZRJQTgOZ46Vjdh8++4N8HGlnRdUd2XuCyuAEX8rTtpYt0eCKZhG4iL5vErniLY
ATWdESyDvkbKOUeLqZHsBWN644mHsACI7hA/jBFOartis8/EKcBwc+YH6DEisyDi
cHP6oT78fB8R1Koap7Es6iJ2c1v5zMpaTCjOeqm4i8tONUr/swHmi3RrgO0jv7Nr
nHhxHaRlmAT/pRk8RusFQC3CXEbns0L2N0ZpLdlzsaDFGV/pp64CU6TXvGx/C00+
2CEg7lZPF3+yXCLkl0dXNg7QyrO0Dz6u+HAbF0tz5LmvUlSlgQPYQJOpad3mUCmQ
dBkSQMYVVfyRh6ihPhrONGe85EVVp17TRkJt75kAf8x8rtCaxLoRBE6fqpsu0hI3
H9caZ0ZwlhEsTvgsqfw/9jJ6AWehHABiqggfxPskXueGGCXF6Kpp4n7WhPHCrykM
etcNHWEOtJ5QKmPm7+DLb9H8b8ZcU7pid76ZW/5lacUrP72v+PO/ByOxEbnAInnK
8RBEbGSUEqc0P9FxjxNOw1G+zWINr9nGKyChcKlzr/t7+9Z+266McKj8U95lNxr5
r3YQj+fcVW7aFZX+jI6nEmJGj/maOdDQRaoYo6e8mePV+/dTV5LduMxvpTM3Rbnc
kKNz21m/sf4uxYMYTNzIHTmChNxXtoGeL20D+5TU1odBs+s2UvzeWeUVCgn3fHUF
RZSWtRw1z381s9UdEFL21qNDDe+RWRpskgMI1DLc/WNaNjzsC1tTiIXJ4XCcBwZl
AA67MMir8jjtIqtnfe2j+HtaIgeijmvIDfNAEvvoG+V/Yg9crACMFc6WacNwx/+6
ji/FSVq9RPJH0oeo9GgH6+BOPybRQBE+vooVZyD04lGiutNY7e0sNZ8NjL4XCZQY
N0Rszr+RrxrTsuHmGwuClYmuFvnolOEDq8Gd5S+E97Jx67qyaUxkDEVwg831/1rI
tjrKyvv0yQpVeJI8vm1NKMvjNh55lc3sB1xcshoYLZwnTxZWpDRAoj+lfLB5M5qP
IS0AFvQwFGStn9ehObmY9G62yaPrRHgU6jAgByIFiXkiTSS4KV2EyMNAPJELszEr
yhw7hC4KAUJDuqhCiZbbdKQxUDOGP/GWcflGU85St7xZOWt5QoqDWhNKab3ACJgx
8Vg2jROk3aBugU33PsjrFYeMvAbO0N+snaP85cpbTjuNboRpY/kZ+d8Lm5E9DxXJ
tpesl1Z9GZlW4jAYdG2kcwHvLOl8xmR0tp/pn/tbxuSLpy34tnRNYamgrn8fgUlo
L48i6r1omAwmljfLwQDNNgk7IA076lW2o5+LIjrXdLOijioaCaLAfSxs4ZqodjC+
JF7Ouy2JH6xUiVC9AoV6vxyjKB5DFBUJSRDoPQLmCAGBG9juyRkjxJ/zhYsBQ654
VNJHm1DDrM7iP06NEUxEf6sqQOmRi1U5U5BDKaBUd563ho6xJG22SrFujTfZNwED
9JvMmeMsdNSmFwF6JM42QArXexAvd//HhLUhjIJDAGktA9S2sGIXDNVC8MDlQRgB
h3SN4TiizU+hapLeTl0KdlOGGmYGd0V9kBQiZejZQperpRvv0RxZoR7HQvDuoMVO
1JsOVhZAwLHFmUsgX3QWfcYHSSJghN9Q4m5jfPlSZNUXJZPMiG0rEFi/BfTUd5V1
mxLY/RxjHngTrOUKr5/iRYnNHSVtZ+9otkCzD83S1EyN8j4Ay8UwH6/8cIIfKcKH
jS2N53+vXll62Vn1MBoxcX1n/rrinq8lPo9G8DCJ/HPf0W1RHDEHFb92TeA81REF
kxUXSI1nUG7IGAgfD/TuUNbcsoMxNP2FiS/gW2TZghWBCO0onBClBWd6Xz9JDhTo
uzA3A/ePz6DCeyctobE8twNKSXlFZn5L/epxgEbBYDZfm+FwcFXtE23hcpEK0Uj0
17SguYvK4o9PmZD7XlzqvJqAMn87dPQdXjKGu8K7aWMkwPGThRMrUHH1BvmrUd1h
88IgyWl1QC2rNoQ52TfZ9xOjnmB/laurNwZBqnUYpps=
`pragma protect end_protected
