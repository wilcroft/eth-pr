// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:12 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BFsK98LqDd8elwSazBeYWboUXVmb1KpAjGxpkwe7PRYIjl+UNbNnPzZEQNZoyWAe
33XV/V1RloeZoUEN9vTibmuefe/JW3HOPdFDNJ0GJcfxiLV2QTo49yYxFtDbrsS0
9wVw0voMXPIvddA1nAr52xGk/fJGnAe2y1rBZg5Jc0s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2288)
jNTlFmXkdK/L9LwpaRu74CQUbXzua1lUPcss3SrS/odQDZfjjLyiwongRTPWH7gD
XibFeNDcCA7x+P7axw9zSgvpgiqBitFq9YHXFRq7YGhrq36ueXqvnjg2WrPMznE6
4SD0xpCln0K6q9Q2c1P4lPXO4EQyCtzThbZXCoODRR0r2wpj+m9dS0Vm2aZyHipR
8IqNn12KCiTMmRZ1Yv/PODK+CulekIaCx5dmdszkm+0XTUV4HZl7E1xE5flv3xpw
fjzgM6jIxHFKj091MStFkz172IbwgdP27eBiVRd9tNMu/3y/9HeLt0C5V1Q7QiZw
qWRFzpzz5jxqWo0PEChY82WfsC/VGF4OGOG7wf3FhSK5Jv8HJKjbqn01yiQQ6oEh
SoDJzUp5qenfBI7GpN/z6C9e0L4Yq0PRYZKAgwW1Da9l6oQd8kkYOKquuErlHXu1
DpNJnD/aKFhgS/eHaXvB9iPyuE/R0Fhd9tlJiiae0jDjDcjYTf9jkiT1MX1mZGvt
ct+rIs9IdOjFXmQ/Pu8AjO2bQUnEciRHNk/yGGWXOyVVLK1+8kSRfQeyxx/hB/HP
06z+qkKVlvRsbfPELkAtG5bRJFhtzHnkfoJk0c3jvTGLQleOWihSuuRdfVSspBAK
vUuxgAS97PwJNGhkOn9d9mM+9nujIgK0EcOIMiPeW360bKPpHsU+yzv051IolwPi
/3qyjuTqXBZBxfpmj3cgcokfaMdVEQ0q4k2Fm1CFHbZdq5lrvrKbVafUwzV1OUS2
N/Xnqwz4U0Iz8Zv4d2/+RKmCCcKfZaW6lH1vAbIHoKRO5KuCWhnCZjrr6oAqeWCm
7xHQwYg/GuNqezgp23vPEM5KIVsDCL0SHZi94/AqO8BNHHP6owjJPQOGN9N4/O+Q
00Jk2S+XPJ4LrHZb58bIZ6HjL0P/9V+H8N9g9W2Bqi+l+oliBQwujRf4oXFAVxBx
7/a9pFd67eETBtOqiuT3BS3wlVTqgs2t8OVLagkZymmFBER23Qb392IhRWL2+cUe
a6Gjtc5njRi1Vj3GmagP2Er97Kxwl64fyE6IrUUICP0B8cRJI8j6WRI5ddurQnFJ
n2cHdkG0xFL25+bvRtuhtPVuQmzee/1lQ+KvD8DfuKHKi9Cz4ybJCBLP+RINrMAd
4ihmDhGrZgs0mcdEjBD1AmHPL397sx+tKO2cv1Qm+xI6ddxXDi0K09+lIyJWtyDD
+IB/xsjGmCCQpViiJIp6x64BhiiOCG45MmevSaApj7D2X74yZADy4TRpFOiYQVhf
JvnOK7SlQjCqR6OxsWnOM3AxyO22YCnZhNsDchCxLgfj8/12vI51Rk3ShRHvx29m
A7fV2r2TFzMX4PBRWBKmH9tw56Z29OF6lovSAHNm8J2QpZX+AbTOVUUTE9HrbM6H
NaZ3e7F9xjzWs1KS7YmxyT4O0csFp6SpaCWAB43fzu/yyXF8HZ+8DGSq2FSJZmHJ
3dinQdOWhuqMEDim34y/M0IaLTFQ/kdTAQYGSRnQKugb4Ulw16UZFrFY/oCdY+bA
aFZzsLd6GYmL7SU2ZVw7o1hy6K8Z4fTj2IEUO8lnRojXAblkJSQFm3rnuyqfZswt
Y6jWEUhqnJ+gnpXSCxrwrP7AserpG/J5C9wj14Bn4pm2dYx9WqRMjSRcM37CHJfk
I5Xzl+kTAkEEvzwX41RlwxdJLtMzwj4P0fTAXcTAJudnPPBOc4r2isOk9eJsQ4d+
SRQP9Vxj8Y69RdFMglC7Rsvqwj4GxLLUKGVQTf6ADNpjV9aBym3+14TBb+xoI9VA
NtcM62EUEa3l+RLaykmmGhNbpYsbWkJyTebAr4j3oBsZHquum3vFi1NJqltbaakN
EwTc9m/SeRx2wiAovP8ZkzNceXMhCds6e2dKyD5RN7H/3uIp9R8/0hLtfI5VaJsP
2q7GH9jbxZnqi52whJ9M2+Kz2tpvcfWS2yjUbiTWKyVLKZrDQ2YJl+KVNDO9EP8K
jqGKdz2LsYXcfpePiBH3oUiWCxETjMnc+DaptNR5ItV7fiJFKYvuMKr0uh6OewSk
4pYyG3iLEM5PPcly917Bols2lXG5l70crNAY+2rwSRzykKGOhUUAzxqU/LBEL+BP
haD2TN3+hILGARoOZxfJLvMYf1hClHtjlU3r72zhE0R3WWaLlrXG+9hTSSe7J5Uj
vjHSY/7AeKcnbW/KHqg3lXrjmf2vxSBvJbHnTNbRG4IsOsJ//5uGJHYKqiNQuQSb
fCi6wAQ5lo5dWciqpFDHE4DlDDX5TPpFYmMFHB3qHEYSpVn/wXN2BntrKqEDwUg7
b8qiZ4y0fWPJZYKrp739OnqG/RL8DpxfyWEJjlwkUAnBiZApFHhd1E80SSJXL35r
fROFbrViOVmKlKdDonE20X0FCjhlHCR5AS6HS0MSmnkMvaUXaRjymEsPUJ9qLnJ8
aao3tmOiq/TNGT4XKTanX762oKaMpOO+aHArxPQFsYdkhEB4erCXOVTNC0EMFYQi
+CV/kSxhEWVFvHJT0F/+qVvQIn4N9Sr1err9b3GNG7+2ZMoJJ6/BmR2qAz3/+sRD
nCMGpFIdcbMulEDhlpiVewcy5Lm2/PIyvKZfYgS0Lbyr2RWUpwaIs03kFeW4PJBF
vDtayccwDJ4nxRlHNt3IntyUkbdkO5wXT8cjsbs3VmXqtxiv5djMvOHGoQ0kA4OC
aFJkgywLzSOH5TYMrczx5XKd3V1tWmV1SR1HmA2l1VdnCbCJNF8nZp/+OLC4iiQE
THsa6W/JRA1dPn+f7ypFFY6lQUQlahm6nPsUSPzAurxwvaAIUJB6j/voBzNBp1UE
DflJk2uNP7J7OiwbgVrGQH19BQTOkAo+oRy90mr3thtMiIyM4fCksZkxzbPqfC+O
EOtt0fOSc6v8qwa26fiXXZMTth3gqiS7jpLENx2n74QvTQupP/ZXROyXmO8xGOEL
oDnm17TH/rYxrcWJ8uci/DVz9ZQGgjJnEI1VQX3khHQbnu3pK1ky39+7CEZ4S84W
Y6XaRlEi8lu7XSDJYBMOQvyeJjmz+xUogKn9BnE+wCU=
`pragma protect end_protected
