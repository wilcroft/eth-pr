// streammerge.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module streammerge (
		input  wire        clk_clk,                //               clk.clk
		output wire [63:0] merged_data,            //            merged.data
		output wire        merged_valid,           //                  .valid
		input  wire        merged_ready,           //                  .ready
		output wire        merged_startofpacket,   //                  .startofpacket
		output wire        merged_endofpacket,     //                  .endofpacket
		output wire [2:0]  merged_empty,           //                  .empty
		output wire [1:0]  merged_channel,         //                  .channel
		output wire        port0_almost_full_data, // port0_almost_full.data
		input  wire [63:0] port0_in_data,          //          port0_in.data
		input  wire        port0_in_valid,         //                  .valid
		output wire        port0_in_ready,         //                  .ready
		input  wire        port0_in_startofpacket, //                  .startofpacket
		input  wire        port0_in_endofpacket,   //                  .endofpacket
		input  wire [2:0]  port0_in_empty,         //                  .empty
		output wire        port1_almost_full_data, // port1_almost_full.data
		input  wire [63:0] port1_in_data,          //          port1_in.data
		input  wire        port1_in_valid,         //                  .valid
		output wire        port1_in_ready,         //                  .ready
		input  wire        port1_in_startofpacket, //                  .startofpacket
		input  wire        port1_in_endofpacket,   //                  .endofpacket
		input  wire [2:0]  port1_in_empty,         //                  .empty
		output wire        port2_almost_full_data, // port2_almost_full.data
		input  wire [63:0] port2_in_data,          //          port2_in.data
		input  wire        port2_in_valid,         //                  .valid
		output wire        port2_in_ready,         //                  .ready
		input  wire        port2_in_startofpacket, //                  .startofpacket
		input  wire        port2_in_endofpacket,   //                  .endofpacket
		input  wire [2:0]  port2_in_empty,         //                  .empty
		output wire        port3_almost_full_data, // port3_almost_full.data
		input  wire [63:0] port3_in_data,          //          port3_in.data
		input  wire        port3_in_valid,         //                  .valid
		output wire        port3_in_ready,         //                  .ready
		input  wire        port3_in_startofpacket, //                  .startofpacket
		input  wire        port3_in_endofpacket,   //                  .endofpacket
		input  wire [2:0]  port3_in_empty,         //                  .empty
		input  wire        reset_reset_n           //             reset.reset_n
	);

	wire         port0_out_valid;                // port0:out_valid -> merged:in0_valid
	wire  [63:0] port0_out_data;                 // port0:out_data -> merged:in0_data
	wire         port0_out_ready;                // merged:in0_ready -> port0:out_ready
	wire         port0_out_startofpacket;        // port0:out_startofpacket -> merged:in0_startofpacket
	wire         port0_out_endofpacket;          // port0:out_endofpacket -> merged:in0_endofpacket
	wire   [2:0] port0_out_empty;                // port0:out_empty -> merged:in0_empty
	wire         port1_out_valid;                // port1:out_valid -> merged:in1_valid
	wire  [63:0] port1_out_data;                 // port1:out_data -> merged:in1_data
	wire         port1_out_ready;                // merged:in1_ready -> port1:out_ready
	wire         port1_out_startofpacket;        // port1:out_startofpacket -> merged:in1_startofpacket
	wire         port1_out_endofpacket;          // port1:out_endofpacket -> merged:in1_endofpacket
	wire   [2:0] port1_out_empty;                // port1:out_empty -> merged:in1_empty
	wire         port2_out_valid;                // port2:out_valid -> merged:in2_valid
	wire  [63:0] port2_out_data;                 // port2:out_data -> merged:in2_data
	wire         port2_out_ready;                // merged:in2_ready -> port2:out_ready
	wire         port2_out_startofpacket;        // port2:out_startofpacket -> merged:in2_startofpacket
	wire         port2_out_endofpacket;          // port2:out_endofpacket -> merged:in2_endofpacket
	wire   [2:0] port2_out_empty;                // port2:out_empty -> merged:in2_empty
	wire         port3_out_valid;                // port3:out_valid -> merged:in3_valid
	wire  [63:0] port3_out_data;                 // port3:out_data -> merged:in3_data
	wire         port3_out_ready;                // merged:in3_ready -> port3:out_ready
	wire         port3_out_startofpacket;        // port3:out_startofpacket -> merged:in3_startofpacket
	wire         port3_out_endofpacket;          // port3:out_endofpacket -> merged:in3_endofpacket
	wire   [2:0] port3_out_empty;                // port3:out_empty -> merged:in3_empty
	wire         rst_controller_reset_out_reset; // rst_controller:reset_out -> [merged:reset_n, port0:reset, port1:reset, port2:reset, port3:reset]

	streammerge_merged merged (
		.clk               (clk_clk),                         //   clk.clk
		.reset_n           (~rst_controller_reset_out_reset), // reset.reset_n
		.out_data          (merged_data),                     //   out.data
		.out_valid         (merged_valid),                    //      .valid
		.out_ready         (merged_ready),                    //      .ready
		.out_startofpacket (merged_startofpacket),            //      .startofpacket
		.out_endofpacket   (merged_endofpacket),              //      .endofpacket
		.out_empty         (merged_empty),                    //      .empty
		.out_channel       (merged_channel),                  //      .channel
		.in0_data          (port0_out_data),                  //   in0.data
		.in0_valid         (port0_out_valid),                 //      .valid
		.in0_ready         (port0_out_ready),                 //      .ready
		.in0_startofpacket (port0_out_startofpacket),         //      .startofpacket
		.in0_endofpacket   (port0_out_endofpacket),           //      .endofpacket
		.in0_empty         (port0_out_empty),                 //      .empty
		.in1_data          (port1_out_data),                  //   in1.data
		.in1_valid         (port1_out_valid),                 //      .valid
		.in1_ready         (port1_out_ready),                 //      .ready
		.in1_startofpacket (port1_out_startofpacket),         //      .startofpacket
		.in1_endofpacket   (port1_out_endofpacket),           //      .endofpacket
		.in1_empty         (port1_out_empty),                 //      .empty
		.in2_data          (port2_out_data),                  //   in2.data
		.in2_valid         (port2_out_valid),                 //      .valid
		.in2_ready         (port2_out_ready),                 //      .ready
		.in2_startofpacket (port2_out_startofpacket),         //      .startofpacket
		.in2_endofpacket   (port2_out_endofpacket),           //      .endofpacket
		.in2_empty         (port2_out_empty),                 //      .empty
		.in3_data          (port3_out_data),                  //   in3.data
		.in3_valid         (port3_out_valid),                 //      .valid
		.in3_ready         (port3_out_ready),                 //      .ready
		.in3_startofpacket (port3_out_startofpacket),         //      .startofpacket
		.in3_endofpacket   (port3_out_endofpacket),           //      .endofpacket
		.in3_empty         (port3_out_empty)                  //      .empty
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (8),
		.BITS_PER_SYMBOL     (8),
		.FIFO_DEPTH          (4),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (1),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (1),
		.USE_ALMOST_EMPTY_IF (0)
	) port0 (
		.clk               (clk_clk),                        //         clk.clk
		.reset             (rst_controller_reset_out_reset), //   clk_reset.reset
		.csr_address       (),                               //         csr.address
		.csr_read          (),                               //            .read
		.csr_write         (),                               //            .write
		.csr_readdata      (),                               //            .readdata
		.csr_writedata     (),                               //            .writedata
		.almost_full_data  (port0_almost_full_data),         // almost_full.data
		.in_data           (port0_in_data),                  //          in.data
		.in_valid          (port0_in_valid),                 //            .valid
		.in_ready          (port0_in_ready),                 //            .ready
		.in_startofpacket  (port0_in_startofpacket),         //            .startofpacket
		.in_endofpacket    (port0_in_endofpacket),           //            .endofpacket
		.in_empty          (port0_in_empty),                 //            .empty
		.out_data          (port0_out_data),                 //         out.data
		.out_valid         (port0_out_valid),                //            .valid
		.out_ready         (port0_out_ready),                //            .ready
		.out_startofpacket (port0_out_startofpacket),        //            .startofpacket
		.out_endofpacket   (port0_out_endofpacket),          //            .endofpacket
		.out_empty         (port0_out_empty),                //            .empty
		.almost_empty_data (),                               // (terminated)
		.in_error          (1'b0),                           // (terminated)
		.out_error         (),                               // (terminated)
		.in_channel        (1'b0),                           // (terminated)
		.out_channel       ()                                // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (8),
		.BITS_PER_SYMBOL     (8),
		.FIFO_DEPTH          (4),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (1),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (1),
		.USE_ALMOST_EMPTY_IF (0)
	) port1 (
		.clk               (clk_clk),                        //         clk.clk
		.reset             (rst_controller_reset_out_reset), //   clk_reset.reset
		.csr_address       (),                               //         csr.address
		.csr_read          (),                               //            .read
		.csr_write         (),                               //            .write
		.csr_readdata      (),                               //            .readdata
		.csr_writedata     (),                               //            .writedata
		.almost_full_data  (port1_almost_full_data),         // almost_full.data
		.in_data           (port1_in_data),                  //          in.data
		.in_valid          (port1_in_valid),                 //            .valid
		.in_ready          (port1_in_ready),                 //            .ready
		.in_startofpacket  (port1_in_startofpacket),         //            .startofpacket
		.in_endofpacket    (port1_in_endofpacket),           //            .endofpacket
		.in_empty          (port1_in_empty),                 //            .empty
		.out_data          (port1_out_data),                 //         out.data
		.out_valid         (port1_out_valid),                //            .valid
		.out_ready         (port1_out_ready),                //            .ready
		.out_startofpacket (port1_out_startofpacket),        //            .startofpacket
		.out_endofpacket   (port1_out_endofpacket),          //            .endofpacket
		.out_empty         (port1_out_empty),                //            .empty
		.almost_empty_data (),                               // (terminated)
		.in_error          (1'b0),                           // (terminated)
		.out_error         (),                               // (terminated)
		.in_channel        (1'b0),                           // (terminated)
		.out_channel       ()                                // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (8),
		.BITS_PER_SYMBOL     (8),
		.FIFO_DEPTH          (4),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (1),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (1),
		.USE_ALMOST_EMPTY_IF (0)
	) port2 (
		.clk               (clk_clk),                        //         clk.clk
		.reset             (rst_controller_reset_out_reset), //   clk_reset.reset
		.csr_address       (),                               //         csr.address
		.csr_read          (),                               //            .read
		.csr_write         (),                               //            .write
		.csr_readdata      (),                               //            .readdata
		.csr_writedata     (),                               //            .writedata
		.almost_full_data  (port2_almost_full_data),         // almost_full.data
		.in_data           (port2_in_data),                  //          in.data
		.in_valid          (port2_in_valid),                 //            .valid
		.in_ready          (port2_in_ready),                 //            .ready
		.in_startofpacket  (port2_in_startofpacket),         //            .startofpacket
		.in_endofpacket    (port2_in_endofpacket),           //            .endofpacket
		.in_empty          (port2_in_empty),                 //            .empty
		.out_data          (port2_out_data),                 //         out.data
		.out_valid         (port2_out_valid),                //            .valid
		.out_ready         (port2_out_ready),                //            .ready
		.out_startofpacket (port2_out_startofpacket),        //            .startofpacket
		.out_endofpacket   (port2_out_endofpacket),          //            .endofpacket
		.out_empty         (port2_out_empty),                //            .empty
		.almost_empty_data (),                               // (terminated)
		.in_error          (1'b0),                           // (terminated)
		.out_error         (),                               // (terminated)
		.in_channel        (1'b0),                           // (terminated)
		.out_channel       ()                                // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (8),
		.BITS_PER_SYMBOL     (8),
		.FIFO_DEPTH          (4),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (1),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (1),
		.USE_ALMOST_EMPTY_IF (0)
	) port3 (
		.clk               (clk_clk),                        //         clk.clk
		.reset             (rst_controller_reset_out_reset), //   clk_reset.reset
		.csr_address       (),                               //         csr.address
		.csr_read          (),                               //            .read
		.csr_write         (),                               //            .write
		.csr_readdata      (),                               //            .readdata
		.csr_writedata     (),                               //            .writedata
		.almost_full_data  (port3_almost_full_data),         // almost_full.data
		.in_data           (port3_in_data),                  //          in.data
		.in_valid          (port3_in_valid),                 //            .valid
		.in_ready          (port3_in_ready),                 //            .ready
		.in_startofpacket  (port3_in_startofpacket),         //            .startofpacket
		.in_endofpacket    (port3_in_endofpacket),           //            .endofpacket
		.in_empty          (port3_in_empty),                 //            .empty
		.out_data          (port3_out_data),                 //         out.data
		.out_valid         (port3_out_valid),                //            .valid
		.out_ready         (port3_out_ready),                //            .ready
		.out_startofpacket (port3_out_startofpacket),        //            .startofpacket
		.out_endofpacket   (port3_out_endofpacket),          //            .endofpacket
		.out_empty         (port3_out_empty),                //            .empty
		.almost_empty_data (),                               // (terminated)
		.in_error          (1'b0),                           // (terminated)
		.out_error         (),                               // (terminated)
		.in_channel        (1'b0),                           // (terminated)
		.out_channel       ()                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
