// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:11 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ax5XUne956x0ohUrlvCu7l5/gsIQXQ3b/xANity1Hflpsn+uOEbBqO8wh8yJoKds
6/w+MO7FWyblaW8qyyXUp0vUC0cxAveGwb1rkK8jYnH3S3LLZjKWBhQs0dDO/xPy
/kftQes/tDg2iOBZOAPfjbW0yA7Sql5qs+Ozhcjqpw4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 324336)
84gSkvtvVIrlZqI7Ce6tmvcNczf/OiHLm3Xt4dMSknh5r3vE+RlyLc5WTEfLi3JI
onL0TybT3Wr8TMF8Rl4arW+O2OCH5qIIJB3KfulWzxP2DTtsXwfKSB8eStxNnf3M
xsYGSwkmXqbzGs0yYDDA3mtWE/uPe+nvC37ylHl7+8kmdDiNhucT+KZqDhtS0y0c
0015xQpHNJW29JUBhjQaqFbpqhuNNrIPT5XLlTL39w3u2k2QJU2pvB+Ekz4XrcvK
aLA2aCYQR5VgFy0r3F8+QnmusoffcUf6jRKpLan9m5Lz1GaY79rrOirKybjZNMa8
MF8ydZt82feZWEKVGDJbswRi60PuIaWhZGCzHAp5NTIVMgK5HJltw/rzMlAVR6fk
YtYQN12SxJ4Om6iYPJqpcQp69qGZ5qe3nlNKsZm4z4rNLpM4wDGuQ/qeIDQroIGZ
VVW5kMMftTcnpyH/MQ+xMIoZ6pR02c2xIv/sDJRzt8o6cv1g027oneQVKaXxm4vP
FyNPrTEBYVJrVFgsMu0wYVh9oLREvC/fDvyclXv+s0lP7gRY3l6NaZadQO2xypgJ
u8cK2+4KJKLbAG6SJ77qbvARJbmVB2VRZWyHZHYb4Zdw27nDa4s4m16OYFHRlTBg
iCR5mkdbtEw62oajqpMt8ZI1vDGJGkinsn35ZeV5PmzO7z+5BqrBtT+XlBWEACG4
n/xELnukZSXWCFdETxzZ4oJLFZoQcTTYSZBntSXynL4VbkePFk3K3WgkxWk6Gryh
FO+7DwIAc8B5JI/FvUHcMx3kKMOjOxciH+0fIyWgj047oSTDs8gTosDWhgow8mT1
UFIT6d4ui3tMJ5i3xO9qAZI/EFJLAi1s5sNT+OEzSGlZNEF9T61QVsp4l1jaqTX+
MKE0RPmg2y3svUGg3sLMoaO2pOxSQUP7zNrTXBl5uYvrELXUj6qA2rjNv+vKiRKO
4/LTvMcj9DvE9gwjtKUb6gprZHrgYzuWoRdzyiYL0qQ1MJck5hl55GFwiM8Fv6se
wfyoQwvBfkWstuy5hZPxnhTVJHpceg0UYAaiWsPadSOVqn9em3rbSnMIDOY56+Bf
ws3WCxuUIhCAq69twErnubkWibB1n5ZPCqskZrE7dAaQ6bi/stupGyLxNhDR73Y9
SIu0J2MhnAKd5v4sODirK3AVxehIGdXQuHHs7Jp41yYfYruBo7kpGT3rk3sG7cHW
uAlZUPQj5QiL4fnphME4cQpdp0u5I183qnjgMTLB2u4iR61ndt4lMPv8Z2bWO5CI
XVIXyeBkaPUhzq0sQf9KZT8QDjBp86EqBrV9GugssQqfB603WrmZCfS1PxrDKHRz
ez8v3Mt8ke8gGbDbQirKkLbUIm2toNCRmPy+A8eqgXqeWz/q8a4f8r9ZLYl8MSO0
Meiwx6bYJePxMd0ciGVa72FLcPyWDgwe053qrRIYKGnx9NwTcoqvSrJO9yvH++gS
oZ57LfSml2X5D8CrGzXxMmaGHNBDlwYUUrGnDC8XXUdq9jWuOFXGtSHX94r8wFsm
zsAMhFong4JfXOikXpwkukE974dP0QUMN1SBkf4u+4Psa28KIGhmmrZz3jo+4BpI
bloIRzBd3LSTt+OtVHUWRYFqjbl5bwWdDXdAP7ToW5q5N4prXVoOO4FxafIKohMQ
7PsmbzP+5ZGuO8kdYmpiIaRGymX9UqkKgAtlODr7ZUu6zejwO4wqbc99NEn4X6B7
R6lBTKAJyGgo1iDhpgjq/64nbLXLtE/KDkm6n78+H61zJzU3ofy/bLNUpBAu2aBD
Mx0pxOtB1rrkYEVo5TrCno7UZxAR35JO1snagbnQu0JSaRaBtv3tYs38hsE5qGtM
WSO2BlROQxc6eCIRi5nMvqN28TGqf1xkj+BIKMAfXmSykSChKPdjSl1prARiGySq
jf/blSHYmK6z4Q7Iph5ff+xFoYyZwPMomEXUZyk+wv4CaAHiCet9g/v7W6z/8rNy
86/KZpIbLs4LFtuWOTwRh8EtrFZQLAOLF9aRAMcz25QFx93DFGW1g2RkTKPVlQGL
RRc9zqtsp24v+TyqlFUhn3QAQk3dUQcS6F87koRl1SCCQXJZd7IPLjlKn/0zsd8i
dz/u5p748tLaC4vclUHJ03f74BBZmN5+7AKyj+1iBnbLiZGgfmCW+MQQtyPPSu1E
+gKlsiUOGF6mWbT4FMWr0yRH+rWcDtslKfVXcp1zsIgqUTVgcrov+F6tEwLuWHlK
Vq2ExhGIEj6wOEYOLoh4n5DuioVLWegrYhSu2Q49xs2sIYoIZYJcdAZup8c02x+U
4z0qXV22eFeduiCrgh21T+04he9MQ1SOAtnngVdXfSPbRqiISQcKvV3SezMqBbWN
e/mAN4Mzz1l8+AWsCxxIIY0LOgvfVGS2UO0vsShDREKnfNVLLjdJBjBBY0xqfs6T
hXUWexOrwr/E2o1tR/rnUzlZylgfqRtkC68qppIIcbcJQFW4q0M3vRzseDwEzbp6
1vpTzvKKNgAIzyNkdryD17OjnwusKp1MrW6cfueOebCCVik1TF3AEvitxw8hTjj9
dmREz3Qt39t1Mmxg2FINp5acJ8vL3Syr51AjcoNRMQc7Xo8LxxAL54VBOL3DbCwH
sSfJzP8J2IwuYU2qruxv8LV/mCdL0TE3g+fbY/C4DiQmoIl8uVG2SlPYi2cX2m9F
aCyd79sH+41plqDeutOKwOKGEAzH4p4G0c2Ta/94qmljMF2aDCnnxGIoZyHw3dkg
qKdXb/J+llDLTpLoX7ijiEFutGLYqPwUekdy9EjYWR5DXl42nmDHiaRrCovptvwl
HXUdPEwKKI/iKva+g6cgD/O5VeYAqM99eUohRZhBxMfd54ZAadqken3v5gCjdjdw
ArnUsI+r95q5xKAQffQNKYQgo0oXZ0L6udCtArcKn/LKrxzbAPI8h64cMafxNFCp
D2/M/7NgZ07q2IVrqA1DKlS5d0tWzSuD1zDuBCNHXE0rJND0JUjqaLqaBMj2U1WZ
2fs1anfkK0KgUagazpJmFh/nNPH4vT3yt/ABCvLLJH5D8XJwJkn0zA53jumKVlfj
Dk65w/rM67waQNCivUcuJltNIZ2TctXV5q5mFLaeahoc8TkaurbbccOMNMCvM/aI
4ojOPPTJ3+JCs1e+IUEbfQXlJz5qFXnGAN3EIISXkQ8yQzivH3T+WJPhhCUXYuLm
DzKEP8t2TZ3Nn5cvdSOHuocKisPn+Sgv+UxLdm3jRPdRBP23TsMCVn1wbTRDJLAf
TWZa56UzofDRqjsj3c8ecsvvdlrkYHyjG3JUZICt155G5xoviOJoH0zyVq9o3YoE
2zb6LLC3ufiQUXwx/Pt2ahzsGHt6kIjgGmdyWYfOrzmalrn19nyvdvnlbJuYbZ2Y
CQVZe9EiwJL4vxyr7Wv19usZrqS0IyN+QidAaAMNKtnHMrkj9l8HbLLiVcFPGPy/
KjggVropH4X7h+HXBV32JW5HDC3cxX90zUfqqLnL1ANkfcGGTsGx9oy+nN49tFgt
OK9dgLqk8gijvc6LR8MqW890dkiM6uFUnRryasuW8C39UzBFfkUVyv/QD6M7zn1e
dpow4CDGFcYirkLfrKh1rRpQIhve0gNryHqRp0kRbgsx07kPk2Ffdb+YFljy/2jJ
efRQoXG9JGX4/GOI28uCLGXyndyI0t8ZEGsMoAepn4WBdl9hl98R5k5NJ1JGB26U
IDGF3f2cLmRPW6Zk5T5ZQy1IRJ/jTwyP93aJfkdYTq44mkP+Xls0As4i1lpz4vFj
MZRwQ7vkdKxSQBn+jzh8tzHVErZ/3FGOL5i8rXag8CJXLLUaYi+m1mMo/ivtEjZB
BulDWOrCOfCIf+y9JxiTJXBh5CRvq0co9Km1nwkKSg1ZfXmxJAYu+UUK4mBFr02Z
LV8lAzaT0nEKcnKDbaz1G8USoRnKgho+Oz8uNjCV67i6br9nRCLdmqbh328cIBTA
itgE6w3PovNvPb09DnoHATjcPmW00JssmoCm+5LYR9AL8ZmU/0JD6D1rYdmiMc9N
j8W6BBeSPELUIwqHSNCUfOWTMUh5p33gEtZ90F8PKFR+cwOZdGfMKa0vV4/55KkO
0J+iEuicnM4H00kNZQX1ShZWd/W2VBkqxKXP2C6UeQs4jmxXr/A+Zk04diFpGziz
AFpeTEmYVRmC3rds9x1wgJXnw4l2oCFjJ/diXxpUl6L97oexP9NPIoDceOxz1gsg
5N5yUJ543TU/ekH4sR3xJ33WQgvyN4Pn3ZPq7OTrrZuJB3WMJUOtcWlB19zPGZA7
cemhzO//wpxqqvMhWpyK0uqW+VKRjJzi9quLJUbRUeYkF6d4MueOGMRdIW6WBZIp
caWKqRVvCd/AlafvJW7EpUeqEYdzqpV9PJsqfqYkFr9c7H1hbEFoEzM2JtF+U7wg
X38/dMtUtqIuNEbGUrxMQ7EnfPGgnp944NAXBb5ED74pBrr6Vq2LDmGomewrfgse
LvqjsTX4RVeFBZtehaeqq25s0wmQ9w0Cr2n7vCBMqjJEIi/qJupfoRjcISm+tAwZ
BQiyNEc6jfADShF7numDwpOFGl/XAiAMIOPJX4EbXxoECo4GBBqN9jqveALEthEs
yqy6UfxsV7c8RTMx0hHOVPbIdEn23snAfnG0lZwQP9HpFZVuhXkF9gvwabHAF8q0
1gQhm9RHYg9DQyPZ9fz3Y1ycS141nVUY396rLlVaZOTelP3ZyXZqSu2SsmjdkmIB
QrWlEzB/hngKCbDvy4YAUTd3S2SrQo/zGqaT/8xtWgYakW42qSY62dYvREUGenIR
CyzuYijr7G4kdQYLhOZDcLx5d5aH5UeSQHVGEAdFn473ManhT1aVhjrmKpdbYU85
AcSgsP2hu8CZ9n9Sl1fBEyQZv1q6jVJDbMIr0Mrwq9Y4M224ZrbfSe/rw1prEQYq
dWgwRH96JjcVH9xl7xA5+07kF5JV3L3yaNj5acAV0E3Qf71nO1D/ciZ0Q4mCUqc9
Z9xxD88gJxQKAC52aPDpud8RfNDm3lPLJ/+EEtkmRxQEWoZ7RjvN0cANdcInoxno
Y6YxXji4xjua0hWe3Y03PYODFvYeurq3b37vR5j7vgyN24HETgjTbJe3XJFddVQy
2n+jz5/XH/91bS6pxqF/8UZUfMFBWbd9rlqjnXPGGU4oUjvzzGmnxofY6Yqkq5fW
ztYERfDZE7gOCcGi7ME6xutq1fuBd5RhntukKr1YCLlnq6A2yQK0fGSHL7gdotWw
k2i+OFp/6LeJnUztC9seCIY9mKg4H/sEggqPkE5ASGb2eepmO8opA09f+tJQcdcs
6QgebLcv2Wlwf4BD4r0Cup8BOeqXP8HtB9NFLe/qsu3+w2WXTO3iGoCTxHpTAwXG
m6DcDC99i5s+O8lmudXX1p+NkNhhkM37JV1CmbwSSd68e89DsxPf6LirhEhY+1rV
UI8f+stDMlbxO8YrojFFH1F9ZLmF3UPFMPtBwSQf9um79nKe7LXGOFLSGqFbSmmh
yWeyde/m+DJljfbJW0uNrqH50oW1nLAehPiPxV0Q4RtS7w/IMdvf4PBvFvdwqcnQ
ajH5XUjCZrfSgw6T18lGJfRDtbIBkfEl4qFCRmgUlJ+xohgUVfaD/KekSUe2E+Sx
BiMXEeaQgRJwj/tcCi64UygdbkLikUlqT9sq6WyXWLggYNsPzmtdocAd3mgg695Y
cjBKI78ZqtICxkeA5/XxlAlO85UyHP7AEia4oSBtXFN52h285zyVSo0rW8Ao/p5M
xD4w3N3sCdA+J7Xf31wrTZoAAASJtnwdF4ji5HqBqcQtOZ1WdnpXwghBnjuYriXG
0wHr3+yC/U323vWpR7acDxHe14xvfaVb6MQ23UvHDdRyDoZaaujB9eFPWuQ0CLxF
9Dopuur7SPAHA6rUUnoR04UW5McArxharE94sdxPOQnL/dgd9kLyGj4TEpxe+5iM
EhRXBTA39otJUaBjcAK3EFL1wvl2ml2iL7P9uHxaXUmjklFGBZRnkWC3uZIUzEs5
ceO2oA30Q3jkf3xLgHAgMv+3E6TdjGGxoQhrzrZlxG7AXu5W2OSUVFtKJ7ROKhHk
UgU2CZMqoQIBcCpXIgJj6EfaqLVvDWRDq0+L4rxy5Q9o+DbaYOwosW0R+7D/iNXQ
p4A6MtkowMATuZSoQu5/HRY1ioGW4ZKR4nOouSLbCmg8s48oY4Wlvvu9Kkt7Djlr
DazLRCidmUibvHHq3rOXzFLowmeYGxHFH8B/c2B7nT2YbAkMenYVZXKb8azVxC/G
NKZemDfhkZqHMh6ixUkTnnSv+VhvsMcZZxwQXGipD6bWL7zkoEhzdud3X1P4dmWn
hep2gpKEghhu2k1oFADEHEgNKDvNNqrVIcUBRkqiFBm29gtzu3GK1J30KPT3+nDl
oj9mdCNsR0CAiMJQXLjcx9ovGh1LhBR/F19k10iDpVh868wglSNFIz+hU12Oq9Ft
GcEkj9tH4dZ5dqVsuB2xirEEbS8jFBixDhwgtwJtobipTIHKRhr4GdpqJ4gAhgrY
hnsDRSVaRcc4zdfTqYm+/NMPf/FY3MzDXci9XdGV+DGxzY1Ej27TtcUiyAfmel1Q
1rkNSD5Ucu7AWrQG13Y+diwFbao19uec31TLyOt9VqGi6YloC2JU5SvI+dQ7S4xB
dtso38u2LZhH1muF4uZjCtD64WpCJirs1dI0xII9O6J7mM9Xe3NcPydt3PRSfFwR
CXBr7RQt8k5fS7qGIc4/u4jSecI0hb2jjcZYd/WGRFvRolkAYNh8HsEEi4CdSqrH
xWx/3EH69lU863WYoUmH2sin3yqQuoFtqpNWSYHkpI2TYldzl3BscJd/uUxJ7kxP
xhMY7tJGXn7bZnsPR3tALDL6aaqGYpBqpO/heNIZuZQ7bOCzZyetNjkeqH5uqr0t
uT1+DSzam2rnlEZOYq/8aKuXfRBZK9loDqCGwuxDPsaiLah3RfRlNDZE1LQQAeM8
fTiQD4VjxZzZpGGzt4/rsH2Wu9sunkeQLNQpZrYhKkMZIqlMthM4dDUhlI4vR2xv
bf8OV1khfA3PX7UD8cT3KSgiEzEsU7U8GUIfxWb0RAO4q/Qme/p6lmtP2fMe78ar
dr7kRNlFUvV7IYLU73yWwY4mBJP0JmJkf/87Mvqyd7f0kzwQY/gzTx58TKCheOox
6ewvV7zkXLY+7S+tfsXAm831eDD0vbuo682rkhUad19KlWGztnzvfp9t4jLQIp8q
thkGMC9Svfr5D5XdR7/D7IE6ecLpVZeqVQKZPcVHUkBJ+CCqPW4Q3Ncpn55Amx/j
u0Y3FFbnMhkzKJtRD/fNHa1Fe/rcyWAYwI51xqdXMMjKX/zDJX5xESs0EJSBYeE7
PNdbt2Wk7hJe+C37N+j8L/pasohNdAoNqXyXtkXa6FRovenwRZmKeLwMr6o1/StU
zE+xwPm4x6LNAXWaFFz/6M9FPjTqF9eFi39YfK03yvIqaXosU8ngRvTaAlnC3ihC
I/WiYEk65VerFRQo0KGRuRpkRwOwnWbkDcDyH3PW2MLITa6NNZzGsBQrvcY/MM2i
VhyddjBVZ7RsCqoti0RLoSHIzxBVBsuvIBndqR3YXVRWpcW/STjU48AynV1/BnW2
CjLAIPaZXakm+9g2/7b6+97t5YlVrniBr26MV6+Ss7hGEgA4KP5+tuggljFLZMSH
Oh2cQw54UbY1wan14tc1eLhNOBm3VQrnIaxogQOcORxlhcjeWmKnhVyFz+R8ZVY7
zXoGXJDfMQ6iGl8rU2X7jO+eGUDt3XHpIyrzuefvkpsvLoJ/4nj22Ndyu/VgRTzr
37d//v0rsdeP7YwmNa5YWXKk1ZbPuqLfyDaQgIEWoH/x9ox8hGMMWCVQlyajIuML
MWwsVrLZjnIFFbDdU0nfu/IZEZVplKykbdJJd2JB39U8mRc9ifvBJyuIh7z1orto
5lMr+Gaka4ZLo5iwQwGGwyo98zkoQN1sFfYFqOPOfLGEmnQjLdC6fPovlooQtT8x
6sha6+SC4c3LT4EnR0hwb1AmJaEhtHjsRxiK6BGl9MHTevIAVsF6B+/UJRZuOc2L
S7h5/r5Sc8BqYanuyjalTFxv6PbaTpHxkX5kZ1FVIA63tu66RNK1ulJQKz+MVMMz
vye+QLhHdIBZ/L8YQC7vvmRdGKav6iCk6/31lozl9dr3v8AqIuQ1+dQurjszRCde
xfqHC53x9FmPpoMhTMKxyTdnchSeKVN/3gQXrxwppW+/YXC04RuR+yvcR7jYMeDr
jeHYshV1x35IwveIp2dS2bwwmzhY+guKOVbK57v1Uye9ah3eKzK8cmyd7q492q8s
2qlurpVK/S/usfnmzkRmur6WQ0A7PpUL7Fa2raOpk22Ls+vbzkmCyuNeCIpobUNC
zJFqTJpLNvNBGD0bUFOU6XGbwqldlXpFHKe2xhP0hRCQ7b+SygVrRTI7+zyRJc9/
PY9+a5oV+bVhDcKWlIxbusv+/WiShsCJE4mHOCggkoL05VeiPHqz10CCDL8YZigv
2UyqnfmWm+sCGiMFjeq6OsohV8M7ul+Xu7NQnF2QLF5PQzl9VLp757NIIt3i29y8
75Qyaz4f8MBrqzYmHP1hKS3MajWUp1c7BFdgUo4aW2QntpI3DVpELXobZp2/w6DI
51R0gUEoExNhW2ycsrnHM6XJUOXqu+tGspPBA4G756kQmvy/PM5RGbKyQZXTGtoP
wqbF+QEQBMgUPmbD/a3nPfCE5ST/IUw91rMZybUDw5FuuITawgHh0pc/qNguwBYU
SAHLxUbo7sFD1Ln3MUn2oQXCFaYDt6kCSD9UBPtWUvE7jU70lhKFg30rqwcWXg62
hGPxQjbZgSSNvxCIKGQWCo/1A/KF5NZxyKpDR2D8ACKopCD4bAQVdZKvG03iqfn1
38T8rdYupL0g2AdTrMBJR0HWg3BLxLx9vlcjUUEqp5XrpwIKfqLOQy0lPL/8rvi3
2Q5dSta+1k4EN/3bAS00M9Lrwyv/6dmRYaniAtjWn1gYzHumNOmeCCC0fGEDlvTz
myAFfKeVG+Ug0VPUL4cLYoSSaGj/WmK/qbJEq2cEcGHy+Xb9P/z1dnPN4KkQLlnP
fDn+tskK7CMh0xBVcJIgn67GHxfe25I+qK7/pBbxcJCjE1Xfv3g/3qJ52sVAZsEP
mOs8FezmRM0O+2s+MsJDUo00mMw5kekaCIL8zzb38E8WI/6Vh/ofIRPbqRyRdQ97
8XSAYL26FWSSK4khpjaWX2cSje3IJdf3FQbYWHdH/890wHzG8iM6CWPNv1eJ0WZQ
iBdRiY+iZqttsSj2NyosE7gdeFnzsfY52ZEPfS6+Zq38ooM9MdytJOU5YcqkMQdZ
9KGU2ljieOmFRtfZefDbQ/Bo3uKtDxQSkX/J3eVIMnvK1XtErJMxXl1roLvfSzkU
IUNfcIYFrlTETKT3gliCzbxtI/Rc9VgqsNPWAIgsd9Lfp5HAR6CckC9tkoAnS2b7
Z210o03LxYymVJ4URRuwembrHd6d2gwouJN9jM4UzokI1pglJd/2MysdKVWUX3Hx
jdiCFsKYKmmaDXaL7Tnarb97O6sC0AzgnP+pVWcIKQmZP4ClQP/iOwW2/HxyAyDa
YLf5IcTVZyhRD0Aeq+2nY7EL+GnIkqxVlYpcutiTgsB0Bz7siycP0J4/+NysyFkZ
p7QfTPIWaQ6O2g1anKS1ea9o2EmhCrvywpYISoMLply2BNEyXT4IBw1YNpR82ZJk
fwjRKkPPnx5KsG+9qccFNA4s5tKW3SGe+CmnoPGEzZBHRRv6ABQLfnetczeQAYdQ
b1NclUKVcr60SvzALpOdyEBIxNXSBpnOoCJHNF/MYE7R9Gbzv9/Us+BUCmLstKnk
rZ7lCj8gKhOI4N9A3UneEpD7+gQFecuIM6J6gy8Bg9IBuuDIR2MQ2lJEq+EMj37n
Ztdb5J2AxdhRMZcXa1QtZTw9SN2lpq2qUdz3YOFNTQ+/g1tXf6W4Mf1zfuhGoay4
L0v+8LmqfXab2rL+XuHux71uNuNt0F5KcEGPySL/urO5sdSu9F3ZqNWAdeJAMzXh
1g1VmUMW59GmLarGwDR9F52vrwpCLZTCgTcAr/AVWnAdjGJ1V5cmyPKs2kuRhcTX
0HU0Jw5uBNO7yWl1Ne6bV6f5WmOLtrXhX9yNlE7599tVhW1YrIXj+PkDKEK0H83L
vo3CFPk9EhHoW468V1LNyQwFxKm/QowbXqvt0afmZJ+KRwDBXNX0C4PoGhNJyYqX
dqbqqCtvYZBfCCdxKBq7IxdDE9FhmGEUZ0D8WPRzXBe3XkpVoJhjc1p94yLoJIHj
Ro68vPcQp7HGko+EOmjHB3DVDo5HzGCm09XF9BeWXzzKz6IgCSDwELcJSwR309gW
IdDoZr44WuZdRlI/xhVOJk0RuhAB4WuAuarhDTlu2EVnH3pZNWZVR1qs4fZJNCkV
1P8BlZCEoY/PMWRp/HDcgPo7QZ0S7A5aWdXOq6RGSsLbjr+lbLk6sPNbZNk5oPYw
snzrUvYOkwmLUGlH7AADuYUcrUIS7BOnXyGlE8z+D2FnmY+HZ/4Hf5NUUHJz15Ix
R9BbU6yhaqGIGobxYyG1xjO7P0lUja/d4JU9zidmy5uWCFKvhl7hHEh44JOxtUMg
SCHPGN5bR+0t4ogyLX3/FwFiOJwIZL+WOj81ZGXqFy0zD4KUui7ZTFxfJdQ9QwJI
qCr3ZR+oO/r6s385xs/TCmLlMiMJxZwTNjT6KKRbhe2MjJymsRSvRmI2BPTsKW97
ZW17IH6p0gEU6WAV5FJLeIS8DKbMNWqND23pJHk/M2QI22TJdKZqiMsACexDapla
HQU55JXW6xc83Kg3oACEIcGjDbyBG+0CJ2gQ5wIxB0re87AJCVWierXb+qlBlyMh
z0GJpF511awdpETPRCpC0fMmUYDxjJ4eCGiHSidZigMmt4+/jfmNmJLWDQnY+Tw3
+2dAbvhlhA4MDQw6k0dzJD0lhxB9vkY5Oh8OKZmZLmCYwsu2I0FKJzrqgfZ2pKR1
eENrSIDLP5bQcUwckH9XTigqebQsXJqouByB2ldnW+Khe9mI+8PGIzXRTAKu2/Gv
va+qtf2DDQ79wrynCwXYRF3EzcEuiuK+hxsDN15IcBXnYEUPuRJz9OuPWmNOW1ZA
3++DeDax8nar3lpn8vCzmeo3pvvh+ieHlD0HhYv7gVhJijDdDuXoKPKKE+45dplR
bLxW3Ve3IHRyOZ2MVrT6QsHf9vr5QxidMUEteOyadZzHWop/Jz3dp8t4ML9Fwy3i
3SZU5VoCBHmTZSJVfO9Ta14+kHBOBgkKSwdZu9NapLg4sv9W63al8OgJudSlrxPi
/8Q4sjRPdfEOVRmgSad5jF933Y8e6ZtOgjqZoZhrHJy3mM8JmWcSlvUSomzJsyn+
11JnIMA1yK9QdxAg1RW2n1VM0yxZCNrnHkNUo9Fv466OqCBITVx7RgpmuBlN3+B8
23fpBnVLlDWL3MxkiH3C/SE7UTxVIpYQciigmLToL8Jwr1oDAAouaqTRQ6vceHrb
hdcvUpT2YYAizeC4B+lwyJDRZ3Q3wjHcTKzM2/tplTQMvX9T2rcr8OPuJpyEKrX3
FKHJwF93MfYPAQwyV2TMkVTVc9Pha5tRc5dcqiHMGsnXq5I9B8p1eQJgBI0LvG80
YHbHH6A6hFOROzJjngThRkyhy4OEH+0BJ29TRp94NS5ihrjUSBclC7oYJkqMtKVX
bEthDUJImTNSMSrbCdFVKU8tzAFVq56X0dPFZ/vWYRAzDDkKt2HfHZYop9yoMXqK
nr5j4lzOQH+bC48E8WjKoLZ2ogUOYEz2xgU2OtVuNb28uK+ZkQmYQiNbIv2ufuXf
nfyiW+46XzO0/tI7hXODCzRt7c0cXKJR9vkanMg7HdVifFNVbqgVJ4Q7v92SEnxF
DBDnhy7ZVXtBqmA1W4h7RMq/o8Zzv5jtDqHjwRrbAfwrksR0K7PFJMSo2nKXyAWQ
kPBuVp3f8eEEwJlDAfVPfsbD6l70shpDv5PkPF7gK8eEHjd0ewhmb6zFcEf1ul72
kcmTi4BwCnTIO9TG2iQ3qWmMGnGbqlzs60Fc84JnXu4Hvti9x+3F4gKQcO9TJ0qJ
jKx5NHYz3rQrHI+6kNRK1w1JOGdP4eK/7WNstQ9qJcjfbyorzQw302OjeFiLYuDC
EMGk0H2vfk8BIcdVoxCOpU/dhX+soK18w+OsO0WhX0eXJh5Zm2RDy41RsbwmO6LA
thuXkvmtKATVeZrOqJlW0pYxN9s4W4d+py+6lJ20b2+UaKbLwyz/0iRGs7b/SJnz
5vrU/wmNQwe0lCxcY8bT5nNqOCpJh/KOgZk4wmpueljR2OnA4jx3vCY4mLRcM8YO
ar02gcAibQ4B+yg2K+RQLoFDfMZp0XA1jiZ1/aGM6JEFiZz5AhPxojSd0gpw7NC/
cEms7VvJZpaZFAAsmyCF0+weULqUHJKa2N+15Rx2S7vSTueBIhjZWpeE2oEQXCPS
yaaWZEKcb75yiuiRP+9B1vlYMQGVg54tD/7XcARnTVYJ1kyxmsmz37nVcCMdLYgO
+U7qwWzUTaL/HWjFghlgMDTVLhmwo/+BDayjLp/+5FlsOsgmD3bo6taL8Y7y8qKh
atfZtKEg1Gr1Fdbe5mIoEvbi29vobY8yx+htHMCUnnfO6tsakKMxtPa9Bu7A9n3/
wq0tb2myU/OP4V0Sog/9HZNCP7kzr0Ffl2jki2W9Z0hQJ2yRJaenBMVMlXAXFevh
CG9VmA7pKBx8GhGVdqUk2OpSF1gP1mhtaeaKovTyWVGVsE6ONvtUt8RU3cyHcut1
SUfHi12FUG0dWOAzFFBxJTuXx0LKkM8J23GybKsZ/SXeITv1Se3krCSZiaqG8OC3
mn7Csf7hm8/ppLsWIvgBnvbitaPSzJB4nhgxHpISF11fox4gzXZdnXpTxwdr9t46
tL+SjQZFFY4/+euamJBrr76U4ip1ohLCyw0gAw7iUg848YSzSfdnyYh8CWN8IBho
iXxKoT/xWQxfJ+zyMXK5o8IgQ5T5Agsy6C9izxaP4vHWDOBDiLEnbe9eAQAQSXNR
jlhnyhUU5QVkwOryJdSsxYl7IaGA+KfIR53nVuXZ2uAgz2eQNTZiCtgKEHb6pnOz
uZZdrHnxXYnlLqd8mRZtGWppGCbhptKDniOSAunVS0zvWpobXMRE5wOuPMVjsBrK
YLaKuBUxAwEemXdGIIeSH0toq4jhhrRKlJMXYAHp+OjJP7AVvvo/xTqHfKUJXJxv
woSAfLjhHkeeYf629wD/4fOPMao9dkxgk3CHjjiSd+qIs829esjdazRvJ2YSc9QF
UHxoq4vZSy0YCdd4sj5Q1w49Zdbn7jMzqbK1JlucKOwmn/jJwx1VtNHxWRm6A/H8
XOMMarqDZ9w10zzesoxge0PGfldoWmkSpJXY/C6LX3sT9QBZdlpuQ8cUkdHCtCX3
Yyz5p9F0bf7tCqfHs1BLvUEZLcby9DfsetJ9gdYZk5FETL5ZPaEOJ4YSHILjIg9C
/Trto4qQ4J0M/h3NvErP2SyC4evnwU6BsRz+ZUS378COwXoOiwJoCvh3lwl5VEY3
YRtlyYi5QwrVVFXHC9Egc87gF4UdWm6yPnkIVCdYLrvdLshTktUR8suLkUP6sb+7
HHbRVkahh0SWUIPrDuDi3uIw8e6Yc0ZZEV/YBJkB6SSjp9cSA09PsULQy44BOfr5
H3LyEh4pPnQDKThCiSNiaw7hIb76Zp6toyeNdvCg3mrca4sTk3dWrLaCTI0jnwUP
O3mnIEzVF5CYpHGOhqHcQPqH2Lu77vDsUdylX95xHPyj3ZbIeOUkthGMS0WIRPic
/MwfM8IFYIiccL0gw7RVsskZRfh4MTmKYT7rGFRYxoZt75fSvFRzUqp3+eoNmptb
g/uSJ0jZwqq3r416rWtDus9gzMDeCuuPpFXCNRMm4KS9J6mHuFMMVU3e4EsEgPzz
r+YQGDPLf/oHDk1lQoVLOm6ynW/auB7lX8wN7LxpVLawZGEe8C24W/if+MF4h05G
avy2olxPmcNRS4iawyCZCcJDIsaSAW97sJyKiF8JcbojZUECd8R0gO6ak1srdx98
fEcvQdsTXylIYqWkvr0+X6lh8repQcWpNHLDflTJM9gzZoetRBRhZxNxR/brWYwA
1rlzy6TeoW0ZzGB1dizyUdnfMflOCMtniZvIsS6/I6wi/fYpLOtMDZGF9t0tSiSj
p0rCI+dT06cBeZNEjhlR2h5NJfRQkGyqmgPk0KNIuD1YrPuOmWCqePI8AD/b+0Cb
rqA2TwYB8p9jXjJpG8oaxgoFuN6zMhRhXnsMd0wJamnpKsA6ygOGvT8Ch+EQULel
AzTsptNuOkEkEeVIrVkKkFysgUp3UQwBz/qTAcZazfj902b/xJwdTrb+fCG0or16
CQORoyyvsU3/8RJppi9fJ/LUjvQACiYQplYJAJKSWmu2lVzLcSW0If3DyivNGYoE
v/xn/zDcikWfy9zM+n0V8eW2lwtslik79ni/6AqiL89Ip4GSFBQl1Swo7O+zN7on
ze+PS1lI+OBrm7n7FgBgsxEvo2rQFo5Jah66wwRQv4JQVlTH8PY7sKYntNmq6qp4
HXiY3xInHWQaR73ciatxmnGtndgMNmQmJKxkPYxhS4rEkeqAGSsY5PS0Y9rsnul9
bpn6sNesJIH1tq/RCT1toazQLADxICSpr6PDEBf9bQo++XX1W8taHarlPKjXkPil
LgqVolBplEFwpM7bo1h3Y8fAttxfvDvi6YOy+pGRKlwuqihO5YF/+R5OGCDInXtY
W95hXCRrX3ehjskOC3eoQ+QHtSl23nQPjCyRb9gTFQIQfQSzYQyRDAoDAfsOJEEs
d+kZZ+gHCzpDzkdwSSMd0sCYSwgcf/97wSQ1wmi6crRSrAR7KvbClV0TBOg7dvn9
cZo/KbJ1epzlzlV7WG/ThQYvV2ZWLnORq2sIy/j6K/QTH7y/Uw/TTG/1KnSaDqhm
oTuUhTfise7C6iXOgFIHg+RgeTwVkZ6oa5kVbH6f8n9fG8JvCprH4IpuzeHLzQRv
dJ1M9/wLEhEuNdJFEPldpQBUt2XZ8SEES5nZy02STgQn8HVyrnAB5O+PUn6APjMF
D52l3lHNLaqQwav+lChHodwEWMhzCDiGHWMo78tSnem1wQDXrzUbwbNCw0uXgAkH
bWiKbj0WM5Wddro31WAEtPqgerePAhy/MIC+VMuUjABcXKM0ZHdyvFOoM17p98ei
a/61n2pXm1pvNWXc5JqhHseFixAT703XR5lRt8kMLpZw/Kl0uQq1bLTPR7X3oAJz
XuM1ioSQ6xB/whB4Vb42vHTVM+bHHHQF0bxHdsAw6uzKlcbut0LCX/rhHRou0ead
XzqgnbTQ+Ul8KDFRnLVAMm/09Fx7Koh6kKyjHUObidY2VY3p9vzWC4DI7jyGwSdf
15I6+GByKa3/ia4ZRVUAC+gwM2CFvH6a9oP8ibQopyABfOhmW75ZcOs4OJ3nEVAl
O2giIx2LZ4Z1X2pQXqXYakTX7G4+rH8Gj+82hvRoQNxm+uobqdN/QS7k0gV+vHM3
WpB4tdEfT02Fvo0M+mNMAXMpcv3YVpkm/LMNh+ru9YZwEIJqE1gKOPuhbvuWVUWT
7nuw3XwMUmq2WwsEjzh8gbWHdKYdZQbSYx41lT9D4OH/pznqIYFHm3KqYO0Zg/Wt
Ky10+11pxR2pLY0fpxqKkeMsjqXZOYz4GTwq6ZYzrmTu3j4EIiU9pEcALDRPAPOr
jcybOJ5uRSCiv1rcY1iOgn5YKw6svINUzX7MXHHSVxd+0Ebd54522r5xMRYgOHOE
MNsDekrppTo20U3/Ukk38fiPqSNcgaRxeGJjiGIulVb/0BKsZ8HeCQ3CBpm5rLhj
yg99aUbUw3gGu+luVpCu77IFD7eo9VPWTO2kaWcJUL9GE/WjTRjvba5tKjC1y9zo
i0EhFKPdS4tZKWPz46a7CgGsQHKP9r140i7q8UFti+2oupDcsmsXuSTToMVlJHZw
LseEEVYkxWXOCp+D1E93JGhpB+GPHNAfr2ja4M7cJncii6c1Cr1ZmGRxyU3ymkK5
Hs0BDp/hnJya6azL8yffqW/V8PBEsGIvbDYGTvOUSIbJ978xnUM0K7u+dCPMkG8D
Ba5XmCziYV00xCxPje0lXL0yrWKaU+8fezmDCs1eQECkVaIw+YbbnzRvKmjD+8pQ
TljK+9wtyqhhFCAGsLBmLsNmDKZeUigGOb6nUyvYq0eyWo2JRXI2fbkw9FX4gZJ9
bU2pSNDarG+riCkKOpPuk44JxGodsqJOq7pOe+KPZrGEjEjzl47VouEEmEu9Iizk
HH1UgxCvbraUdCE3vaq4Tq6P61iytrvozrt8uJV1P0152AJpjjeWkZgrAWUauIlV
eF3Qvqu0p9dU66LPZZXoB8nt4RvplTKyDidZMel3iHheT++5h9nULHRmYPp86ktN
Ykgzplt/pwAfoyIHGTGKWEgb19OpPgwa3NPfi3badKMvVQAvXdC7kSaaJIQoPMvd
BPKR0bkRL8X3evA4QSH7S80ytrbKQIg/kMz/JdLiG8smKY41k13PXKo2sha4r7yr
WpAQddsGMnhrPrsZQHf3DUmWSDp0Wjg0VzRoZKQ89qmO8ErCpbh3/vxkcIlenqR3
zb4GfwoNH98zs5s1sFG2z7QcEZSWanuW5vg4kdoZ3KivM8SxuZ8bZRlm+D4LctKe
wuFJrDv/TaZQ4uIHM45ZK+lvAqzdezPGnILHzqj7aZpqenfsEa8/oYTJ0cELM60l
PsQfFuFcTN9rCN2VyHJC6SYbxTp9C9ZTWsmCBSDxXI3ikn4hPOS3Bs3fOGatWzxi
pBUiSmcUpZSNIKZf4rqwaPbQm/KpnA8SO+3wBgMcC8u3WU69dvQHqzcWyvg4KUcF
ZAV0KEeOBqrQC43RB/aj5A7SWz47EA0dz7vSOiLqhPYmZ6V1kSXynukThBVwSvqr
fCXW+ImuLfURys0NNcQsu/g5aDff8QZB8P/ak1EMtsvIHvPOxaZl2DQuWASJVfxe
OmHoBDsrVPfRotiQ9wpDGNv+UY9FBIQHlrrKlsSiEWrJDAEzsrXiCSqrz2n/+TlD
4kQHTGMVD/vcYSZPi5eelci7ABCq7Le/rsSRmW0NXZwQhzkyd0c74c1HzGHSQv9m
vW2XBSmdPlz+wzYe+Oq812dCnMc1HIQiL9pqXuhAIPHDiQXm3O+k7K5Shf40huOV
AxqqalMfE/cDO0y3KZ6JoQl/7TBM97OhIM+3LmIf6oIZr6xjId5NZ5h9ytBOmrI/
iCprbNUFFcpxPKZD/F9RUvgGGHwX3zEXnHoihikPFQZ74Pad6HZkeiQlowpnmFp1
zZQRgebP2OXqlu9o+QtjzpnwwfIPmO+IHo+pwg5mlAq2M3NP/0MY8bYjZRn2K+PE
/TbdzEniThO+7l3xQ55VSyPi5eLRqfbASzgHhlnvzsaPbiVFoXG9O3TW09YXEix4
obYuZisO0JTPGT0Wb0kUEhqOVQz6+k1bPtHrsY3VpfPDMAGjM9HqesHvZUIPN85J
I8RjLLjfy6q0wKCtYGB/PYWQb0Fg/EJif68RuxS8nmrT9yosGmVCk+iLIeBxIq1F
dNUhXgkfWRU+PlAbUEDuB4x1kAAyz41ljSqW5Aeja2tbwUZ39rLIJBu9hT2Hd0Hu
07ZvNzif+af7YESVTRZIMn+fNbE/qeRDgsAbxm7ESSZ5ly4yOpHzeMxJVqj0HL3E
ZY7LJhfn7Hep0xG7lQpFuDf67o6u/zYqP22alGyCzLR6xvjhdr8cJH+3409LoObt
zv4b43Ot9g7b0qFqyXaJEKNAAfrrHzBxZSNWFzH/jteIVfQ2+U2E0nJFOdJPaJHe
JtmaMpVVg7Evp+p4560bJhY3aD0AilWlLz/aH2/0Ji4J25ue2o/oGGwsPx5thTh8
ySlObjMkaQGC8rPvpU0n3df3nEzsrhB+d507BqbE8C0nLblgCTdZwlAXxiHQHpAg
GZjQnPRhqO0IIxUjppkZ07yv2LhYobMrj1AjENo++lm2fgUanL2aeH5ryyVuSP1j
wUOqxXwB89SVwIv9TTnGR6kWZ70UrTbpoJjXmh5Z5D3ZJ+hiwQEs/F2arshtzXot
3TAtyjVRyhhQ4XTv137D8qTLxLGZPo/cHIQEFSsu/P8v/V6cxAQWrKmJGrR7IEqs
1egTRr7FZKYUMXlE34WeTqKrEZ+ecYXntReXa8TUcFeztZc6DOXr3rQV+QX/xHk4
g6GoHrcK/N8fz2RLYAorEEog5RrDkn80VqpqtkS2lQWmmOa+u1jdGj39/E2XGq9d
qRsViotuRNz4WPK8VJCc0EcnAo/f7bH3DDdkv0oYdU1yVgWxJNXtYgaUHnn9Iqm/
DTLpqjq1QC2Re51Q+pmhAtb69WxbeeDry+/Bko/Cquv1yfceQ/SnblmIPIZspR6q
DXXxUfohwiVItPWlXiR79hYhj2ca1TuDTfTwS9xAjVzLuGyQOmDqYsILT3/4Lqrg
9m2PfrdMpSAoXOareu3ld8OTDIYjL0vdaxmpUosRgCSl+jtMo4gFIOc+jzCas6q6
Ft5hEuq1dcus6LRrYtRBA88GD3FfAJYk6qGnPizG/AMYPVGHtrkt/hR7j0tS2dCd
fWzRVUv/JkIC/xMQVW6pRDWruW+sRLITy8xgLE5L92WERtF0/kAeDLrPbH8lJ9SK
kVj5LxMtGb5m9KKJINfUJUIGydeMPHJfry4T+IByGvXhKZY43ry5a9ihtSnav7rs
dGsrnqQV14SLhsNi0+EWgt2xwRe3vDYhENIbcQz3cthcUFXhaRXwQYVo3w+WvHjs
AwCxtQPxHxxBd1o/vvdDRwrKp0t2yrCguLkhXDrfJ2qm9gxtZY/3ubamr7z2PSo3
YKZubUH4QJlBPzYHn5OJwzHkmFqEngQy3Yt7DYtSBkDWHMH1ew+YqQsfRFLWvM0+
MUY3GH3xJu2Z89W2pfhw2p0jaltpg1w65KySISFSD7Sc4ARVKY5u4doMVgwzwZrp
ucqXIHUyQvuawIO4wtxmQHP9sFIJ/xvHIJDByTunLCZitlm25O1qeTMyKhctaw0A
AH8uK2Nh0cMJCvU8GAtxu/g4ttpFHpTvLlTlZweDAw1xXZVJxqhgaNZLlf7A+MPS
Nh5v/+GUQy7e6SGwcqDrT8yNSjPY+sapELxjwIFoL7AkkCdLrRAuuzAq+RXMj8VI
FBtTd3d/YCGIVVB/T07f9or0HsdSfkEW9pEW278WA7PaAHzDDGj6pGIuYjpxKB8L
O1QQYAjnsGI4ttd+6oeBd4n8njaCsl/SJc6JliF+ChrWuq8HGTv23TaLYvNYba0t
m0rNkpd27sPa5K29eRt+Nk2vH08oO+QhDseI37ktKNimUdTN0PEe0Fs0ofNc7Kkp
WCcksJ9Lm+Qnq3Prujqkj3WVkLHmahbHCM51+nHZtN4SFb+5KE9ZvzWRBEy5Whpz
Rn4F1Pfu1m7D5TyMX/RrU2vq/f7KdqLKuH5YXMmsCeIN4U8Wy7ewYXk26AIKuCsT
d29vzoWyDU966D41shRxv0PkTFvwSl0MwfBn7nUYYge8ssFICoOun/nTPM8bW1+4
GxC2jHbmGK/Mzces5KbPJOzbcpRMug5xdL/F22KZFKTdSf72faKbG7lOnZEmFjfm
zAxb08rXzXg8mOCluaIjil0RhZwe29a8ofywybUYL+7b1kpraI73CIxYVGcsC71R
OWDC6iTrlgboD5+g3N4w+/mCSor9pKBmP/L2xry/abqPf+u214oTReov2W7Ax4mf
EcKLhHG5W2/TYczXr28KI8yQ6SVVkLauLRI98xeiI4VnOtUNROTO1iyh5xXuWMy8
dfs3P4FFS6aXxb4dXaSBa1oidju18U4WwXKExg8qfNk8UzIMA0yBOYJd7EmuqUVr
VaxCO5NLZmtq9wByZH980AaT9PCuzoeGOi9fhKPOPOPLsmfJAqPefqegdN1ohFao
SBGPI0SedEBedmIhPOOVrd7n3rYYGYANEd7WN7R73hHTIIFZjuIt8BQpOnyqra9W
6QPvvNM+h3W0TnBtHW5ehEET+GH+7eH6ZF04MKv//jCSaKSWWU1ODNmIdV+zxVw+
tT8RrjkEcAYnYHAP4Mp+dowhRnf01nMQY+JKC1YEaKfBZUWOy0fy5c2pEIgOlHzk
iaVxtupVxePNZKRJbA5J+g2j9u+bEBytaa0J0rYo0EszEt60xzglCWyTGSjnaqO+
sqb/ECRRl/S1zW4oWeK1CbDIBBQWl2KrGKzg/Ee1GR9ttB7TWntsibErquUEQNEL
hb2ABD1G6w9GCDjhaUAsqsV1yYoVgo4CYiEvMBOYPkbveDjvzyNcKU6M8mvZoThE
F0Ks3FqVgK0I7EXwi1xG7OdQ3hEIdntYcHycaY2vUURGSO/C/bkVR86cxet/tsr/
KZquR50nIGXxMWXEqdwFybd1Fm1sHhV/Aw7Oux3xxa3WjGTLcWhZ47Kilh9dc07O
z3OkdeLAfasJrV9g5gR+ZzrAB6BLHarS9I9kY1IoHHu2jS6XCjJuQeHxe6/wyUuh
f4jwe7sZhZYS06ExSVJjwIhgeTq2n3EMFaNxt+Wh7xFRG6i4ndb/QJxx903nFxco
LjuPWguockNbblaU1K895hOlr9X4RLjn8ORaL0TShcXqkqoMlIQbWXV/07EYl4B1
hN54J4bknTcdNCz3uyf6ptPdrwuJeNJ8Q5d3jvAqlpQeMMzZUiRuwt2Vg5YlMq1a
wi2sFDX2rYUgVinVDNjUt2xsvRjcQUgdIOuSgycNS3ugMuI9Rqwa/Xe6s5niKh5Z
MMutGMqUkHbIo/yAb5wE6+yOPryxX8bl759m+Th2nfAv+ZbMKEXWhcXjWxeeYHLK
sgmWleJt8GzFea6WM2/0zsajpvyy88Oxlf58ckpMOokNXCosQtQedvHIgG8SOotD
rPVV5NOf2/4sx/7M33Wr48Dj4S/KUJAaW+3j+EgfhZhPBVA9BkD8i3rDVdWaSuQ9
EFmCbyQ3BR1ojDbY/lHwW81GxtsrPTp8K3K6Ku2gYFu6XmIETz2maYmjbWKKLs4G
zEFHLb9p74Lz0waJ2vPaBVB5ierjBgrWccp91Vh0vrmLS5pOW2nrVHVR43uCzaww
CQRbWshUeI66tUIXOjUymVx5Z1A4qh+HTuKLwlm1GgimWdkdqoS5ay6I2tOABzz2
Xz8ctj/kTbpKCGT+xUfkHh99tSzzySmgRcTOuPhcVIMXe8AoBFixTigT/CBOOSG8
dVjOQS0G9NX5+lRbkbKK/1c1yJW39BMH7+SKlnQLlQy3EOcWnJL2bivfk45lRbMk
sUDi7pyueuuHURG0FBXNxNuSWFNabDxFJ754eAs65hTdb/pBDJLN3xB9+kt893VD
IKJWoUpjH7aoyW7kVpIN9aYza3IJcEWIZdw6p2BQuWfV+Qwaq4JC06UWBErmiU0I
OhqNFajHwUOmLKAMSxo2GBKCHCGBoyMEzTORMjJillyONjR5uPfwZmxww722Ccae
Xiw0jYQJ8shJTgzYuj2ud0vU7NaTe6u0hv5rPtW2icBj5tg5Msk3L+veKTJxr13Y
jPDC789rziADCBcfmrdPrISahXPKxp6dddPnRsNwsWTH5e0ctI9WhXT+i73okvbl
v8+u0dlieERFUndFbENn9av5ZzZwBe23QMMO46HmPzakDs/52b6xyP7RtmxNY3ys
icqMYHe8MQTNhE5/JTnw8hv7M2ju7URUirt5cVecT+FgHFIO44yDkm8AhoAcw0AC
eKaC2FMwLGO29tsepLlEPuSWY/YeRWgVjXieOnevM2HLc5ot5sKmGAZQD9NHGu6J
zi2BSjj2kZppR6kP4XLVi0kbplxS/IA1IjcOsSSPEEYH9CzdDqKRokkvcoli1dkj
B7tArnjdkOADBGQAS4yBPS4eqEFZdoDerYqhHKjwQV91LXYqhmb/5ulQKcHuAwpc
eRzPOT2Di5iLVnlhAP1RlmIjxRsOgIW4R5C2ZDbKazpzitunm7UbT5jZDn+jblUK
8JOyOKD/GdlwbW6doTozizwZva0bVBBxdltWalZD2ZnPKdYeKPZkOLcvKA6DEE7Y
j3utPvZ9qLjP/mQwZ2b+rAN91swEoBsWcrW11n5Ok+Uv8BOv3XTJOjt5RwyhU55o
tq36pZAD2Ne7T1NRaBXmGmE/0+dmBEnNodrMr9mpS6lc2TvYO/ke1M5lCjXwaT6x
qWGfQfbLRpyTnnyxQgBbLwUodnj0vOlStsyPzS7SI5Vmf4lEbKzFf9pG1IFgEBjP
Ssj6N+rLlnjzcqJCfbq1Ao7koWVBDA+XN21BZMhuEMzpxB11XArn8zyP+yns86Oy
HPFheLKFLhDC9J3B89qThn8+EM0+efIfkD6Jou2iC7waQi5xGGfheQc8WIEeVFSW
bZcaFET9G9+Xy1jK50SV+MeLAjX7NjKtcVNL3pS6vxemawfm8R4GHrS/kPSNx1H+
kdRnpys1gc2rGWi71jZjLx+1vzLexJZ+iApgnGcL9vA54L5FFNzc8m+ovirCaIP0
pwEZC0YxRYo1PcITu3p9ipR6OG1yeFE3eZi61jkE1UwJ4xNnpogkUKXcrIMAGYRN
D65JyLXWIkTKpRxVmuYMF7bLO6BCPMFGwCrnLy7kvDh73+LxvJd4tVtMtRroiOyU
Sgg6zdn+5lHxmxfxotZ1KJpCZCLqVKU66IWNHPZGdKrc5CKZ/4rvQe0Hr+KDL6Ls
vN8mfsUz0GqgQoU9mbabbvIDItQabLo4ZxkcACNY5Q3wnM8UoqPrdoRojyHqyBp5
7aSVkP+BzxyKpT0QV00DKSK2xhcFfBXEugHZDvEgN4wTyo/7qyYgO7WzsqbaNTRG
N33om/eBWGFrqhNUb/mGtPlDozAkHcYLvfExm5i6Rd/XnL+EZnowh90jCLAy+byH
ObmMvthU6sYOFV4soqLHPUWxlRMDSt+cOQlsCI9Ii4FUNpFJuWyemj4v8tG3hOd3
sipWYfpBUW0RsePIFjgXXQ5RJm4rcAYLrHj1JjdDRFwm4uEJJcHNFrtt1vULmnVh
Qv6soYI0GEFhulezVm+yLE2Z9tf/eT5vre3devkEZFcEwm7HtOL+5vR1ANuMmO9u
+MkTOKSdH9zPo38q4LB8zXXz5uo45WRAQQW+nVRTgRDWJ4Ej9yVBP6IeEmCut5iU
z1N/t48owOE+2xm/X7jOTBg9g6xgLuJVW4q8vkclOkmg1poRC7EXLE2tbWYsd7nf
W2dOKXoHzLWVkPbasGYiLAYBUxFC176fgEJn7wngub7XTFXcvMPkvXRDeDl9zfIK
cLNJbHB+SMz6q9y/gxKLfMmHJwz9RlC5JNAsoGZ1isp1fjCNZw5sxx1Wi0TISsai
faUnwqIPzxaoci80teuFanXytEmiSd1/djlC0ka0jGkaKIYNGBUbbvdfmrDiOaa/
M6Lc9Ro6YOD4W9oi2qyiU2+ucgZMbQwBcogLhs3RLjgrNd/eqUVina+bc6exq1rT
+Z4CUCB6qK6YYTZhj8yrjcwHJoQAfjFN/822Cnsd4Mwo1uEDQKz5Fkfatn4IeUDO
1KgkpJr+yc1JuGjkxD2mJA5WiV/hxWo3YLbLywNR7BCIJVx3r+kGn+bQwamF0DaB
u3YrXJgH7VagXDBFX6/IWa483v9MwIjdvLpPhmWk3g6+kgYi9xHGxVldqrO2+9Ba
h744JpQDWW5QiLo0Q7wvT7ZcV3xNkQ9BsyxgT2kDguxM57Cfe30m0D+gXEH+CUW+
rt4ZQBx1QKd1/XTsvUMxK0QRvJM7bPr82S8lqm5oNGvEhWdZzsF/JQ15eegW3r4r
yeYtI1Drc/Xo8iYUrpBsLE/CabaZJd8E4F7q0nkortFw9hEQBCedBCQJG7i6iRHm
ZWBwIx/M+4LbJfoB+qLPag2I1OHL1iEuIw2Lg8mt+2IZ4q1QAplbDTWaNk+jS7YS
3EQohlL+YTJDsgoKEE/UQCRVaCSlORhCDrTtdxb+bknzCljrAjP36tlagTj9PgkV
X1Fa3W474Tmfs09spV/0QQrbQ2PGOqEG9L5iBxErFHgPGrJty69rRvFWjRGIhyDT
AHfqKb0daq/8Kow1K9A5MtNmdMSJkmEPUWDOm96HJ/KD3ERnkhtjZMJXa7e3fhaA
ognrz6c6hTWdOL6OVO8h9uO/iHK5hnJmqdPiV85R8LmM6ILIXkOmuGKNcSzYp0ad
uyQE9mKJNFGF7UAxSXXFR1fS4c2NUfkqqMutti1HbuGwhay10JOhWTVkwY8xx0tl
k+HxYtau1rLzI5JX2Bqa0gxC1Vw3G/ehsTa7GI78iSeHBvLqnDN8RA1gh9zAbBvj
noiDkzcp1chMc08c1VAmDqr8ZElwkBoB2EWP8rIFRWwTNRE5LEOVHA/yCqCaATTx
jJNcEpDijXv8Y6joJwUo8eSq1GJUeK2VALubeQ42EI0tF7EvQfgX5fec0jTmEtBj
nygn0sRs/wfwgSjN6zXEPAIMHLsNiZyjStb0oX0k8oBZiAxX6rYUS9gUnikILHuk
cmP44MTWyAcZq/bFhMbhOdRYxnrhtGtp7d9giTpoiXzueax94fq6N0X5oYiyPkSZ
ejajJ8YBjzrN98ict+V2HRm1TpyvPeHXFoRSIVuC9K7JB4swHNvqIqbyul5/FUAk
9NfVuIDiTAIux5y2SXN1dRgxyu1thGzu4gW8RCUGCpIG/UXMz8YIK+4JxRS9jZaX
G3VYM1b3w9VfIbnXeIPYbZtQlq0I7YvjdU/tHl/fEP0Dqp8zvFGqqmCNkogd9bKd
CBwYSiSowHgoGVmMfKyTgJu9D2C1p56uBzBcs591veNnxT5XZ16yuRDgjmulBo2J
mMLLoMaX6v5RTyewmXxZyWYQr/L6G3Bl9+eevGXbtEtZehoylfalrbVeWkyoRAtx
5ImM+skGU6yUN6rxXu6t3PvhfMXxlmJ1l8KmBr281qLKreHoxAo8/jGxlXUfVi0n
CjwtE+gKoW8MXsGvQxNbGrXESgeWdLk6v+FZItHXMGGcOjX7vjXlsjsJUCsh4My2
w511Nxg0KTf/fdmklcAbjjOAWoaVcDCSKlWQjBl0stFKmtsDjskJsV2/HaJa6APE
eTxKqJvxlgb8UxwuvphN411nubiBX3R5jeL5WR3ByCrdq/O8/IbyT/367kOPEC6l
jNa3K4GUGkEVG8wXfXubqrArZzOSR87pjJGOenAxAcLaJ0E42pppotHmzIFFsBnW
McNGMPQ6SPf4uN237r+qovXgKEVTUxidaZuc8PpUZ+IxaFcWcnxJrS1u5iDNTVZx
in3nLRHx117DRED+aeDobLONRBDEr+nv5tJRmKcAVrvEH80tXwxQPe1CGDmqiwWb
Nh1jCSIJR7pWbd86QZT5IWSjluAf9ZbRWZVsfNtj3WHya0KuP1Ph2N/cDBwIw8kD
0pSVyA7rkJAbPaVZ8FOzQNINOKAjEkZiEqe5jca8OeKIvM5YcHVJZkPdUBVTEFh6
MW1ZtcSdxHrCcewOI8+q3prsKyH5dFv/btEnfIm3S9CaRbxgkA2vylhNMigVYU7w
HQIO8TQHgWKPXIuHdJDlBARaSNese6pLBwIboetdCHM6OSKaM/bQsOBzhNw5f7nt
rYILzJJY4RX6sV8rJqhEnEUQN2GY7rRqqSm08q4sHJ7BqHbCZaSkapi7JuM+6RAx
QODYE05xOGKtvHM5dryf8+wQeEjA3YpJrFJ3bLB/dgQBiKrHizGWr8NC9TmazI8u
ZiCoUfASLMsQcYf2hy3UinC/q8sEgJohGc+CNogsecaZ4x5NK4Z///s6qppAK404
T31fQfeN97dDdwLfjXURrElb48sGsAdoz7XblQfr1FJjxb4tG+crjIRwV+X3Ju0o
kW/IBesYJa0vhTbqgoY+rcG2vdzLAhpKXT8nunRxBH6/4nA5LI/l2w5akvOlDmY9
kMLRpShgvbXm7dRjqaool+ZQK0uupTG6JddFMD2zcdKiOoVKpuF7KZsMEYS3iG9e
5DnCqx5vK+aeYOXhWrOuHS320uLmc+Om2XJOveD8kTjOD0pg1PkihEVCohPojT7g
ZlkjpduyM1QYaXpp+3/wKjTRhRX5IuT6RmE3JygJP+/9Ozg6yQP9KFymu44j86/a
td2Nb5N8rJch9gWIzTJfdeUgw4zA9yCpKFNZEuOOLe4t8ghIkIe5DoQHOgUMdl4p
AdKjak5ziZw3jM3ApLIQ0etebBeprVTSUtdCocFHo388ObUZWPB+DZlRqP1gQRdL
62hEeB9hq52FFFU8RTPGurKz4Cd8DczK3f7FBtYXz8HL9cHZMVniWD2r4dPWHWE2
F/Z783pelaN/CTo+DhE2Ae/1EAzP/vXkxehc6V9HqTa8VcJkEaMHsj4g39mNrH1N
nlsDZj8xhEQt4je0p/t3cv208n+nWQFAJaTOGkQLeI2A4MjQuZGre4gT7oNe+yiS
P3wHdqZV0J0fWVa1cEiJaxQOWuPsTJIRX3NisFa4y/l6MQC+yuZyDKr/K+fAj76u
jaW9yVuxXp3Yso0EK486ixdIw5R0RcUCSX93+r+gpFSWnzI6yJAhMJUtiIteNezO
nZVmxCVi1Oc3k54reLMaIvqlDRNM5EI4rmJUJ0kDKaJEprwzc7kQtdFRQfKSh+PL
lB4O+Q98oEzEOGduBkraOcdz+hOxPORYdzkTj1pVNG4TVdO/2D316O5Ah/7Kp3QQ
c6PfdUcIAOhzLrpcaWWqHD9uXt82YLSiI6i/b3ofcK7uIRpH+ZojwvSUwoma1VHL
1S5G/HjMjHzerfILpyUUJg3iJmgft/Aw2bH25JC+Sou3TyCDA7knzoatI2l382m2
84nWe1Gg0ZkmxveCNO+4NYCVn1WSuDnea9ft428LiCubSQ+5+ALxssYzMD6TUHaK
zU4M3qQSzmYrAoHWnNSmynv30SEi87+k5uin0dmHtLWtOcdBjx3ZzWsH4x5x06GX
5ZBjINvy32sQGUBEkkDRLANNlau8zi3sbT04UlWS873Dkxiq3z81FN7KoQWeF0yi
yG4t1eN9+nFUVQZrzDUdKWQonVQe96gaMQXRMmgr+nZXaDCy0O00FkwaCkJKrQQj
tTzvZgCwtA2nJRA9mR/tY+bBXui7CtEYv3Vf/+UyFZRJktZ1wVffZA9MMOALimfd
wReZJOqAHVDJAAbKn2Jn/1J6Ymbw89DbezIboix/sKB2lM6b0OuHj+5d/C2k/6L6
RuShwXs8pV/PLEToaDHCHETZJ0sUL6Wpqsly++Ml9zNQ3GYBqAUIw5iVjJdAr3fA
J/H2wMFxxVAM0YXTNiVEmiOWDdhrUKW2OeMdEshbHDNoGIfODIPXVtKwhz13CIBZ
D6Y5JP4ZrMmhqO8QmA6QIhAO3kzu9Q6No2e8hlFZ2k4p4xiH+RX4TPdqkCtpA1UT
U7rWhKNtSG1gFDmZtM3gBXbs3v5qRaPgE5XrL32IUgKdli9GE5boxQYEfvtwtel+
SvtFUCPXmwr15VkBrSVO91OvT1/Yuwp8XPrUbxvPj6JlXhMUWQn2HmKD2KDgcLTp
XhEm2EgUseT1gfT6hHETzMitQok8eQqvZCVSZiRSbxcORC8hKaG9ca2C2nnKbmjE
k2PAL+V9/yTYfS8HNDJRdOUSIepMrBes62Hy8SUt3tTY9K5hKYP+ETtONl6s6rhj
Zbui+312NwfKZ/nQjU8YQKaiw1nknRgMAHiwkMaeQvGEyAc66FmtMXSWtFvyLxVc
bA/heekTXZmtEEmTwnSWK8b5+x9CyPx/xVcFCjim3cSeBFm3XAFuTTUA4j8w5hHm
+Y9nY3rRm7qfeMGmIK9iYZ+q/Ot5FwCOkEilK1nBfbi28lK270kY1Tsxy8g5YfB6
7geeulpyiXmtX1ma+Xq7v2n+vRfCverT/S4hIkq7NHwxNULy9tOSrfZq05E6X1ch
YxWCByO6mQWTBgmliiVFt33z80MceD0FoVgOcRZYaa1Ed4OVcwgswgrfrSmmqAhB
/VFDOg7qXGKiCgJaqHVgn5FiwlBfaWWI4NFk7z/grMjRvaHGoYaQvVtFvo8/Gp9+
jQG6wj7OVlVPa6pjvwm+5DpYaBFPj/YtcOn9OfYAksPy3M7FEg6bghECQadHpWkN
99P7IJq58nqMuXGG1TP3xvn+W6cqq81VISqk2qioG8X9iqxPoi8CspEZuIUm4yPK
AG6h/xNjTvMVo8+T0pKN+XxeAWKfY25cS27EYw7hYEUoPSUaEdBJCHx7Z4xZrzhN
Yp+aGK24/wt3m9TovUYATSYERhVd2bpa0EUPDbsF65UDGTOiLbO1ymuV1CrBxgxn
dBS/1VKDZtyBXFIeVkUgwLjw1zKUFpfWHLLgjArtm9tEpyVtUn5hFeVI/tnoJFuR
jC0hQCbBmDc08dGDUvnbauSX43aUUtwtzlkEby73W/LJeQg0N93h7y16culmf1rI
0m1SrROhDlpAmpMOw1T0NeA0IkZebtjlOPBfqFJnCRNqKSE9aGFAEh2/YQCtwk23
xVAvGC0iFd6cLOFXnCNh/6q7u3brgV/E4oXqS2fb9LU/XTa3+gQmhlqPHbBgLB0c
FhpDvmzAWJn8ArsUhMw5GrI9TDwMOjn7gIKAnShu/Aqte3wvQll/WF79gIJgZfNG
YO4+QXd9pyMwlIUmb8Ak1B2fhSxyOL2LlyHNJvWcG9CJ3y2VTI+ljHDLkjWVg0PB
fzi3I7+syiHeBW18DhCyKgRgb1Xiim5VkUkn6ZB4mGb9igssIk/3j7nWsW/v/aLb
G5kFfxxwsnnpzCHnahOj9J3z29GIHRiaiEN59olERwkCWcDiZz0gqm3HpelkvajA
tjSscm1SxXYLaBD1ly6y70t7sA/PUsz9Qe+DmjEiIFsoWm1Q1zT2Sta9nuPYPkG9
4HzUpZfEtXIolHcCumDfwHBSVGDNQ0YsqGshbVlHJFXLSokk7y03kVQym8xY27kM
9L/9TlxyE0pxa9atrXvxxWeyRzAv0jQCnhIjzf6e5/4QaIeyfHzR8gD1uXs25fe1
rjO9tmFUNXfoBnVbzF/wF3pX+H0Ctc2X59MRx5Ckh8+9KAHbrgDeyvrMXK2UOMsS
BN9IV6c89ob6hIEj+K+pP9DjUzWhE9r8eykd4opv5EVhy3nlCMsEgWaSfGGO0pMi
kIfdHZI0kc3ZKUU5JVIHgGJRVqFkg7MwUvHnajDrfAD4z4/+ywvguapURSmacxfV
scH/gr8sdQPuFUJJ6llSO9zToZgB3f7wyGrij6Lb/Hu+EE2194agdSLxUV5lL7QE
Iyb/1khUUSpR/DNzNWC0Q5gpmxC7ox6rCTwgXRNhPCWTW2z/h+l0XV4sdmVSLjLk
XtxstYH39UdliFzWzzZTiX6kQZkTeq0qym89GVSmn2Toy/Ygc8S+NQlt426nv80T
mjJRR5H0rXZjAl1P97gQ+y3e1XR/sE9QKR5SVXD67Y3/nFVTUZm87aTG/Xn1QH2+
3+csfo+gvJE7NXyf/bMtcx1B4cz29WxSg1BcG5GnVgAZEmxwE3SYh/rpzJMbyUuE
vj/Pax2KE5N3M6YCfV0tu+WVtm8ucAFJQEri1ntgqrg3Smt31rSGIi6POBMQxjqC
DlPMJv2A+qVSOOfQaF7C7U0EUCZ/ni14E4kOa2NtAbzpKr6nu0yp8f48k0u3Fjps
6UxcC5KkxRKvQn8p2YhHk89zBotqz3V4gV+Dd9tohVkuBRJFaA+ZKOqGg+9Sjx5L
z47qIrker+gkoc4FNkT+LsJYT7xRbRIzG7UyIn0htCvV1b2a1Rkt4IG1i1oXJcpj
AQI5vkEc/pfYlNKJ1GixfN14FgPfZVX2/eGmjCz00D+IoZTiRW8txvsI7tM9K1pE
ZlT+51XGHqbXsMvkUTyAZjGb8jLp5IzRq2PvThm3kDf+xO470YLNwbHA49Sup1EC
R+Nh5xJH44BaYOTfk9UMUxlJVxganzZ9amO0J0HDFnx8UKQmqUN3pFAyxGsENRZx
K/ZPWZ3AYTepvp4bCRMO0VImfokGfmtoz5+fGNfBNDn3UThzEmlYF+OwAr4jh7Wl
ItpntZOPBGSXIeOnh2HcFgMSKZpSCQkBMfNM34Q6OAjG5nEKVJktES6bYPKgrHMF
8T6vkmYHI97buDZxuf38p3KULyXNbIihIY3QcFiNydF9Ce7iHsXXyek1t8zWP7V8
g5jacBM8GxqNzdmhAmNQeS6/VaZ472B2kDWNiP0PandCowzqLFXXbqpq9SzavmRx
qb1wUau4p2drPK51+JakRUkHrU11ea/SktYwj5Kf856jimY9utVIogQSqrhledd4
g04jg22v8MROQB12oJC+MhWB6OTauszHMC1FVbjmoOqC8eTk7CyDDfklMRtl18Tr
tkrbuZtvJQsI+WpSDPHwfvvYftwWeomUn8N3ymkqGMt0WSN0YgwskTY/i3noOTZu
263heRrE8y2S/uif4h9A/A9dl1Djxd5E2dnM0PPseCjKtyJURsxultaSvo7XIpFy
bRjpzXYeUNIux4zpH/2q4s7nL85rvzYm7axiyLqpBJBttbI0AyHWOr+LlBvhkMG/
tA8yhVihCp8QUdR3/4ScwfQRafesnBXmMhbPDYPMeulSz/aR0bUqFqw+JD19pStk
WFCYdb/CuBciMkivEmVkvEfTwi3q2NTmnLvjP0Ol7LwyK3Ib/1BTM83E/j54bbR2
iktkBS5lU51fTc2TA4k6j3WpCBQ2dTEtA35BTc9qOlZWME75MpeDdmYQ4LpHgfpX
4entPmaRHaIkEm+Tdl9ZCjubg2PLXkVpmDVc7TNQ7ApAvAjXZGvSKrvdAYS7z0r5
xh/Lipvtzcms4WQlYZYTQsvkvrUXRBg0bd0kJgvPhnQUEWKryYpKbheZ7S5LJZk9
G0lzSoUAhj3+ZGxvJyG20sT+EZy5HsSzBOJt5RqZzOaQ/M+W6jbv77rfYQ46DP8t
S/RGiadK9PJtY/4qW3D3UIXUF9EdL5jZzcBrb39+dMAcNtriz59G3nrDC77foBMh
0S0zF9igEzDZAcmdnSdHHp+DjjNJh/6NgNj7Rzr5FnBSablcNmQTif+iUePnUPiN
dTDJ335AttdJZ7Mz8OYR+zwmHJ4GfnxQmGVwSSGMoUiaNIZuKj0gfqRP4BMIdBMK
vinLhCMQ/7MuRagjII/yDH8ntmTg93yqxLB9qM2F5J/vEXltPnHruLOWkLF5zrC4
9O6jiU2vpj/cWigp9LtMQ8at9/qqPc/JB/O2RxV9w3ubha8t0rbk8qumIzgYvt94
CYA3jKYQLKsMxJJ0DSsxmSsoqaF8BtNuFVuJ5gY1zp7jY0+pC8hjM5zMW7LjPBLN
riuyHF9PdRqotSU0uN0upF8wsFXDm2LGkQ4jUwtuojsxen4VPZ4WF8oJtLYNAnLm
bw5coYSB09UyPa2tNNDUWsDVAi8ZcuUGft/xJ0yVw7/GLMZIkDgjMuIyMm/HxQwt
UtAoIigQ+grkwNu6ypQeVK3VHxOppOgPfmoutRH575C2miSx5p5fP30dgIiZlXfn
m2DVZyrIPFpFog8gQ0T7dkZOlrjF250BPmkf+Kvoa9P31mvIzyUCmA8HOL+F8NdK
c5tEq7Dw3mO71D1j5eArogfjjwfQnFFIWouNj5WIIH4wvFRLmjqdmFguxyz4kD2b
yPfRtt0Lw+nltj0bfg/YDePoA07qd2MtNVx46mjo9xIk3tmymkdHkfFWeAslxZbE
vy9s38taULI1iMlX+1rhtjPUjxvy0ZCiN7fQIM/hNX62R/mqAaB5UqSk3i+Du+nq
wAUTxOKgwUduAS2Azr1qAbvCzbeHvNJwczVIqLpEu8xjp6NPdTW0fIMgUZx+eWqz
DAyy5xu6UcQqd7ejn8sxzS2S7mXrFf5UtJHhOiwSZwi/gGIfUgVf5eO6o+Fz/l1K
Stxc6PXDqKE2K6PE/9ifML8f34whpNDsOTnl/cC2IoJPpWNoo9FoItQBqHrB47MY
o4IYAQirqjMi3AlmFUUwujUBjjI3W0bm1O/9xOhVysa+MDOR6iADYOycF1ZJmK2U
1YHRXD77Uj9H2DkIHmC+Nc13+5ccpOKwAWfJEpg/Hli6G3x2svNAshls+d/WVeNG
0AyhPP2LM67tf9az2oZvwHt/6685FYPamkAXR5SBnMX5Tat2EvmGTOiB3YbVlR5x
N2zQ0i0yZtI8CoV+xIwSAulJMsRWFFb0AcUsMYeI218SQGWi1NaI4QyZG4d8lLsG
ovf/LPPR4/HA+QczXE+t2zhNVm0R40YKSXPSlhljOjLKty+NVcgYJ6XPX629vIYD
tupoXZTXCw62BEjWO0k1vb9gK+ifpWX+Cu2wySjFtMEc7n4pkDa/ZGQWrpdTjLK8
BngXuxZ2+/o0kK4SU/kzbjQgAWcQq1CV+yy3dCDeR7pZUSxNWOrhpJVqvDu/49dQ
4FKK4dMjgS75mMue8Opb9nTkrGSHq4e+VD1DXrzbk+s9Xmt4JJF1yt1MKVsifwMX
s3ELpBFxxxQzyqpd/xBZrVftnck4d7+aFerUA+I59PR8ChJG69t2uFnN7Mjb3cSm
+mjsUjDLtJzRyqyITbdRrLIwgDrw/b+xKJ1dSmpnmgcazAC8cLos4V7CUB8qgO/D
enUw8vNBlWWtxD0VYWVzV9A33yU4syXUqrLCazrDJVmouXeVHyrrs+7S2CM2aIWB
youaPuRoTDO9WDzP/dXhpUvPdOBp43EPMx/nFXYqvTVLr6NqF4rf2Efuc9i6l4qB
4/rw8LdR3P2EgEFyb/HyAJHZhi7MyYqrafa9c7cxr5QbfvDHaocPCyYuD1yy+Xry
Qgd9+B9cuT8GPwi1D/eOi3dNvk017iRG/HwD5SGDWo3uenShtafU+Z0WJlFk5tEU
YUAoS3X/xSRN63WP/oqblFG/JdS6rut9KTTVCZnD2MJAwardnzJzgQdw8aVXqu6p
p/Zoij1C34gvxf+cuA5B/9nFxyM+DLHiXsKFEcP4wQcr753tkdG5oVjN29SUEvB4
n+auAVjbofRNgBShWVAQpkjwW3zdi5BPGKlI5bdw5/Gs6osV8E+xCEvU0T/JGMC8
5qVXSASslThW3eP25dZtCer76/8PWmqmgOKGZ17SjcvVLoLvYpPXF8FcEqqYlx/Z
t6qb/nyAbT5dbaIGCzPZT5udfVKqFg49LTEVT7bclBLJW450JOOKsKZucMfx5poW
P5sEGNs6i+x9LWoDrAqHHohXg7qg1D8Kl9q/LJzDwZKLWuAdYRJ6aIYiM/rkXwhv
UEpKnn2U9BL3peUVf7IjPFO+mtAffUY53GTWQHphCDUrJPzZVElOPqBpnW5t1n82
jfOrIFLZYNCTWd3EgQyZCWVelQ09iKmU7VP7Bu/VBGBmFLHmgFcvwAk0hkyvQbnz
RmPfMbWZHo8Hw1RlaxxkwPQUyJx1DozG3PBDXWd8v8Q935m2D1vcFO+JJzh+bR7j
JsFdhI0xUsyqhZdrQTxmE4wp3c/j6tQOW2cZDGFCy6jZCLVDLuZYeN7v6yB/eSlO
Sdmz3Hk6GdbCUBmYKlKBdSzGP9CGePTKavvhGOEcSl7VIMTd/nQTsYzdxo/1VxjA
RNWeHCwO+oYYZyOayqR2gWyzez80YP4GB+yQWlF0cEZJBRVALlZull8FN3XfoGur
xnHMlHbUlNDWL4ye2eGE2HpabiZotd6Z5IiH8kMFiBpgzfCErXvQsjZcpxj3HIGv
n+8jR4ODdqu5kXQG3nz/8/3DQrdK64tSk3cKeUQWZFtC6ComHlhZTDcpXiA12hbS
PJcWXAn2IgWEfI+/ZfQPd/a9LOzcGWYRdV/B1clbdGHI6pKwPj1XLqbIfa31XF0J
Ga1ELAgZxdZeXaXUtX2nLvNRn2qIpX2DCFvDrJhm9sjqe5exU8Xt0lYnCjvCHBEe
uMwcEg3dLcev1ppShhzRetse9/aMbjtq8iC9y7PW44eB8wOIxCs6yj/P5eEyr3c2
ZWcsfzKGhBJ5GMaEZi+tRAxzM0MrXtC0gZ9sbu5fjK4jGxtsWbRBiJayv2hQuk81
ZpG+j/0hQch0HNs2/4aJTeaG8bU8ItTDJ0AjzpdM9+RBV9s++WqhuJWXGwDiCG2G
NOBobURgimhAma8VGISEPR3mFF+i73Dc0TdpPH+ZXHxOI2L3OAjuCbZGnNq6botV
dtG94M8danIXyEo4vGeYZIOcByDWFu9yKOLq2nFob9RBWiaIxTiMbDeIKToLu16q
0k9EHIRGfRex+3Ew/sZt7B3RTNjPCcJpNLCuhpB43GpM+7+m/hlaT0HBBt78JMFz
MrV8G/XGB7bIg/BYhkLKtPk19Hn1zY7FGrIa4494zRwA52/Knp7uLn+QGa2VebwF
9jBgMIQayX2QqplozS0AbKhfGCruyCwMZBuQNaFGbXeOmGrnRf00+J+IR23pYiVk
Q+TQQeakwCUPRpi29j/rmZWwLYVM8fAxZM1WKwA8Fs9LEtGy8xWeN3Kk3B46JEIT
TQr11lSdrmT0AD/4pnVs09pxcRwl/WngeV0Ab6vOI9JiYUZE1bN4Uo6t1yUhfpSC
iYdzckKqKHYUaB7qokv/WJzk2Tsnj7cyp872/WxMY7cwYCEirz99AUUoKYOsqlbd
FmBxW73+faX9RE3HOK/46bfHo0XC9Iqa0PE5YsUsyelWuPHdFXKH0cPpprvE8aI9
l28h+8oD+LsWsaRIQ6OnKrvqM8rRihnyPriEP5JGfquvCgndMEMp3rcIHss2ZzlY
xX+lDYTmxb98cLEQ3p0lY88tgwANxaGPohDadr9ljbZBY92X7n9SL/IfO87LO7py
Cux1Vdvnd/rw0IVBtvXyGGKksgFHyWnEcSMYWdlyOjnY4n9c4KsrIAZAIWTIPqvl
1/5e8ltLkucZP3ZLT5AENVPFZlYx63KYo2ksPR0l18DaWz3EW2pWDIxar4eNA62/
0p5ikI5nA9E60NHLrQ3r/nNevRS+hTSyrRl/stAtRB/SzmvUoCyLiJrnrzj0Htk6
OrWElXabxg/oOzdvZUJAAo5W3DitkEq4+XO63CjBvDecBySqS8egs6vK+ePVkZye
06oiG7V8+X9VDlJX9BTMV0FMj7Gv9PL9iwgbvDhEKlirOTDCuFzB1xTca/sluDiK
DJmj+3uTZbBLcLivwsAd8jCmdTh1S3NQV1L1YoflMPbSdeZgeAl50bxeW1EoeQG3
9iYRLSTKOCNi24oWXWv+WbZP8F6SFD9HmBmYIsTUsQ+2SUHaCU5eTYrdhKJZunRN
hIBtF1aT5KsEvglrzOfEw6rkzMlg85SzwJzPGywZj6WitB3Dp+aSDn8eHEG4tFrh
Zl+BhRN0SVMOtOvUJ3zF8MjHBoZTpr0M3FCn1ICdp20VQJL6t4Il98FlyT03/EBH
45AsO7q2DSRhS/Og0Tee4NanJeUYmJUrJ8UXq8E2PFdoHySAeZC7vBAYq606foQi
0wt1tM7g9zi6dSiLyomN82ELdvQRzVO7epIuoKPIAv/QdNtmFdDx5PBfuFjUzRga
ki4FIta7CJ3j/ADDvFTxe3Y8DN4n5idkmYly6fVnnLwRPHwESZeNSUjMcCqrs21Y
wTU3ekY8V3vVyMIrkntwytVZ6NJy6AqeflGSbq0uFsUnWGAiw8UQ4JAnlg021Eyu
tR35FinZgPec4QV8wJdCVqEGT2F9IdVOqivBx7N6dZcBkcd5qCko5I70w1SJKipK
LM0NcXjHmL0UThc586xHotuFmCFqQuPw6b0FQq54KlN+GATl4/0CNcV2lITnK0/B
yRmxC0j4zhj0kK8Ldh9l1MJeE4iCML7x/WPjkvudGHwhTb/NPDUGw6VY4IazUd/4
NOrc5WNMaNrg3xU8jbn3/lG0R5qb5piUu7shChnKa1ugSISx5SEfvdbNd8WGnMWz
l0tOEmNaEpfJ9BNBsBCKLO+vB4a6cK1m5eLZsNvfukxVrvOzjPEmXBsi0j97mnGz
ph83N/XJsQfD/sAcSsMg3KbXUl6u2y/5A+Aypr0Qo/7e03e9GrmL7NlONqfRMFqH
y97MgqEnvMwABKbPPZEw7xwJlhND/asedBbW57fh3/ziG99v8nxf39JpQBrIgW9y
LFM/cdMny1GpQhpMO0oVWIyCuJjzyY3LxopEdxWccgCuiI+UahTAQo/hpav7op8f
wrjRKsYyWynYGI1OhsgzqAaSM4eybnjCSboXjahUv+daKOqsfQNE+LPQoLHxTmuc
H4nFkSxUs4OakRYo58fa+X+Gr1A9hhefW1pCa2pSdj7ccHPDSfIOUOIzej8SNeBv
dUqrCVzt8Sbt9RRQHdvHY9iUMdO1ExtyTE04Q9s1OLTzrRme3M/xLMkzn+E5h6+k
QtlmjNH3Pfpt0lCXv53BHU3Ts0nIB8Inxv4HorfhI9ITjguVl3jLTiJz+yzG04sN
FoWH1LgfgdvsP7PQ5YQ+KMlCbr3UtnJtw9I4HsPaXEFQqL87W7PcLhUvBGicBX+Z
NImwi0XL2eOgXA6w00UHEHmD3RMRNlUOWutvKh+dnhGKFvbUNdJBKctS0Nb8w53u
gH/Qr4clBtHevM1NbHT+M0iAP91SDcZFgahHwlpEMabg0azytl7I6TVdrSnnKEtC
VLIbdHG4uZzLgzDwlp3UKaCR6z1axO5vow18SmlVShPUh4nSP7dqOESUCVJDNk18
cD13ly/pxX9sZm1cctWVYil4ccrnakarALkYLRI0CL1iWBSirlgGZGeVu/wlFU3e
N+Px6M7z2un5sCETg+5FiZU+x6662/PEZJGMbrZ1SiUwQz0qbz54Kl2iBN+3OXtE
DmLNndB18BivE/Hn74+Jgt6UoTfi76Vtgz8JMPDnawUf65tRdusFHXeem7Er8u/b
+zJWGj26I0j4D44GhJx9VuMJTSDj6ZHPHHqc+nBy6LxouxCFcW52b2wPA1P8uGmb
4dyB6EoxQQQYeo0R8GWitUymGKn0uJ2K7LMqXe466eLzVmtryDi/YqZZPpR53+0o
vdPRqCRLWaFMgGvZFYiR/mxc0tPRFBhs3QtfbcpNMm8652nOYfKTPjIzsSc0RuC6
JF/kG07KiJmGKb/XnVt2I4xWWMnl1kA0BfH0M540e7WZKPvoSbZMNFMOellGQlcL
G67semVfODpKh4FSGiRetVoHWp24M9NXvba7yyG+JGk52/SqlSfP4Nu9AWMzPfm5
GnrgV26uqC8q4n7G/r+/OyLo+4f1XZGrRxwSOn6z20QF/olfvQRX1DI7hWl6RR29
9aLTUMGh+ZDLKe9O6/VFz6qeNjxj3NLKXw+cCF315s/75rHXwzdVVqe5ni/oykcZ
1fAnwQBSTyIuucT2M5EWBPrlcHJaCwxwECWJf07pgAD6hNFirvLWu2s7tlC+jWge
pgIMZoxfGo8MM7qgUxPY09M7DEx9knXu7gRku4Xf7T4ZSgWecbmN9v5oPeHGE7Sg
5g8+Yg7Nzs0p2tyN9bXAx+aKoh2GdwxC59gCd3pA4SSf2oZnNMvaIZOoPdiEMjo6
tyPjZ7lmVAfwitqP/cqWvJeJKJmCWHzVTEfL9hw5tbSObKjOGof/VBDZb3VEkbzh
mAOl398ddEm915YXoRtyN14g2OyooKku4Jff/4+L0+zuRKP4AOcsDeI2QSmS6V0w
yODKniIFYDtt0p9/eRs41pWsgLBOGY+ZEgkwod+oCBRaWp2UcPU9wpqPRhck1ea9
WNKnxEjuaa04h/5zrOyOk4sk9h7xLgC9I8oMnLBF7mT1kkOemCOfvycE4Rk43MAu
VnoCqHzEhoyqvn6+65ikuBgiVz9QFW08O7Z1ZRcdUPng3tJxs9Maqf3s14Aa19Lo
CfmiD1dfw4VuuON7Flpo0pIWxURqKuA3j4RhGFDBHiYbJCyb21KVHtyZXMTKHWVJ
oPFjnlSGDurxlV3Nypd6YVp4fjwLqofCpZIOsuoCBSlbL2k9GA51dT7hcLZua345
wDvcuQE3BgqIf99ZZPzqHJAnYDqVxP7lUb1OCYEkundt0aENGj0S9nytCY9WvAMw
nGPuGk29j6Ayg6zeqKIuTn9TW7rNlK8vBGAKonVyKhd3kGp+NLUFSz7r8xhA6Evb
H9a4GY7b47B51NHUtfTpXG+1pEySgWu54evVfOQZGcWdITCFftyxR8DCTgT385rn
oVKKpPHs1lMFl4TBHNw44qDED9HLDPER2DBKDphW2dcAW88rgQzitGj3HAhdNlF7
lj3JR/ORimRKL8XIr3w9Y7UXhVuBhlD5pJfIyKyz1q4lZzq6mIOblTmTC9zINZiN
/XSJiwajD4dyGG2EH8h0urvulABUIDIuIdky2BSfvLaQFm6U7SrcDhXGFKZKiF2u
sf2T7Tz8NG2JwWvvgWnAReNgDA4zKtTWMhhiYg7JvFydiivArWkFeYBYeR9W5eSS
4RoxpZj3r+KKMEwquAaSHqEXxZPonebJFd093NSEFm68x0etH/W8a1RSPXC3cj9a
6dZTrGYlaO7WfWul3A6+CHadAlKTr/lsiizyECRUWUkM9TltKBpwSgvxQOcmjjYp
q601rFg4mNbs0hTJrPU3FEPfOrG/CKUqJcr3dB9C6v0wmbRYGG5w+KHDDVJRK2gT
xmfwU1koTUpS+zZlvw1iLbdLK9a8ueGlSz6dm15Qj7wrz40leQCE8RzljuSaJKeo
QrfYZYg+vPNTgJwl2/GGkzCna9ZqlBnyOg18/dkOUV6whXYZqUwj9GIpi4Wugv4H
F3wDIQUbTFkAKeoe4bvFsib1bLsrIvzsd2lQddrnZzMhxcRH6uUuawcjNlbWV6jx
t5ebhcsILtek0d026RN1oPdVksYg9aFBv5MhU10zO1VfI/hiofvbUH8wl2E8zumH
RE6Yg6vl5+5naNVa4zR/+oruGZasUdqiUXDzl7gxilIGVb3sKY4TNHthS5fp+DEb
pnkpP09tbtMFzYTj8wQGBn59kT4eSXiwBfE9K9C0EloncFlgFZ/tywWo1blNTjuy
X+/InwAs/J7Kda7ulXkHEXAoyPg+/H4castOjXNtum0aSB/mXZNi0cwRCSXYJLIZ
u6ZeDaH0d3fk5fkebBXQtZQ/r/ywdrq0GtRtyZMVjg5cgf5j/n30Dvi2uHqiJgh9
j4rSBkOQTbnxtV8t8dt0mMx2R0egnjypVcrZTdO0mdY5F81XcdkvXgHaofJ02FFx
cdsvCDnujHf2NDn4ow417NnMu4bKhdZXwGCzLpYh3bzFNUJoGjwjQ67RHb+kNPLa
2GQQX5S1Pp3oAw9tnapoYq8c7g15Mwla6ig009M5ldbmxjphkUZSogC2rBvjV/yQ
ybIGwNtXfHPWdqySLG8bgpo3qDIccjgu0tGvCIKFjv4ayAl8cUhA+FfKMyWr1d6R
fHrKhIu2KxQTuL1YH5poApRhFRvHtnEkQ/CYdVu/h5lyzkn8Rx3hYe2PqcXuZg5I
Q/kmd5X1FuBYhxjKbBGMRdtqnoUVxOS1es3DuHczapYx2y8GaX5ye2ipG6Adxu35
88Vj1Ogal217UDOCDUtArG8xSjAzYVanr5nUfBfgeycJqd3Kxkqw0PtdPaB9GFW6
FQxe9tueyxKRfX8SetUndojQjy0TAOQ5/YVeUUiBMUbNuvI+B+p7Et41jL2qdM96
pdklG7aD2UQrh6AqnVu6zwfC38aoWP7VX06SMUXnqKJ8uJj3ho6EynHyIiT3a2vL
dkcT0CgXl4HAZBHz90Y3IqieAdGK5uxOFdk5XB1KlqzDAv3UDZpNmff9njlq0kR4
flPpBGpOkbck93hbmo1xynM2iAYYGWfdY3LLGS7jDJUpJNQeurgrm/CLTkTs/LZk
CD/o2mJ0of/vPGB770Hvpp2YJ4lm74qQtsKg/bPjKKOr/qCFIPlc6sc/2TH96n3n
+M7j3EzKqmUunVcO+IHnW1NIkwPwuWULG1YN3SHFFTMD5NV0MClIWgjcAWqEI/+h
ArZ1BDoOPqNxriNvcnDzh4Hh3AVU/qsdNZ2KjpW1ZWKEjwnbrmumJN9jxrgvcj1C
fRWFywdD0YaWOtr6y7u0vQDzOkk44zudYb0glbHz/p3r2LyvQB+XwmpiZST26XeD
d3EUpWMSG/Zm/WWrxvC+PxsatOi1GUJAnRFIxz9WBbHXUNKz1ZBOxvb3GbwMaXAj
9kFrmbcFk8hsXXw5kL465t5e/ptAeQSi3xEn/vwnoEtJnJYkGV2GJXLXi+8u+d/e
zK+ClwEU5TtAVvy0f566TquA3oQ5ZkIaFABXZHHJZCT8z/bhV0Mqe5FdDJ0MF9SX
zu9ovIVkbkGrsjL5cjC7omH6Z2ci9YAzm42uudkdX3EKCSUmEtrZrU9Iz5v6noL+
7CJ061ADl/dETb+UWpy8JhypI9rzT4IrIGFSmvrfYPQs7+XommMPSNVVrGInAJRa
naxS2LNcIiLsqnt4vxTX/ogNPeVVNDQV0Zmuwh9/j8u2AxLCECF5xty2X/rr4U7d
M22cWjgPW/J1dN6lODBgj1Sq5onXqzaiCjtBxlSmSN4hKlSBTlXgTTMBP9vMpukk
pMB5uvwPUICqEeRGibZ6GPERThozF7F4bwzAtkXeZpc0aTvhKU2QvDoa1nA3MEHU
uIJJVZQ4cf5B2Sppm+H2W7Dz7TO33tk+pePqfemOY+tDLjuLmh0BqKdPKN1u7N2J
Pdmf/kbPFYpi2cJeKUyehONpf9V75Xh5fIe3RKlTyqeWR4xl6V8xzy4m9ORj9Fca
38gyH0Nd2KR1xDtY5HdJg77xrtKg9NJaHrovohdABo/O+ITUHurSvLRFc0FXX1O5
dElBKZoq14TrsV4NPZckNeBXynE14SSHjLOAocCMsQ2tYHUc1SQS1mhjIuFrmzK4
+G1n6blrg0l+U7gn9sLE7P78tJ5bTK7CsQmObLsFxf+6VmO24oAr75RbQ9ARLSeL
VQwrKBdTmhK3dqrIhtlDtPK6G3neJx+AQQQWh8RRaRI+pekWZ1c+d6blBIxLLTme
0FWIpzi46CHW5ys1OPN03UmykYjdhiOTEYkmQq6dO9vims5+P8c2fPFAokq6Hv7E
myUkhaFQGy5xABRsHzxYgfpQUQagVKq3hWkHLOyq0+j9p9noMHkkq7cUayGtSZdz
HVsveph9Jo230K0FKXNEbFA11xSTBRnmQm8C94hBdDJbtztlPn6x027Yp6b5BU3u
CZIWfEPqsrdMQ3AzniVHCXkVh8aBZyROarEZXrIW8nvmUKBYm1IKnZBFb5m3EWx8
6mzrZ+gQfUCKb2YE4H58qruJHm5CvvkS9xBg3ksiYS/zTLnI3kblbcEYRjp7p87E
NzBSNW9Vmk3i46BNy56JgVUXAv0XB4Bx4cvdpWLUDFYcx0PAk8bxCBRNPtVrhYCD
plEyRJpazNY1KEmVDgWcp02TDwYPmG5tojQdCzTb1VCZ/xJDg7B5/Vaohnbzfu+g
KILvrclcsdtlniasscYa7wsi7xO/HN3ZbgweUCh/bhEAwz9mcQfc1rLJ9+2MNqJL
77x8dOx/YOCWgxkzRTpbAIepasEdqbcMvof3YKkCGjZJ6Iw7KKX3ke4VG9I3VHDi
nFEK51iBnqIxucLBxNrZCcg846pphmRKHkwVO5DjdeMCMbNagDUdrR84YZE4/CO2
wc+DjfJr1p5KE3/ioO0x4jttRfbuXV/nLQ+0djBTYTf3NiS2Xdt6g4r6j9SU/+To
bs9+CQxbnDH6Rqo+rVDUkY1a/4y9XUs0nih0E/LR3pRmdapBF5z2Xqtadn9GiyhW
xaRBZEj07IxMroyZcDiBExvJHdsNK9mSgwNwZouvDOHH6uErLqZTruXp5gQh/hOq
uZ1Dr1oBxK8UV3ro7UmqNV5HwgXb8UMI1RyN+O1qp6FHKPbpddvwbKS8W6nGtWSG
8Fb3LrDVAi8NnYGhbSbQ9gsSrKf39omsfRQq4Y8NeGcnQRDhuUIRGRwzHU3VOzsA
c9qoB6/cnK+rKr8ZiNyw8Ibre7HVJtMFcOxikrojZIuKpK+dcNrFKcLBObyYfeKz
0EwK0rJDkIoHTM6wXNgRiMkXme2l40CcJXMojIH3wfbvMQLYB6uJSTBJ/JWgHVR6
wKxo+LwP3pO9BMoFyWb1dBQUq8wJTBGXs1Xgw6+WbpOJBl2D5Wy+uJvnHAbEx23z
GcGTcGD/s4GOeJg3K/kDONGLDFDCf8qBoVR3r+bYmrxg47ID9bfhls6G2bEF4bDx
grz6dXi+p1spI3COdmFa12f1hjvPdpWnQAYnQRljuXNmrwf+gfhHK4cu3ulCzwc7
EvsYCovIxn43mC0nrEvKoOnmu1iRuDwJuo1iOMoJr3pffll7CHfYH6pmaUgUXrSl
GlOSVAJAnPqp6BJ/jKZSZMHEc47VCEawvC+H9J+saFKrvzdE45WQFw3dIhiev/cg
8sQa9YZRvbYGapIVLwDdIk70TPEGZShAHgxyRkEcLizbQPGaOYqHA2clZx5tbYKL
DvwJ+hAJ7oT8R6VegpZplpODi5EumkN28I2APMXykSnQgYMZRhRwMh68REa+mMnD
NYWchtpRFDcJKe2EE0jCDFo/3/PFNfEuL0k91+M2uEtuZIK0qC981rZjYSz/fWjH
jBt9nDMg6YX/Qg6Zf/TmJ8xpaCtXrAcSb3G0Gncq/1EkYCzuxGgsYYhGJGIcWuUK
eOIQCyfu4gxPDFdgl32b4g7Y9D7R3DBxvLkb2u0OMmBFFKUsZwc1oXPumuf/Z29/
+pAkyRwvfYDzayOWUPAiEv7aiSZUdX1+m0aoNP2iAYk3KJSUK31gRQGXG1YgkN+v
HcNjpl08Fy90LOxNoHH+650/PdJrdKtRIycSWpT510xxm7bfLS7AreZP0qON2RcZ
fkDUDWySzOVV7JwL6NzMjppNmt0oH9LWuAlrL9hkq6WKhc2Yeb/CCo+0oz1Tu7/g
J0JXsfJFNIzuDnvUMChkW5sl57wPDliao9a1FWiO3e076Oc+Vcvz8afPoIEx5e3G
C0jff7SOe52y9+diKMrs9UqpHPOGybkvny0Cq6PvSgG7KJnoBUfQivG1IyXaX/rV
Vgp3pSj4G08cg0UpACnVSfJrRUP3MaaOZoLK6XGsIVWr7dH60l0641HQOteaPhRu
I/Sj2gpGSiR8lDmAHtpoZ8TXlsq1ZlKr/z3Wvemvf50Tv+JJuJUaQs4OS6IgGI2j
/LNwE9tVX9kMP7LN2iFLXCLKVDoOTY/Hn9KloQt0im4l9IFD15qnk/CZYQdLXWrq
BI/tLfFAuDFRhivfYNzWxNuHAxnI982xNK7M27ZJEcH4rI4fdAxBTjQgbvhqee9X
JU01YDEtiEYGP88mwwv6SoOrV5HQEvVDH7vEjMWAj0YTedBa4GrE9+1JzgGrUeG/
D44ZBMaSBxsX9pwMOdq4K+LJ23guxu705IkTzHxuU/qeP6nHkfo2sQQBFoJSK57K
+VIC1JCvkkSaBpFTRkrR0MMlkJug3JcchGtQs+GeJPf+je1c9IsAFfu/UOFdBcKf
ZBhUK9zTwUDNEQRSPcyqLkzSfK+CH58ntDnxWUGSz0vQQF4F1RoXxVOB8SG5VIZD
wT8rYD55nAcQYxl5IeNS4+iYLk+Ugwrcx8cpmI/MvfRCAoL9GaP0+fIuXEDmOjGx
CMpQMcodhLT8LpFLCwjYAWjHovb65YQ3rtfsvUYppDS2wASjIc+7gm8oh7ScGOve
UjMImVQylag2AtLZNC0aNEA9rotJ5mjcapn9bY+eqA/paPszkgbnjZ3Z6UflAcWW
asX8Exuz8aRbO1CqrkOAM2tFRBRX7ipmjyLBIZXc6vQldXFpLESykOcT8+UfNof8
SL7zr8aFky++mAbHMEDPolKseDW/TvM8327v5LbLbmNMYOmdZoFcWqqia6g7pH7z
CA5MQ6r3hdap7iF7vjodVUFNJBQvazbcZ1VonEbTuBUeNe1ha1iB+KZMbwXpmNCk
AArM9nnSc9zd18d5UU5BWfZavMhBaSYwVRENG5eBOpUA1emoL6dzxFh2lldSmyPj
0MilB1KQNrpN9tkzSvOOGUMYDn2l2K7KYYBa/SEFBcsZLAwsT8z+d/aMp3ZAMOFP
ET6RLhYVxwpZfMt1z0xlilb+ppIrTPyJr4pQBfPd6alsER0+iYz4fOfhKNlfosQG
DH4DfiBe85mTEqnmc0sieV3nbfNIa/em65gh8o8qOkijgCmPE+fJavTc2tGxdgGU
JIKTNkuRVWtY9vwIiagfPcg+SWOV7nQxBqx9OUfiQNgyHctEFchOUqlVCuC1sh9s
cYz/jEzDTijflrLug5+ZJ9vgnG9jFZCsBI/jR9q3zV1Lkev5cwWrPoxdZVbqno6X
upFoAiLi+XyBTTZzx9fqPxNkox3HbRYOuqtmXpx7gzQJtUxBDk488mqknxS7SUz2
6NZ1mM3e85+crwTh8jtQz9wjW7pFGhvxlKaFsKO6rDjYtXfBFfFF0EQo6UB8+rmf
yPkq1ygQ9rNwhIve42nUtASfGXa1FlE32ar7ucQUH16kSA8/YyLLIJwmuf4jcHBX
I3it24r/wq4HQMxY6zZhXvH+D2L/XyXONEQ7ADrZnBF9J5Dcxemzrbi5V3HIwF/S
azjl0UA7u2usCXGZBVYwMOklQUF05tIpp/oc4rcTpVX0/2BBxeXEm3/HqWLCe5y8
t2USLr/VtQcZNZ+nlekFS8nYJ09LxOn5+Uvt2xW6MUK7sbpR5N8iunLnN6uO2fRL
a7NJNFU8WwBRo8ZzkQv+R9YpLTvx5uYIl6EQehhnlMczQsP6R3w2fs/BUpJkJv8F
yHpVnu/5TyapIlB3YwLKVSaejjdKJbWnEvePgCIpsRra7vZvC+thAGcp/ytaNiwe
J3d4bgY8gFOAVfgHZz6nxTJEy6+6rGe+3+NI9XP/8VjDCsrnzFxmJvXulXdRmMbU
ewHPJbiSsy8wJZW0NvrvzzxayORkhIYFPIY2K9umI7PMbnMcnuOXjPsPnYhHPRO9
QDNPf6UxKhwwGdr4dzMnQthIdGOzSXHkK9hu/OfS8oRzfwrDry2ph449/JKZDnlE
DtNk1Bc08NOCe5fnAHDIuIpuRJJgqf9WFXphkXEylSK+9QfCJN+JG6iAfdL6Mk4X
vfHKncvo1PMVmyqufUQAMZ1cAtenK5X3E8S60+IeAdaVoYRfcZXQn7hoaazT2Mdd
igYcNNWY8nEOPMg4s4iSMkRlPZKboqsnK+NgY/VUQXWFkGJMhSpU80pRQZyz+WUt
9kQyjoCmBLwZ7TSrgszQ4O6mssbHWOYT5sQusCTEobu0QT9slBkb+bGqMkdrpRMj
bDN6JVKy5Ue2BaL07nDnQag4RZq5Gr9fi6uJNQPWihAPJa83DpQz1G+ER8KzwX8g
kQb2Cz48LxJp0CF5yqF4eTuH5VdwJsq8g4c9IyxxE9TvsYNEWMXUvc/eOmys9MA7
pyqlZXzaWo6y5NXqv2mAqEt0FLPqaOoeHVMMQADlz5NB76jzfcB7eBALSDKa7ej4
a3WmpvnSYCVTWiqMsB84ubv4GwWPvOnnBYOmSWi5Io6WHTiadlxlHpJoU8rS2dET
Fwa/ntjyeMaIxBywgxZ2yhx+pIJEpXfEQDZfaw5AdrUVkGDZU+8HnaVSg95OoNVE
Pjp/8255DWtr/vGJZHqaZwpOnoNSWhSXr2T88Rnhr9V1NYwusuGrwoNjkHaFNSKu
QpjeYBBV/7Ay8ft3IcsoZ5QZ+nR9MwWSi+TGyH+N1M0rTYm2VsPdNWLRC395Ni1g
YZyndsW4xxEjMoMPHKuaa5bDpyjIRw96fiFExB97SnULWfLuIru9A1U9wXu9zLa+
bEs7m5/s3+HKOBm42BJKSPb/RTpLfR0mKzNkuBEBm4PynUUiNAiYPpwPvteF3Fzb
H6ONF0EMwizG9kw135sZSEb/0NvdaVyWZKhaIA6/u5SnwpmRTWdVrvaMNoqjwR9v
ueA2FzFodf7X7ssHH0ZVM2dRItAFaNK1M8vqSEn1KqSFDS56IrHRbHiAsg6ZPh+G
UR6bePCIsA1rKIbwaYzpoL/mGnzcDzakXGhvjhpHifE7ZReWsJaZbgFZfVE/oUh5
gr6/mpg2sS9wOu3/dsjgd9ie6gEr6BWPxBsNqVhY2nIKvNcQPFs+SRgHsDNaMS8I
uYJBIntsqhVV4W2yPmIjhisJJPWeSkewk0FLVbqEP53aSOTCLPtDh6VF8P3dFLFb
tA3McNrvJ1rsOPbubSGYz6WRmUTZY8dDb+O1xp5xHcUPQT3a9T2KdUSJnDpHddaY
cEYZIIwWkyiamw0IlLJzd7HF/GivpILHcOV8kb3HQr9iG1iaVfDYpkhhIHG32Xfi
L7El3Wn4gqjdDSVqZlFGCdnYPIP90O1fi6TSt5+Cvz+iym7/GJAVSRjP6N/cdU+G
YoO8tPhUXbRbKy4hsZVhYsoeuayC+HeKQenuuOU9JSv0vITvlFxcq+ucV2e6pnaU
D4fuCEyuaY5rfLT+RyFjYIBb+CjklZnID0AgxhOr1vGcmUXoYSmvcfrcVA5HIihT
uJDtdPVyVSf+nypLqVckHrW8UcdrZBt7MGhH9YyGvoZ3HyBXR0SutRmG+GHy9lIn
IaI1oGgSgAmi0oxlDzza4cdHPc5APcikteYuehdr+gjkmlHtiHr6/0sHwzo7EmdF
qgqCCkpvGpTIFsgytttJ6PYTkLP6sEkRnOmJDdot+WQ0Zps4UliyM8L6WUAAkEu8
TvTK21INEd9zxXRMKVVYwjXKp/wz3+povk8UtqSgQiQtcw1xF7+kHBazTLZkl1IH
rj8O7adnrnVI0L1eF5T02GEMYMCSf4NnPD/Sp+0pFcmgTo7UEimld9EExd4LWYvc
D6BcNUlElX4xB5/AjPFU1/JEZYlI+4VZHZ5s1DsrxGp/t+NRk6rldx/oCI0CsuwR
MNsTxhQcRpywHDYgMjohn4O1/qdVjuOhHhxYyv2G7goKU/aqKI1t+EyeU7+FfAt5
CldlJlC8zggcT6Wdow8a1FXBVxDZdRQvvVOr+biLiWDyhGTH34V+lVfPcrWQxeRB
M8tu6Jr8tHqm/+XXY6/j9LL8OEEs05oq6wNGl6BSXWiz9fQwU9G3TvxduPFcI69h
KjdAnlDyMN620bKvk3yk0qFVnCoVP8rFqCPzjKJGlvn5xIxGnGvfMoeoeGh5Gqai
JCRelx4uDESTh0tLFnMdRU6Wr0qN74MOLmoBDqb0d4CduDoL1ZkUPv6Uh8dobM4T
CTs4UPDmZJAp35FSK01RcBsEQqqCX3JoGKgREiUrsW2QV736EaagkqisbktsKjSG
5DwlBA/vAgOh41PwSzAtHAE71FT4ddtLmkLxs/FCyIeqwWRhkz8mlw39+VmzHC9H
XkRsLnsnp19FS1D90xB0lyW1ic5Mq9hd852K/Ys5GznAUFUfA0GGoRNBKMeebzd2
MNIwGYUQfr4s7UOEBj6egcrJ3JJwy5iq1ThWVSn7dfWr2T7UmLOzk9juvcqbBjIW
tl+pPgiLpwxgwsrESeHkH4VoScDLkXcfqilqfA3WWfgFr8cgIHcyI6cokI9xqV29
AON9ei2TcU6sVbUj11cAD04L+mERtBqzy0tv8h9OKhaQsEP2liQZaOUK9atIUuHp
35cHVcEFFNwo3MhF5VzpWxGnE7rTW9svDufEydQTndIwZrGcEE1OSO7TL1RDgexb
O4knXG0xUuihLeSVHdIK1n+9bhbRetLoAbmri+b9z9K73euOAPLxuE8CBMKGBU6T
4ZvGT7fzaCoDyFCrOq9E45RuCbODYdGguc8Y1z+rgB8w5KM1SGbcq7akSxFXSOSy
DnyTyhxzj8nTisGSPvTupcA/XnQgN5WTEy+vTSmHU2rl0w25MR3EjxYM0fZdkfE3
y+jUkJCRnobKmnJI2eQW3TL+C6t9an3BlgaVBsTmITdBIsY0H1WxdZ5YgJesE1aj
yn23myDVLaGinJpVpBtDFiNmFX6rSCtJ0tqSpq6m5WB2cIUKcjO+JHdAXUpKPCB/
5PVIZReDlttcIq4tJZhUtVnlDc162jXJdLp5Y/k4+RdmKTrtqkwS3bEoOyA+H2o+
EAq1SgsbAT8QyJ7GIT7pQnePYS9j5GSmyC+SBNMx3NipuLEyRNICwuVb6iFvKz8h
p7Rj5i97vnI0cBLluxt2vJ20ZTObpg1V4dCitXlmFh5sYDJg4Of8p0PO8dbPCBH3
Y3QsUuQb1XI7QDX7xJTwLeAuCQGWU7b6TJ8Dxl+1CPO7I0INX37EnBnzvBmpjaUI
MuyPCWasMkv7uDvNqKlfLeBjIzKsPxTacRguwnAdoCr9KdZsPDMu8ZbQmB24ZZIh
AFAR/+Vc1eVskysC74QClWp4EaLt+qZce2NcnH+DIb9wg8Tqp8e0UhPRTbLi2Xla
ARnaYn0e9LxeZlqdGrsPPe0aEA05H7Vjc80Gvc3IFH2ebnWvFLiXR+AFadq2C746
gZXNsemJEkx7bvcOgaiED8lA0m2TV5B1nOlWKHOjKvTBY1jaIauWPrDenK8OPBjn
6rW3YOXjFsolg/lC95j2c7SjjVTn+3IwINqqKzy3LeITg5YbPC3hRT+zZ3ReDjwR
/GTwAIgV4EawTTXvyo9nDv4BPzC+E/WoTnUj7btZlO0oA/FEEpOypLqLjksF8R1t
zYYO/xQU0esV+JXWmKOShcW6YVwzFTr3zaQENu9Z/BZm24xKfeA/PuDm+YReo0Dq
cvmnwZ5rWkxyyrV0SuJfwYNadxmPOAuuIpLKUpiEeiqvaSGTudm3lG1BfmCcvHlD
GUSqyTiXMVlYXc/r86L9xz/fjHrS06yylvPYYsBfmj6t6Warn2yz8mkZqTV15d5y
C1tHys1rcmZjjs/gPlkTVqil6eYolqy3GkQO9c7ULyXgzh9Y0dnKOdrvmuX9cehA
u5LA11xxB8rpYq1OaJhPxKT+dtkgUeBxiX7x3WUR+AtI7n7rLM0cgiz7HjciKAtz
xf0SmXKCBdEANh3S9ayB1uDFZR0tISaE2x63iBDSkH8+Qdp0t1tM/4dHowOv5FY0
0giOA9xPh/Jrql1dw8lI8t4HpQlSDMQNtR4iLiHCl0uusO6v2Ld5dcqa6Ic8+bi2
wAgbhA6zp4EkCfgYXH/X/iKDzlMnlgEqjDLYcYOBX2iBaHuztH7gOPtmN1pA0wrY
Ah77njCAJXFmxqJYLGathQJdJT8Y5EWwHVN4wsaSxIg6CgxZhITswl+S5uDB/WxR
hLOFwvLE5PjbQs9xD+fX3Eac6Eu5jLPBjpDMYAQuITqyfgpJLmQJDk/Ps0dWBeGE
zHDyLABTQTlglU9IUwWeAo5NghClUuJLe5F1WyGk9kkTBVpdA6wdzJib237CZ0C2
vjmCwucfrW7wdRYGjwv+i6ZfWi51Xng095UjUI9SVRTuXHOH7Ng1YC/KoE8X0cHe
wnNuHpJ1c1S9G6ItR9VLyX7g8P19ztBnFH+zL019dWM/A7j9lLl5hNuD4JsmJBFm
rL6wyPpoibMT59EybSMbaSml2tFzA3eWtv790DRk4P2spd/0fY9YyL8uqAjNvKxX
5LlEM65Cy71MwmQqtPLW3tq7YIvdvG73B5EgskkM+bwh0/B15+i95ddujPU7yHsL
BmiCGR8yk5H0HgDF/UbthQh4hfTfNbSGVT+lhWYZT6MsBZM8zq1cEJI0b4HzMUfk
dh2ksbJhtXTWW+9sDjoYEjnZfKVMBtqPIBnkVoG96OH3C7KTK2zfvjIZSCDHYUIg
Tm3suJkr6xmtHDc59jLIRN2bbgMY5e4Z1lQ+/S2q0qlwT2zIsFhpu/ogjQXUprxw
rIooUwbECuK9X34UVdkyyhw192wjVA2uOngs3OFO28Dba8F03GNDFFTKva9LP+RV
NQDHl2SWvEG19v/TDM7cpL8kd4wsG33gUCPfToKeHzuyQgoexMEueOjknGkX3+Kp
mqDaa4n+9pokkQOrWYYog+VEIAuV8dM1+uMGdu8YoaRjRwXR/CZrcqyX1k2r3X9k
DNXlSu3SeSZAqKNoofnHJumnCnhdJIzlDrZ4LQgo7i7kY7I+iEKg3xdDoescNROb
7K3cfzbs4+28FLn/By+aul0Q7hD+2AOwYTTPJpgIzL6k3eABSynXPnhBMhU/nUww
Lxwa0v2GYPmyPOFxG2pqGspLlE0Ra6nVl7Wz/HhM7QbgCCOyrUeQ2vxSCQLKsX9Z
dBhwOrG70w/pevzw2c5vps7gWM3Cy7gAEknImwE/VdCvyJoFcgOcNexsLzwLi5iG
N1JMw6LqIvXWnr288EfekgnXcv6kZM5rKvZn9lZbXWagvwM2S2zHTLzN9m4pnwmw
OLqrgEMeDb5n2bqCqAcvwCak+d8SgMO2PgmNl/3LefXr6SXYybGZdf3ZoPshnzXE
7PemFUWmvqbsEKe1tnwnZkmpj0spFPdQWc210Un1WY4nfJAcF0tnJRnhxDwULtJD
cvQzMABNjiy4osJsnzJErsvnxr6jAvdJUZ46Zr34FRKSXq5dScw9tDbjNwuVSfSB
Kv12DfZQl7WFMDwsydVvb4KK6Jd1Xa/8o6f2QjOMc5y6zovI1zU0WprJ2VfmTj42
JU4aeFdRfr+tVG1b19nOBlMRe53BOJlMLnT4PP0qgetut21I3HtOjGBAuS6SW9m4
bLhYDEHVeISgwnZ0ZnxRk5MsVPKxLxfn10HM81xx9A4DdSRGgeHRKNh+Cy2ueIF3
LLq3H67mtd6dqURPZZtB0KPXdMOVtyF7PsNsvFRT19yI69dTpUFxGsgpQAGVdbwa
kdWXqCQsSrVvOLXLI+zV40OR5slrxH3aQsVDdaukUOffT0VH+v/9YKEr/7F//zMp
UezMLsZ9Q4Fh5gwPyc2cXgTUIZ9Djmkt64lKs12d71rEveKMve3Mhmh+hr0d8ayS
Mp/Ur4Km27QdubD/BKZqMMGy1Y0YziNcnkBC5n6aGhE4AEmQJdXrpM77gi5GsTlp
y+9CUinzSGtPiCrcy8IUkbNjQ38ITdyoaupV2j5qyU7VEAijh2T/sH9N1BdF/9pF
rJljqgYujeg94315uF0Nr/KCKP9oDow6VcFHO50kgSRYnqW3D5NUFJ1t7G1cSmEE
+wPDYvztEV+IbvSZ6DpDRb7BFsi/NxuFb+hpn2KMPBj1zAeGoHXaHuFnva80i2tV
RUHdCdsqmHBooejl2dkuZzjJSuQXtolZwxToYAln4jN3mUzHwIIPgqChsPrUZ8vL
4zE7i7gzb1E548NpgD6PgZzhz91AvpYLTqt1MwebXoXT6z1xodhZT5DZiLQBTouu
BiMHqFdrl+yZo0eVpEc288UHo78yPNw4i7bNfNeoym7lv337Pkj9cMRlQFHICOlF
riQm/iulwCga30iLOqRDHvsBW6MwjKXijX3ELpTuOMcsuX5Z3cQRvCTE9Bkr+yov
xOpkKXEbbE4979gH99bKETazJFWGq3eRjj5F/SiDcKhGTS3N3iBKll0IthKnGY4b
CILXb8xY9Zn0Jm/99BeGu7DTM7csFMApByWEs/U+lW3gxmwkvOqQgy++qwCL+jpw
E4xdbBe7oTBPvDpPtzAse7e1N2VsiVMfnpuqF6VCnM32yPTEYfwMm+bd2LInnnox
Kl3avyIRj6j6sExHVHmg9DENCe/PisN5Q9ofQkYjJDJunrSSZCS/ZbJUb2hOy99K
Lk9HSxNGODM8o8c94cJiM5DWBudgYI+GpUKed2Vp7GYgTpwWr0yLv8lhNfSAJVhN
8ORYN21gg4yNuWnucVpr7VTnufWqioetLbKySlkknqgrWZU0mIyNPwKXnc6BEbrU
9bRQe3ZbW4+rs3Eryo/0kERBnP2fqe4ZcscGoHE5w3+Nsa0q8TFCpJ16oPl0pMpy
a/JNeqqZtoXMqYf6kpcs4ourNkqjq7bjTX6NMlF5JskH50RF60Cy+XjngEiq+IjI
neuEVkueLzqmvTZpk2IldrcVNu43rhX2tsIjXGjYEMSnwV5MvlY3g7zwAafLBq7r
se28wqNhQfl9nouAj/OZ/l9KR6BvFmYbS9zn4f81GZO4Xe2q71tiOb6KM2hrHaZK
nzFzukh5k6wwBWoDC9be3kbRpHQQsu0WI+hpazW0DgEINfqC6LHG3GMCw75RmRzD
7pzMyTttYf7SdfOXDncOt0Z98gz4pHceYA+FBapApwjQZ4do6686n85+azLcpI/R
fyckE/Ok+DZn0rby0Es+LhmfNnDPv6K3K00KUoMFV6aNee3x4v4Lqcg0klFKBi17
MAjwfQ0kDr8Z2F99w+hGr3uWdQX5J8VAbecmeKo5Q6WO1KJvdsaJ/E5UglGATBpM
9y3tWl1iBraRbKqfDtqx961L1yaQ+UC9eOAobSmTJFPyjFezxCRpOPejLv/gS3WY
72AkG8C5xOUW6y1/2hJb5w/0TaypyeVABokZMnymxn4GUV3R5vlhGzicw60MF7Ly
smhM7orr5lU104+QOgo+du37VFkozGtlP1Ds9IQX0HlE/cTlSdafWa16s27be/qk
tgcDcarAYenIpY9A6uLtuKnZoKNSH0uGEpHzDBy/gwhWL2X2daM0XXOvmhn0P6wh
elIIe6yRTK6MxyetH/npKQxNPY/yiV97EDlm75o6DsUsl5zBQgOkOhEj3uHl+vAD
5vwNX/rQzkFmAuv+IpwWbIssgvEAGe+HCZOvdoP7DvYECo6/h6u6EOafesor4HFp
XufS5iIdDWa+7uuOlAYtmmSRPsRVt4GTbupSaUSbE+s1BuZLarvk1ilOXZsJquDt
rvzbugyci1NzrxlVdqheMGp4QPaYwCotH2Ls1LfhGYT22ZulBqOvIsLSG00gQQ7t
BeFC0qPrtc7duSk6JtGNMLqi3x0YaNHUgnKbB7HGF0Nvlvg0xMykzivp5laKNThq
vlVcokeww7tHrro0Pnmf2RXKVzdzd3GQNBd0FvlkwqjUqiWFSiY9J5USgZRcn44J
IbOnawkTWiydimtJZfp0ABT899gFsXZzddrR83IMJSnagzrCs6GUBck1b7Bt8Z7c
KwJZztgzibMs7dvvAQpBZKgeJg/Fxt8uJdqFbCuEzyuRkfvRB5fqoJdpPYn8wMWY
yjTZgaI1I1SmJsYyDqjovqBBjwXPMb9dXGGO+NVoJ+wq1Y5en5Q8NWmm5hRSBzN7
nIHoW3aPbNSPDJi7dexOUj2CGbBoRZJtv1uJnvSSxH7YOoyDGkvaM5HIkSeeMgua
z8uXJ3uMW6r1LQu37/aglCQiToAVyk5ya9SlVpPO/tVq1uETtfg9NF4p8gHL1t78
ylOMhSA+Y5hI6QrZkd3+MMPerQfEDxrOznX1ByfhFe7JGlA7+g6x0RUJhcHK6l3u
rTUd/kJRpSqcQhY0Rwn2wzK5DRBq5C38E3EtZrhvaWBMcAueGK1Kc3CPaRz+G+ze
uJ4cmOH4/dr1uewoZ9wgkvcLO9qrU9jIPZqZ6IDTOyveR/L8Aow0dnMMJGBtZmUu
S+lt2JTSyxl3w9e30mcMDn933TrF3wyaUl89dE4xufbUOCXF/32cnfjqeUPEeLme
qvpDrh8AlQLT2vIKZRk4kuaYai9WEOQ3pu1ok/bH/dsH8WtKgxEmfY8Th9vvjv1z
2JwmYrlXIiwcfUYK4Ii+Kx3zqgr2ko16nmNViZIuCthY1Sr8H+MmJSPJ9JmoBiE2
Z5eGwe0t+NC/ecdJIY91DkC58OGZOh6YzF9oarbQB+Z65BYMc3S+jJHNFkAYbMUG
1KOan+Wfbvq7B7q+cb/oSgnTOst1TgPa7y3AsnDPnGvGMUo3guMENwJHP2hAzzuh
RMQ7Dw8mO6Cw0J4tUItf9Y/KLMi8Wf9cnupsgR0nhaVqAc818/i0zZ/RkI9D0wOp
VkW4eQxxccx1GmKDe1XqEjgTQlPD/Z2f3ssPAo6GZIjqy9h3uBd1yYJUnTnElfvG
Ob3yuYaPs7lnwuC/rJFHU4jBV22P9Q1KWia9uWeSS2RFEWvem/hYr8flp/fPXWPK
5UzMxulATzyiuDGie3+R1B4zNZt1/h0v48F8ofyJPRhHUqDHFgv2sfsM/rLBC98o
JrGoEbBpARacKLf5EArGa6m2e/cs/XaaasMeL4Cxf/LjiUXZI01TRd+vWcZdZRkh
SgtzaywoMpxUOM/NCbfIwLcPWInBu9857dORxQomonwskvMXXa9KxK2lnU0j6PfX
MN5Sx8wEq4GNGouRvKfK5qxTk8KaC+tL9u7VQCm7vArV93lGikdqc/LDelr0w/bA
L2rvrldtiMIrho4/3bTjxP+AdJbIo8jvNt9srwSzClMCG9dvK7EEwqhA+Z9jMwFe
jN1GlY2OK6XtVDulOPyoiVqlMbkEZMOPKiPlhvzP9jpAVFGPULvBrYxUn3D2WxV2
UMMlIJrWM0ZdyN2RSFYOtI5ysFl8uMBbczd/iRNe8b7IKLq5atHb8MTC4dQ413WH
k4ntlt8x0FUx/rPyDjhHci/zmwSCQfm9cmehaskmzJM5wAZejb+ZT+/3aHmmR8AH
Dr/uevWQv2UXvDcya+Ok4BuqLd4jx4jwsjYcSGZKgYmh6t3E68UkWott9Ip4q4J7
eakslSVtcZ11d5YpJ6MliqKo2wSbSao5LK3sfVec2x4j+Sp3Hp31gmKS2suv9eZ9
qs2JdjyHfpE5jeB5FUJ+gRTNdNBDWM1TrtbxPUxP53SgjdjaLlnz3qo5nksUXyOi
djLBHgNh4OlWN2QjfYf7bukyr2ijb4hjLAxDHlt7foaOB+E3RE4tVTnNzkhVQ03h
SbTXUgK9NCWwdGg+a/xXzptyvV5brB5J3evQ/7Q8y6NYoXnP72jkvH3guGUbItPE
JW4dBp2d5FD1bDviohtJWghv9WcjeroT1yB4Fb4vU9ns3vcAoBx3MhtDb4a338yb
dGArOPUTV6WHZPwkfhki1QXj/kf9Wbs1kKdpJSJh44asVkbTdPI9aDVpJ/ZhTbgO
kcbJ7BBTklDHlhYHSw51KHxfYR8fsLE9MKg5Hvif5j1B7SRrhZY+Vadn4t8cMs7S
JOFFMkN4biwSeZI7xI+Twf5qafhLKJt2jJjitKLIpO42EvwwzD+6YchD7rZcwizN
D02a+xgLbyPaQC/fGu6lkTLDj4sCP/+h3rCif3mEC8N04GNS+/KSjCkup07Co1O6
pJq9N/luxE9gf2f52NrWJVAZPLeXYo3RvhZzN8ATNGytj5rEwQ07xU31GD+vyvE+
IkNEnqxFFFRJ1S9JAsmEagea4Rgl0Db5NM3twHbuKDd+2hMcllIagvP1ncKdS/xX
HnSjZgKmx2WsSLTvVxtYbwaT3/yTTOaNKsMvDKUnIyQhCgnk+TAPoe5mQRJEbjOO
TPdubwu72W/Rm3X+W6PAc/dzmnANamAt2agrMp4Be2BacoYMAFDFnJhJOiMgyzFG
JTj9oCk1qNr4YjP8QThr47Jp/Z/8yxHqz7ABtP5QbFqCZxQjN+FUToq2t4gNE9EG
1RQvcut8Fc7CCf85sKbRwjDA2R6cLJ1nJN7EYn3gs6T1tfEIedyGUxyrQddSP8Pn
zvyS/J4j2QEGUz3A5osVkPP+0cuVosro+9jXnQk/FYB54Sbqw7XVwDdWNenk6VDu
gWKOSEFPoZGFt/UGa5XOUlg2sEE75mPsYK6I+JT4GbKyw+rz7jd5saD89rvvFSmh
K0ZzAk7s6pKWAGGF+eglNyxUfl7j9H+cDks+tMwnud6FT33HJslyk/mxpmD9VduW
SqkmQs8o4BHPa1Kc67bzjV29Cz+PJ6kEgXFwhkkZTIav70WU/w6rWd9i3fm+N8ic
UKw3h65R2wDZiPQQRIWNjlheFxH8W7UOja8QXxaq+PtlajcodcUt2JFbnrkaV9lg
yrjkZ1hc0kKJehYmNEvqcNYNRpuCrSsoU2i2aI2fSAno+d3G0zgI0zQYBOnpRU3K
CUvFjgpXTHMVCLkGWP2BDmtZEq5DqeTFIdnJIeldxbDjDCCAtcXbPojI2qiLf0GY
IhSYKjzPRcw8GJ5zAaWBIKDsBXSkzhnTdL8kk2+YmoCBd376Vb2O/hEeE8amyHVf
mM+TZenvBoQUYH/vjENf+ZlcNLswvff1EtCtb74lldz577wNQxa8x3OaNbH3Frmi
h9mn1POW0hZsTMmWymnKc0EDX/rUsmHlUvg4aQWp1HxER92TXpzHIiEs8eg9Ialg
tif0ihllnmwFpwK/d6QD9EY7mPvv/eySxg1lRyPDZVy+dVadBJ842Tat5umQ1buG
LwAFK7trAMirxnWpeBe9O5EmDgvLFVtEk/3g9+6tpipVqI0iWg6RG1c/0OrN3NDX
aDeUXWMfEfPB5PHlziwgZ7kceGL65RGssmPgIlFBWSzGLIjKj79tt1zbSmwv6obT
Jfca/ShuQhVliaESBKvSH11U+pwCur3+9xag8sCFKAWQh2ozqWy8qGm5UAwysEf6
PiwiEkSgeGV7tqBlR4vmHnxiFsqVSxoK4DzIStGP+2Kb9J3nIi7tvDfH3u+ss49G
mvca5+EH1dPitgabu1uJWXFRWD0g+UnDG8MceVgOCKRPrZKZIrPeKPk9NWQdQ4W8
hGsjIsy0k316Lnjd3BfUmiPFJKiDKCWExYCLTqD62JffbeSZf9aXgHYaXAZKpwS5
Rto+s6MnK5g/vF5S0UWElba8lR3Ba5LtPZzK1tZJ6sP3j5jFjBI97ggp1MqZDs5v
1GokGx3zTxJV/h36ZJcQ3Pb7ZvAUmQkh3socgGD5HKNiWVLNOJZc8T9MRskbAyBn
TRtRUvQgm1a2zYGVzPERTBB/r190jz2cIRZxOdKZsaeuYkKFiV16ljKMJNBLeBmW
9bUtpenxIsy0MlP+v4dmTHY7U1Hg90d5OMqKS2LJH/WvTj93U9DsEDU8FjliYRCw
mWJW0opLPGfWfAjCBWWxBSkyJ2o3yne9Y0i1AT4T131KBuPHzUjqFes6PdVz+Dna
DoMCRdno0UYkMDEHae8NG68DIDL98QPEVG42cewipHjg6HvLeu9Vu+0roFfTsFrY
UdcqvFhwKlOvaK87kaobdnwmmmwPWaDuwTL1kF6Lw8c905srKm5qz78XODrpdH9W
D64OaIGFMH20XD0vMO0TdIESsnh5eceTguZsQYntmqLYRQHP5T72OzpH2c+9trjs
lyVisAo96HJJOjSzV7p3e6fAuZ/nys4rOrGKg3lBNlDmK9YU1/KbKQuscD3tvjYx
AtiYegmFrzdjTgcc1sMQxpOg2s4Y1S05wot0hPa2YBO0x6iV2Z5o+ofgrdf3kUVB
+xp4hjr/BUawAqlBg0sZTN+p+O+JXZJbeUge9GpACs3K1Me2pGOJs8pp4Cv031K3
3Ff7YBXYbuik2uQ2rrufZH4LbsbXQGtQeXfeeVwmHt4hY3hF+aojtwdtSCQkxUYU
ubZzSkWGCZyUaqOklpp7n2rP210bTdCjUr7OALjDu8SdwwReqU7o0SP2sMtD38DJ
j7NTv+zyp3FTSYWmQXnp52MkqVR4VDpi0gOsXXOvmtMUbB2qN1gqe2JZEHVbrZxS
NHxbnRDaQYq3SBb9wIDldxUO2yrzebrBXVegSU5QQH4Gp9LG8D11QwsgjfrlOyqm
Ukm+FoWWp5Z2/p0+di2uCWBgB8A7LRKK2+NHw5PkP2hK054L/kpQ5r5yTuvEr5wo
GT/35C891JJ948m8rIowad+GNzvV/DqvBOcXEoNo+w0wXZeimlgCaexk/0zfjz26
Ust/ZLaE+Hm4XBCeGE7S+lh4HjS2O3HzPfzZ4+chgJxdrt0DC8plpAIilkpMxhon
7UJO8WiYWGbo70c8I+7jgxzkjQykonsa8/sy5WCqKiGbXXkiZ1DERCpYy4JhAlIS
Irs6snWbOs9TalsFLQpMHo1V9DPh0LCF8sCXZgZiY9IS4SdV/NtgCIBrCeF+dyT1
sBnDWNN4IYW2LQ8E0HZ4qSOWVj7OInxEznOW2XWtwZWfZ0rpOAl4XHh5fcEMOPHb
oo6Ef1d47euJokybbrLYxJhiVVlO96b+VOKp4LZ1WIGuQqfstymBVu7sV+MEeoWn
fKSusk+o7nTvJFyZa+mCKKM8opbIY0sdt4B7dD1n6cuCSDK8W8lO7A9UcWnKWSJa
wXTLH9ibYuSl0WbZGG4F/QWGbFrl5D+HUon9YfgnRAPsjf+K+ttu+gdAHQz3osYo
hSQ9vrspdVxNr0F4vR6MHLuLLO1XFcKU/jDWNIXisi2HL01IsCMSWm0qGpspedjQ
VUiBJep5pd7UxDNdzYpz/1x5mVBQnh/cZS92pA+7FN6Rg+4D3/z1pMGl3qwK26c5
WKjSdsbu0yhZuUhgT1bHMDZ38B5STaIaS5Ps3NMjBQfp+Xpqz+QoktNYBAANcFCN
sEFtiCangT5PfpZCUzUCcBKE3nGChjgkRcwufeNUkYVrvNn1gjFzD9lu8o3cKjdy
8tHZPUXE1HUdy1cUzYIwW5LAsQ8S32GN0kHM0OKDa14QThG3IFeaYIc3dDT9Tqxy
Kgn6nZFHgxnFnB3HZWHvmqwnnw8I9Z31ht0erirV7BJxxA/rAnEnD5DToLJ9pRzL
L4fyZ7QYCsnUFMkyg5JR2/U8CSxmQlgj/CfhSRI7Oa2CvIASEACcpjGtDdby4Z96
RQDo7yoewPjuwh+mjN37DE9pL4q/6SuZ4sBcpXaPIjGHnYlaPl+jAHNsKjfplU1Z
77cz1F2b4cwLIiaLnCy9QiqsdaI9fDebc921Jy8STcLNUHoLtjkx0UBk2xoIq+c6
zBhM1ssyQs3TJC5e8eDmlSp51/Xq6ELo8lgnXsh8xkw9ci2zqqo1yVtpcF0aLJQv
n6egfOzwmEocPM7NbE9tDx0HDCnlJvhKSmPHF0d6f+y19/4ixzzIATtjw8vmGdw6
Wl2qOJNZ7flH31lbR6IBspTpz+tf/jvjbKoiOIcpYL251nWCF8SmQ1yI2jCKvyLG
BQXDs9kXYKWsegNy7Ied+6ny0N+lZVwzjGLSQnI3kDBrN1pXKjvMcgZ4s1oxofOH
kzaXe0qeV14OMGCRwuofY/+BGiJJfSLn+XuJuUlX9bpULIv97aZ7tC6MSc/UDMsX
34wpMblDxVIbcfmhCjDnR51h3kZOSUvRdSh3AhxdJiBxhxiQuYuWK0JOtxBhI1AO
nHCxuU+6xCcUlIeQfe5rj4fGtzJVrQ9AiI+uBw/huuHmLZU8wrC1iAY/HGw23WVk
/CiF1RLpFNJwGjjK4p+JKwBkvCfXAlJrUTuJLEbhzHlbRTadRbNsLxe7zRRpwXFf
LftKxO5eTJkS0jQoTDYO+ygzfyGi1x7wUu06XFSxdNn7SHsKI9ffjGzeWtUPY2iI
ALgA3cA8QbP2kcYeDNNPzbkEBhIa7mQZllXgFCHnzNHprSPeBZVJ1qbwIIKwAbhp
GdiT6bCIkA6pb3NYMcN5ONWZdWFaBcuuGNlqDLdQ9oJUF3ey64FR4PKwCb3pWL9Q
I/FP7jG1DeDlGFhFMirN4v1hOsxadRPCK1+oJIDS7peCBGsHrmvVZ1CN/NnS4Hvj
UMxtd5+O/D4SS7zrQMkJBvO0tXfwhvqM3efogFm73+u3zM5CnDybfvkxW03uMPg7
ED1U95pJp2mH2oXqlWkORRCbuVgb/C+Zf7W4ox2NDpVFzByMiiopm8B1X7JMuY0B
E2D7Gt2En8akW6fidD8ek6Hlj5AbyUh2eDdVS/uCSe8VubwVjYwHhBuKD0zz8wky
LidOnuEJXrflvEWWvoBbJKakpAFgGxMEP3xRQGTVUOxyDgULttJLa9vr/E9retAJ
6JJpdg4CtUv+NlzogGh2aAH79P+ASZbH3V/b/MARkqM1AO/fDuBpCW23ywYvqAqr
p4aksgulT3Mtew/3+50F+b905WAAoWlWS/Lp9WhNZ2ZxnRW0x/YLimtxpfKYLlCs
4iqxZjhGNkEabZFOh63hEkZpCJQHG4HgmQzIgPsPzJCGwC9uij9oc9sSlWexorpD
+vSfiRzpOtqSI81pAziOTJkCwiNjzSGq5ckxzSWY5DOIvVdW8cXRuQIvWsrNti8L
9mrUOyfPni9EgcOF3qxMgJy5+so7aFc25GEL9sw99EibSv2vytoWQvFTzZFe7QHR
h3157K6F7W+ebeW4N5qgnPAiMLomx1tureEF/lSkvQ1evWLArGlZ6wo8T0tC+oo9
aryXV9M8hmuI5tukIEj1VhMsklgqIZsy5dI2POMHWO4dlooKuO5mL0qG/R/9fYyx
LJkhRamRXsZVuZCo+8//PkLArrnQ+S0ByekpAcHMyvE5iEpnZ5aU0amqjTtY1I9Q
1QMZbRiUBMwpVvhLY8WWMzwYy3ysbnQcrLlZd0Nhbc1uwTXQUOoOM4kIPtu3ducn
cXmLa8jNtLqNQRSQU5TZezDfuNpn/Rf1bICSqYXdvXCW7CvHXfhNy7adEH1gIS2p
5gvG0sVucPtLiGhzr+7TbflVM1aK77486thRu+aseNiDD4HZ9RbsMDet4bq2iTW3
Oz1LLWqq/YtzHQEeZMd7t9gJkojsaKSlMXAKopiyQ/MCXLphH4geZEmOFhPyYm3S
18yx+2rOb/29Cff3G2z+FbBCqCDoSmN7mTqKqil50NB9ez5xAL4dWKJL7QDeHaT1
C7t0ceVtkaXz37Qe90hqtXm8G7x4V7Z3bkT25cVXxXZw2M6p31lk5Mx0qlU78v7U
zuTL+ilTLvEcZy+uwrKUq37lGOXlhfMGU2ETRhZJKP+W/GghB4/bx7x3O7TiVSak
nkX3mq+lwRkr28c1W8C6Zpaca60/qSV22WCBVScfe6RX+6pSqG9idv6yuxeubm4d
ZMlEZCJKnS5fzHCip05kRJlTL/Oj9NZgBevMDmE8ZTNBNSvQlmiqoWdim+z8RXZu
cPcYEzqk//HhXdU3WmyNfTMiirKZ1nUrhFFIy70GnnCWzUV+amN/YCGV54gGLNGh
IDt74NdsHonkofyAQTelRaeBQoEwvxbDtOT9FDgm+mk3hoWsf/xHLbvj+aTBMGBE
1XOAFzOCHMrtIMfrMY1WZvQOV7ZD9GDgd6/Ii+SYq4YOgesIhCvt9f/6Mg1ayNxK
32nQrvCD+QhImEdj9cyTZMpw9cADZ4KUqLPcCqfRyVwrf4GXrBxGgnXora5x1qUv
ZakVw0Octu/yFIOYX7ZUa7iOMJi/tthWa1sx3jsQITYHePrtG6NeysudaxaTG5y4
dhqcOAp1oGiTHVull86+e6cKUxzMNsRhd2texZTARa2eysDvKpOutv/88F+onIeY
+KqBSSKszYp4Fm7aqmoZoqcd6VsIB4rrTRVx7I6C715100PhleLpWSzyjWDS6Qk/
KInu364aptUiqU2AtA/ng+kD6zjMYH0cht9Wtb+N5OzAec5lMbzJksqwEaKDHpvU
dIcnD7Pfeb0Pmhoiyx5DkZ+ARD2cGLQglefAT0QLYhmIMVVAfp2qsq7czo/B7h73
7b2dpDwdyugYE2QTZ9zoGWTG3Ikbg9ljItdetHUUh0LIv/VnZ9UYIshy/ACV0t0W
XBoBY6wpw3nQGdpGCy+Rk2oJCUWiR6+JMX5XbngftTORWyXBSI8g/FD+B4iEPJrT
jhNoXlTRSjfu4pNM5SsCDuxPlU5bE9en81jV+HNXGe42QTQhLzktDXelLKSCandS
oFBAotjLlNCHpfRQ6apd9m5k67ytFzJwEKDHu6NYTXEzBZNWECVXcGcWnPOgrYjp
BpI+eBYLORMTxu9/N654tYI8iTA/u7UHu5YQaodrNp3UOfzyVjyRCXs7DZMwk/60
vCHfyulspnWtH6QTXoWj0mQoWd4aI8VmboWsDamMjAH03oSK+WBB3oGV24l5TuwE
OFVnsw1kgheF4TIgcFTejHKRTd4HgMHT9NsjSIYCZzyGyowAt06Ophf/RBG8FmaN
trAerGBuEwYGf98QFJRjFfq7Vga4AYoutknbEHI+ZQUYLIS44yt+lNY+w3NasSBp
fOHPiQpiBfBxMXZIIQxzVNIn2XIStp5SHyEqk4jmaSbV9VWCry8QsPwJ9deiRNIf
Egqmkc6Gf5uWBWOt9WKFEFNELHBP9NmZ3RI5fLJx+ud/7tr/hN9/NfivH542PHmJ
kgZkJkLHIzpALC8Rl0fCbHNhBPb8Eg0vgJY5Z0WaT0r0t2LeB+YJSZCs6thVObeX
gpfOqEiCg6duWvQlcmsyrXqZ8hK4i5JveeNw3ZgBUWxjMAb97w1Vk2obzX9NeqzI
wJ5Iv4I263cDeJFlyLM6B/uKoNKumy+9w5mBYGqvmC80Wc3eL/7lxAOYxL8oINwg
s0fLsdPNEeMh41Fe3sd2Rh8yBO7vJXd8k7sSwl97+CLMeqxF/CZCwye2g1I1WfQp
hM+++52uNDBVrRTEmKjR/hExgNv67I601VPvYIOvnZhpRYk1j3FEevSeGRA/Kopl
ZEUymmzGxpCao/C7w6YxR24ry2QAmj/92gyWpECJWnL87s+ucssLxExgVH1QJdG7
RLLOohd0CKebDBiECrMZM570/pxeFHUURFMtQqp/y9rEFQ7sPGdMgwChrEUbEI7q
m8wv2aD0TjJPSMkfjFS4VoT9ZRgj+zuHos+3BvKKDKMKwd5jEa/CPpszWFbpfpUl
nuwTHomHZ5iulZAjRs+z7t/kXNZNARJfCBJJujhTphgfEf589OxcjwsP7CRdaz1J
YOYHmbYAIEj9iEEuEzxMou8OG5YVCxgkioAtcIXfm7X0/heISnX/jzAf7kosRbis
a5XnKEM04I54D/goORgu1RhoddgklxRFFm2vbEZM5tFsYOH5PI/NO+NFY97VaIeE
I8YosJbgA2AIHAD03aDCCsdNPyctI8kk0o5oz7zhMfg8EZr4sYnwo//8yyZRZvBO
hga+3J9PQq9r8EL4l2sEHGD2h0VN/mmLCr/zqUzg9kklZ8+HrXj0WdP0RskFZ02L
kqmAaAjnKan+uD/pFcx9Ug5oxHFxlzaAGgo8oAIq5FREPi84F34eHQQQlg+lTsKU
imsLg1aNuINDQOz8Eyyudu7mSiRiQaUSi1B+UdZLQ8fsJaqVe/BQCgAZCDfm9KAX
N3cr30ofTv6GX3087GqQsNiOWi1Q2hBzYrcFZ3ZDJLvqDN36HsjXwEGrJasH2jGI
575m/s8zOtRAF7DnCY+ACazKX3qzw3znhKVV1ktsalOCvSpbxhWa/fsgBCIx/ALn
cIhLbdhUed7R18/xV+4CPSwkxGzKWN9uUkQxgaNKm1yZdHH/g+2HcO/+OmHY5vxF
8bQORHPX31B3aRrpT40JXmodyc5eB2cO9teWnKK7+0cqdurc/8/oDY/U1CeFyy/4
nxQzpoLK1EHyJ5uS5qamuwpAy+RTDNCAgeVzT6ITbixWLkH75vDX+Xp5uDpsjn1I
SFw2ys3PJhJPSb1/CZwWUvFwr22FlVZ8yShzFhAc4vzSeqayE1cSEtYhl0xUZpEB
yEUpM5rJG13n0KLa5oyL/Q4aWsFr/9/N5kFmYPAZ2Oy3fRHisH0nSvHlYJP0Q9x7
55Ld4M6Y2nEmwdJlzmfwDSFdEMKkEZ5rdkvlDXyRXPuWWK7Z1ITpvkUyesfk/tYW
DXzekXZ+9I9coj4AnYw7qlTmHO+BPYnpafsJFkuB6o2t9XqwcKkSTWLk5a26fhAT
OwfzadFxoTEhi5IBpoKpf3EFlasKNMakOYpSVfwRpuYmMCbBCt2ehMSFqenviyuK
hMVDQ2hQS+rBjUscOnJvBJv2mEvvYqAMq7l8VIbNaiX+Qu/KSMpv18pXTZiY4Foq
6//FML27t0TPiRJCXeelI4RDVOi4greY4XxMB3A/n42c1JqqM3hzM4MK2YZTtuCV
VUnI59aRROVBrcpCHjIY6mVOqsExzg/PFKkbnFRpo3vJEx4K9PQSxj5jTZlBE4nk
Xxl3SNGAht0z3BaJHR2UL1Vaq8hFDJDScg5jWmhwHhwfU/uKcwtZgmVS46QDQ33b
ecRICr6j3/cj639Y9vMcTJDBXyfB2OIJd4agQKuuONwjgVrBIpwACwTu0gNs6t/P
vP3eSfIsoklwnbwrX4+DzA4ArqoFv57u+EkHo0+Aw0TEEKdW4333LnT6XPJvMw1h
9IY5Dx6qfpRlygz+UECfTWEbhqdJiwiS029hH9WD8aQn8A4nUsvQ9Vi27ink28ES
wD7CNzazb2O69rgGFU6ftyQMGDrW0ser7RiVE1r6oBwvZdbrR8rOpax3wB8oH12k
c0MAej8R7VyNHdjeZ3z598027lM/mGAP73e/uxvrkoB+XngM6NhdFPzyYLaLkU4M
/RH1vqVd21GhJGPE17bK1YUGfw3kWTR+XNDpc9aiu6NcPArEV5A+PSYyz6CE4RT4
Lrr2Aq6857eZYRqxy39Igdl/Bvul/xPusvtGm5iND34OpKE9GA/EBlfWvs2cWkRT
89iUmef1BG0SScPKkzGdKMxtNnW6i+Ztq8pFi90wpMGrH076JU0flYDXDApBtlxX
7uNUEAaRvcn8dWpuW2RDfChu62IsM8yvSdonzwLKbR/rIZAuJtun0I29OvXzTeNp
8UFE3kNV3lJRZYvADHnMyBjfXUUluZjQEmLdak0HE/9v1TRyTk6Trs7yQ294s0AK
IYCXWIQuCczMXIqWGeCFfwkZd+RJj0W8tRdzt2KxG2L444a7d3t7Mbw+KpH9eDZT
cbiGlWtSBlKeuDZWuIZodll7eWsfsViffIFAzRlcCy1u4RdfvPKOfpKHuUOlv47K
G8Sr5wWCNKkZ9Q9gFj9PIVOG9H1jUN3bFt773D6pxxSRkE9WztUOvbGFw3EfLVVy
jJqCqXVgAajalMu844RnL3O0QI78y/tpNa1ZjGiA4diooeXE1mlfa7nswWQ6lRWZ
6ISEf95XCyOQJ6xTQIovbCdsFgOuWfPvZcO95q8aWC1hlFm1FpWYpUDlLTMnJQ7D
OvwAKoR8ZuOER9PvI5Hco/O4ApnffoQsCmWpkZUy/GrJ3WEvqlRzG5XVdFzbEMlj
0nDNkPDGhgeP9Pwi6avUgvi8XboCvtdRPaUzomDlvGdsM9yYFbyQa3w0Y4lB8AX1
ZTGmkDRHEhV3TFNwn1ZboujAopx33yA5qpTbi5jGXYxyccMECj8IO2kjDbyiw8k9
dMsbUbvXLXy1+i9Fx0Egej9CCE24KHNA4HdugkwDr7uSnv+Dk5pRWBMFnx8mVmg0
mLMtxUTxSupq1yLoCTsjk8BSblqgs5Y6ZTvZ86m71+p6ISQtvTMrAMhSGvP4D6s9
wLG5q2WP1U++ZW96I5qJICNqYif6Xb8Dz+kka4pQgYN89VrHV5Ty/iJMWzHIkRWb
cYpfoge2CQTFo94aBd5jSRCbDdVk5vvxPYlwG9BHDl84OQRGDiDwMMuK66+8E3Re
XLfKUWWqYg1t/GH9M5oT13UGS0tZnqfPla/TQwSdY2usiBUH2/df8ubyCJTlghrI
tjdLYGyRxNDDQV+N9vZ9x9/hhv/8XunOFFKEtFItcPEDzgNBfq4vfL0DQHwbw1OL
QUN1/L4w0F5brp6u0FW4Uo5D6EhHOevKZ0AanWqrMziD9YLTBtXj/1ni8dqQJC3f
8inE53clH7t5y9ByYZAHeRlR9uDdZI7VhG9R3SCgqcrXcY2CMBTOOVJzsFRTsfM4
cr8va6hcyl5iWwrN5GcvDAGNIIPR9RbJF65X5YAaeB+O4AMCJZA3maqkED8lgI3i
B6bPd+JZ/Oue3hHf0uknay9Tjuw/m982NrbpIORQJwEppM1hNsC2f9kQ58gESO5k
V2BsO//WCzvojjOgRrmDG0iqKYvk0OYwHN6gf52f5SmVB/xZwAsITNhcNJfqhUBS
iUDp5X/DFiwYx4t0Sm7nMP1pQfER4syRMgD+N5rQz0lvB8DtSkGs5irHboSL/aKS
nW986m/4UkXezRlvJCnjHBg+JwyK/RkmIu9mOkUyWDHO31tjQdcr+nx2oIN85B9B
3oLUgjykAxoU78bhBYl4+ELFCoEHlbWQwxuML70faym6pVhDXmFzLFhqXb71vbZS
L+3y8VeUDjbMQh2xvDVPhfLrEqVZRFkUd3KhQJBMK97o+PcvMSAbLfCPRo/lBRFR
k7hfZv8Zfr9nZvSRHHM0vSo6xZvRj7HAXTRn73PbV/0u2Whj9HegznH0fyw5ijly
UYBjFuQg8L9O/L7FMZ0oXOKuQ79C9ONFNdaaaXyDeFpJkTGulHcQd7S2zzKFwSaA
CYJXkiqJCaPlGiwlHQztVa7tLYKRWziXueyOmqBLUiGixlUEUeibWxuJOmEt6vdN
yv8wn+19jScZek4wiCPmzwa254FPhtiBlAEtwBkCAGz7r6/tK+kPbMafb5KysbN0
yACgBTN7GkSIclP/v3VFFrCl5K/TbHvqluyqmVmKosytXNq4DA/pfpXA4oc5vMWf
eQAoB5z+25Duwrp+VsCtfOApwqTLjDmIglGDnaa4JCxmMo3hlZfKD7sq5GXNu8wn
2LqeTpq7lMzUZBquTHrLy/9zto62BvT+N/pNdMCOKJBzRLMxBzY3AO7SrfXG/+nW
ZNVhlEU44DvjsS/yi3u2T6uM4hwuDMOAY4E807PuQNPS5bnIJE5jd1xgVoif0QuQ
k1omRDRHxsIiGO5A1pSs1KcCM1Hm9M/ABSZ0qZoJqdTnBqQZgp4rhynFG1W8L+Ha
25BCcptwgYrUEbxgKeaGvnhOzxcH+m3UAyVGoXs4E6/HbBQqv2hdeFSg1QlmybEn
T3T+h31z3bEUSHqKW5JVdHnKOKMYSsR/r0QXl81dfzc1VLpvTsEOApzaSZFhhoI7
y8hSms/9UStDQPPKOIRhl+mNInzERrUhwNWwhU3MphGmrOsh3+nb84JxQJduyajW
Bc9OLFKukSe/ZroR8JgGJmfvHUEPMqOC3uFjtzRhJ77i3ju3F6LrsjKELQcxNgOh
B/zha+jnfezUUYMVLgFQdzpDYlkYZahiDEvuxpJrAaWzpTXBhDcwr6fD37QlgOlp
uJrAoEcxoXd+01aE+7cfF0lsSoL3gWmzYSjLpexviHJBcrifn9H7XQpeDVtmg3SA
rapcpWdDpYk4nrg7LhUur3izn5zdwcrPzcxxRDKaMiU4rkMxfEQzt/HOFCD95/fs
qgm/HQ+gZeVpg7igY61wysCS/wbRmGh0LWZTSqMb0IHXGzPZpAC16ySvxtCj9YOy
unNzcUjdbJnk03L+xQ3MEjvJmz/pFwH5+3u86f+1PKYVBXspQc81WWQXCU33Vxwn
gbXBWblFu944OlOq3M4vhYHP22+QLbFN3ExLv4TDiMDzSbdB2Y591QTVHPOb7WiE
MeNH03NNGBExORIKbC4eGlobpMFtvAYd2bNjIIZlOubetFURTPNHlvquLcHS6TkP
T0YcAyvPGSte0JDUS09Giz45wWF6at/hGDTsR92ru/qnaIgvMw/JNaZfgEST8rJp
rGGPzVtwPsTVJ3xUM5wlCLbz9Q87U66ubp56LAC/Vb8U+aRShg6t+aeBuE8T9sKa
n9j1MROUoogHbVHtffjI0AA8yw37uUxkTFQYYJHCOoNH/3Jn6x20bBvIMmdbyPli
Sj0GeLR4Zoc6KFb5qlCto7+06dIklmKdJkQblubbQ051YaC7VDBzNvmBv3MvuQdQ
VaEo8ZoFwx0hUQf8qj8VmssqSKmzdQcGN6YRuMgC82ThcYaxHL0ya/DPjcBz+ENx
eX0R2ZCk9XglTyQx/a7L8EUSqaATloAPws/2od9UN5LSg0l9nALYr49mDs/nY4WV
7iw6JeHzlWF9n7y0L8k0npHhyvSA+NDkSNsdj+ccmbahHUu3B9l+P3ZyiXewDktP
Qq29/dgBt87XRJNst16917SmrBmQjafB9c0wEkXfTwDrlXxUJ6wpB9UyedLxARIE
1oafw6YWvA6sN/zvT3T0R6pKuKHHHDPoMJAAVcgGcDktYxRiRzCsVfchLC4ZyUlO
B7PrVvGHIIjG/UHgGyAuv0hdr+poJWKBx41EHUTv2QhgTn1osxjpCPUQL/n5Ldib
lzbUR26Vieam6Iy+Y4Kean+VnmyZCp5ZZmzpnRd8OFv7bYMqDtMT32o+MxcuFlPz
Msqfv+fOmNUxHYkw4PAjuuA8JsZOquUR4qaGl6ylxvcCGfPPd+ZcEJq6qe62JymH
Z1U3nzoQ6+UZeajlTZ32WwJZGozwyldrjq8xUpPG+X0+KdGc/msBPS8MXmOrLw9K
WkPbmG8S8oxLgVsmpYZHRuwF/MORbBZCiJJKOYBduQ178FGpafQ4hm+tGm/odw2m
yNzOAuQJ4GvIow7CjC6uxfdLetevkJq+oqGJQ+SAdNNB0txUXlM+LGSIP/ugkaz3
vULESsDwPb+QN85uXGsgRumaMQPdKLWeArjCrXjce2/a6SRX8dl3Lt3As0YC/zG1
xFr1GAqWVEeINjfwf0Pl8s0GN5xqDDK43sozkGo6TaGmbONFBGQHS6XXWYPhG7mW
+l4NJ3gmoL40MD1OHkj6VrrfUqaIHok4wZuCHpCr1pQ0Zqb5SLg83B0jVwuG+JiE
Bf0ouZIG/UL3Fsz33s34lRWwIosLKLmH90HG27JXPMYjSsOFn5TgrYj625wDMY51
YEM4K5NS7XZtfOP7n8S7Z/G5UJLtEBof7kp7yKpPj3lReRa/q4xEol9vOEaXZsWb
GeSv+XiSJdernGbz2evONm+BZFV38vluj9mJW+d9uTkuCFJPAoO9SZBgI3AeY0HF
frVT2Ye19WueuOfiDhna8ozc2bjuNaORBNvoXxddll56xKhJMHnyLN64LHrDOMDT
ONiG7WxmpPoy1530Ncrab+qFId6r8x/y6tQIdzDcAM0LONdei6Fg9+uB5jiZ+Xfo
f1MM4i2OoQWZL5ZB9Jj3CBM6tF9kt51SuwVhMFGa9IKoGt2Y4HwuQnVmTHBp9pTr
IvSZumCR9YKBhV++MtA9fcXH1MLWn2YYncmqYeE4MWpFuhgRDdGtdfqECN+uxMJM
9wpK1JJKSIp8OGmNRs7ABVI68r1+yGxcAKyJN7PMts8ThJgt0e/hVjA1wDNQmJxB
1lYL9MRyG3tOddPXwh9iNxC/J5PLgO62EfJ7c6gJ7FHuozes3r/0I0Pd4JIOhJ+Y
1V9wOPDkK3CNe3VopN5vaCnmvNoxkBErhXBEOXGd0RMhy9JRz7A9iC38JuV3sbGO
17v2Tgatmc5WPQ4OlK2bdcyNUmFfj91aVeX1ZPJBcGwO7R/mHbBA+6EScr/ZR8NU
FNqsR5DB0M9oh7o9WkGQah63ifBjiiWJERRmfba6Zdd0ywomufNN/oYzVPBylkWP
hwztFcQGvz9eLKcW+YC6gzuRaFtXqo8FLAf59ujEhVudW3l+Rp+ZjYVRHgk/uO5Q
FVLbiCQ671TvkzzpfOLwd+rNhtazd56PzprjdcNXmYnkylqoPHfucv/89KBz0DmD
pt/n6qnerbiNumhOSgKrue36Ufm3U1gqpH9PR3zpIgn5/6/RtpWWdNfMscu4zhuI
G3qr0i9e2aKUfbX03LLmnSwQRR8iDjNqERO4BLByNbqY16QV9jmmC9GM/cr+n86b
I9vhygcdMqXNKhUsZZbCV15ZrcDMuzB4zc2EAkpOdpAZ6mYtsPF61ZYPfciKy6Xl
fVd6hGTEgSGaYSYxUzw2ozznTDZnf4PKt08VQOTsHdhTsFfKqprt5pjIDB+cjbqF
5dOjo7YxrRlR9B1lKo/ru0IC34UWf6Kc/tYMTVyCNwZM7ccFT4+QUDNV387psFQD
uqjLgRTY/K5ir+naySPudsPpF/djsMEpRKP/3tl9wZ4n+vdHzMAr31E1ScNzyROF
qbxe/Mr6CulH5J2CVWuvIprix7vTI1Kqbp9NfUNjR9M1OgNEsfHqY2BjYM4ruw+u
csVN0ofMf7yrjCFBrk/oFM6l6kBOMvy7Yy2FGzOWb/nCMed7lodTsIDa4j3DSP2L
YKyyLkfWSf3ThqybQnA3KaWi40H5pw8vxdnHazz8PQI48yvADro5GbYa+wAYkgK1
g0SxkGbXv1a5/DDa+QWkO1+8XO6YyngGstWw0675VaXdJ5+iZhHWZh4TnPoHBa7e
RUBUeuV+iYNnP1AAbyY9e6kCV5C8z3Tj4phsKGvtnbtkkYLZx9oP8zSDHcuegrU2
uoaY8ZDI72KFDZXgMyTQOpBO0u4mNF14niGoNJbyISBmeFJsKVdkHeIny3GaWqrA
T8sDJRtJlTjf4nMbbRAhJ4s0C0cSFLp6130lcU1NlCqKu2CUY25plLyB59EJfJmW
dEne4ID18spxDQGu8gn6l6rRHmUnZyud6qE+B99Z1AseE5Xn5k7eh6AUJsLUS+rK
RewQe8ISaJQM9ud65dAG+pH+SAwNKJHjXIGr3dZf9zhLATDsh1L2reMe3/RKm5z1
KCQuZXs9cDjcw+QzCGfD2ANxOs8v5eg6QeVL2j7NlxkBi8JrxsfUJ9R4WXHfiIhj
NqBNxDIwjs/psALu12N6mRLd5VRsX2Pol+o3fed5GW5O8b4Uw0mhISGXTk/DRo0m
Q2L5tyrRNi2bYlvci+OtTVRNM8vk4BON3R+KkngAGzI4il+uLd6uDR26cYcSDUYD
I7FTEcN69X5JqvLZx8oAch15WgBy5Rs2ZqgcDLjROOMq01TMq/RjgBLLpLeWJOpp
Zuv15vbmrXH2xKkLWGgeS/aVK+bYhDDgidiGjQ8h8BKSlAwJrDGnHCMubRCYHypv
OEgYDmfnMzRYoCHYpQZwQcg4yUyIigCye4eXz8icAngx/hHykVdt04qTmY9fzSk5
klD6KIn3JKwd/JTi2sPZgfc5NdEpm/T73nzHGWkkCDgoC1nysAa4UsnIzW3vZVLx
WMToQVU6EhkzY7RdaapzBuAZkQ5i/bflQ6pezBUDLLl3JRkWxaBeFBipEb+5ihH1
AIajJtMlkUJ6OEm4OhhAMW5cA2dzC1k9XXKDUYAft1omESLkEqIGuvDVPyzhLzMW
8uCC4S8RdIzp9iE647a/WM0IshAIK3ODHt+qfdToUdAl07NGWoX4yPK5KhbCJ5uX
0gRfgr3KymXFPo1nInbUOPFAerVc6K/Dy02lleEIwWxKqOY0EVPIZJ5QPz1qvGPm
6J9ApcjwDxtTdKTmP9bWnCxhbKi1Ij4nL+DXhBcWM+HDmdk4C+cylwV+ZQdrhSYM
R51fRE7GDOunGAzPmabH3DxCCdn5muiHNiSgCp/hJb8kwFlcVNJAtRs1L8rn/AXR
3OWfdIAWUfPrXFN+MvZ35ET6RbSOwoD6Nz/CsdFkjCvSc7oC6ez5orbPJ1xI0x0X
mA3dGlwisKq3dPdaYTb6wCtmG+2/3iqxMStfQ3E8ojy6KQb/Hcq5fhPZcQv8ynZO
MkkiOU8v3gEXoF30F4FOA/fA8jIDYcWIw9uMTMSTqQhsC+NEdiMwdQix/A1z6a1O
ZQOxVjDWz7ftAxAdGCI8i1cC7C1eb5t9DCcjurkdCgUsCzl5YuZzpYwGdkyZ+BOu
54vm/4NW1bz4qKbHFK6DfaOOsOqnlzT5nQMk42X4JM/GAduLFN4hLd2t4bqheYx0
FNnIVlQ9ShaD4MPmqe34Sumu1LmFHy+Bzmt2nTaKeUaNnI3o2tlhwhVqtOt7ghwq
WIKkPRb+jyJzGV+LdCDXCYmy4/EJ4bfWYUcNOj3FHal2TkYrUq8bWvsf8zxjWGDS
yPpQz5L66DR1iKx7t/57+EtGT6ejADqWRODAEnxbWfOMCWt2NtRqVP3hpI+GYknc
qcjcnKXBGl4DfEHCCfQtAH6orzaJDIXx8tfodoB4WLUD9DZYjYiV5q3BK8I/lUtC
myvkXlKVePdnZ8/Pdi1USic8M5sbF2RBeLatR+JnZBISxKBTzL7B8mxzPWbFC+56
Pim0dDoUBjY4VFpBk9AQ82OwtlhSvb9Uy7n3ADQOkmJkE2YutBsHwgFpXUFF3ARU
aybFnEeMWoxc0f3ZDrg+xoxtosKzZi3bWmPMXW6ou+E8RcwlEUNfHxszeYZtP9wi
Ipxfui6zRcYANrcC6AWedE8itZ9SYW3o2pNzsGnmJB28Y+QKUKy/xTaEmwG0umnv
iGamJNlyz9g43rVCw8PNcnKvKobvnM/C2BLSu1PRgjhiBy03wMtifrosOdDn04QX
vPKoQxEIwIsRO4VJRIwt7xsqp8N2XjVZ+KJSFut2k6nH5sppOZrdLACPy4qVQGRS
6MEChb/bVDHz5QCarvRRqKfUrPwbm5aiH4xG5cV0V4xi4GonKUGPVpRHsiQZHrpV
2CI4MVSYvPGJfWvv+gxjQ8D/b2y4Cm7kAwAJtne/tZ0EcLNJYz4VJVhullQH2Qay
Pj2YIjJziBpy5DMDujyBcE5x69jTX2SUUfi3ZbctDavBDLWCbZoCXqL9EQwynQC0
e58NU+nPvOb2n4ze0J4OpshvIhfl6QXktkI2h/aTZBUthZCtTCahSDzgbEHFMzhz
NMz5rRu9/8jXQQyolDm+iWsGtjYITAUHifXe4JZ7HoLlffLvo/A5E9reDCaT5XQ0
Lw+bmmmA2pWuJiJuRw75W7m15CxuF6i8xsxemxqmzW7wpdk0lNoXvCvaip5H3dpt
OQu7t6mdbNgmAWxi4H8mBxFzBWniVsU1lUrk+JDgmyanbxUfrap+CGdvL2jM6HWQ
LW/6K1SxGRnEg07TR6mRJBYG7LcNaKjISpkCwup6qCCQooiSYYxel1lKJQo5KMHu
81OOnp6T8P9cSwl6smiPMAX5xroAS3W8evY8JepuUhlB5E5JjZqNCfsz//Mt/CQ3
irUHRJMIxF6rRRsOtxm5LuEmawOgzhjJYX9En478rw9oLAyluikEdWLGHcjQWJOt
1gjzt0abJqVxo3dXO5d1mty04S6EsSYSXcheiTspcjCF27NaRSYPyl3CBwi8OUlk
1E/sVUMPW3Fqgv2vi0PaoyYmNwADzucYwMmPC0elM8JJ+Absv68z9RFzmP2Ntoky
ITwnSRE+TgpCAJ9hfYumkD+61CybsDh82L7b+ASrXvecvSKB6vBEezTXU5WY6OvH
K+cyQT6hx7uzOwqjKH4dm6PP6PjwpbmKTiu8KjA4R9ANFhvd04TktAe8idGOkTaJ
YKy0wxOTlTmB5WASt0TclqgQPOMFRUyidb5ty9E6VsVmR971s6j8n1/ei4vb+2cp
gc0aiJI7YVClB9rOiCL+FCVFlTdCVGLYYU06wC6vRT6cJKd/U1ke/MWjV9iMwYiC
d7l0VnclVuDSkh6wwXhO5Db7o4ztFDZu8IuSh0+pXwQpceOl6Oko+VRjWHHYlr8B
qT7CVv3KUBGm1xhlutkLaiJKDiGXYoWOa1WI+yhL+JkFDeSwEV1jkXE8x02o4+p3
7iPkZIGjc1j9ookF25Dri54CLIZTwe2ayk+Ar8cfukPvnvwykxRjADz+V0WEbZYa
v+brJUguFeKhkiPwmInSz/BSqQNSvQamO41adAnU0CIVKxTXlVjyTdBioG6uquBo
zrxfVeJWjDQ0w3vOZpfKLEHNicbEQ71n2jYn/CHaGIm0j2/IcW0i33GeWnJ7Hmye
mXkITiTKgow1hfUU6VrfNUcxkoDtJXX9hWF6dwmMtX8eYdRuFb62g6WiHawzTQDu
VGPzII5EjLlrsDv/act3fdG5AE6XNk8u3aemA+uZabqsN3F5sDmG2Gq5wzG+7x8I
ZBdBnpkn7QW5jmkFS3VeqvP+Nst7PM6LbOD3uSUmR4dXTCJopoYV97cCvAlshJtd
S8qHNQByy0ct6Kkc//aTrqWC/E2GWtKrZqmaYbLqxDoFrV2ZkxvAKtJuRyCA6JHf
gZRijxQsb6GBmlk9MHeqQsFmVUJtBO+Iay6ry8e3gTSmnIErYSV4v+KZ0P/PE/T6
Wl/s6cNrFO37q8soLAbusEkfKj5CD836QRrf2BetSGNxqsOGaUIM5q6kJY3uDlGq
H1YQOm1ZXjD8p3NK2eWMUFVm9sh9Z7oUvk2sLHqk8xdO+hH1pC9wA7Mjnhb29/BR
Q/6v0/HsUfpHfVih36KLNnhyh+VyGzt/Ku9wWQtGOrNNjEcKtv8rnkc+osEIjDZA
Bc8irqTeBWJ/SjqKJWS5pgRvDXdLNZsB9T0Y+syj5q0ZWs7CpyquPBTps5ZsuvUc
TSM/PqyVouhTneMZQy8FHc6bBtjT+XI6G71b0ygQb4WyVuHk2emRJ5SLGEPFn4xC
qTqG5qXqFkNsqO6KlGvTpF9vPtRCeZMn5K3jdU1gqVuuxPI9uDkJOfkcIGgX4fTT
zvZ3ZFuXxYr8YyoX1qUMTaFaF4ZhQHfGPuHWmegYsob79Eq9F2YWGo23prDVnTGA
dZ90J5H2hhNb3KvAJOxAiXvD5NfcIDZhhbbjOREW2ty/Y+SHV+HJdTNSgFbi4Kxw
zYek3bS9Kd3CbITYxHrctHjEV5qMKYd/gvx01yC1Mj12Oun09d8M9Z/ZCtDkSkL2
Olng52GGlmo+eUq9zkGSaIXTCsivm6MNEqpbilJlfQb/DWPWritIJojJZyFOyX5U
leRg1863LyT4PIFgRYZbDKcq8JxST1QiBGfb8uWlqmMcs1tJ0OSWWkS2KZ5sIlh7
TTZGEyoTnDC76h2oLGcpZY4k3V2ZG/ULN8YKOvFiNuNadpk+gCDNi3RW1G/oT1o3
bsGFyJnDZCkj9mxYzESlUylQGnwmGigSCgF0A4Ac7NS1sJQJi45/+1QICzvsJ7Ay
+en/QfosSqBNn7pyVfwZyecIg99Fjow1HuVQQfIwFJfM6o9ctERSKQQffUOzGazA
8YfLVBIRXCxiEAf4Nkxlv/C5GW86tQWvet6cY+m0SJ043ammYQbg2t/LeCoeCbbT
BfD+L5izLdqGmn6xhAOp/EXCsnTh53qu07TEhKA5FG5N1CQu7umB67pveC3UIACr
9toaQz8S+FVmUO6v03r3NbZeBoyOETKgijyBkxmDOwi305CE5vqrc0acPqPEmpcQ
FZqk3+mWEmd44jLNan84mxGVaPrU1XS4qwyTR0fydICHsoJMfBWuhyBgM7Us5lzW
zyPXToCNIvBota9IpwwsVzKB20SotiVsC9DQSG/RcaQsDZHx++ksdDLPCIHcrMGI
avmvycg6jfYO29azxcrAafEFugC2Zm+h95rk7RANm9WFSi4LguwUie2cgz+i7k+M
NYj2JXodgYfIsu5RCXthyJbOVpOQaa7gP0A8PFOQmdyls8Ud0gwCBAgHxqisry7z
rN82E/Ekh3QJX0XUyBqA3YetjfQnBzVZO32dePk1KF/9RhVBtYsoEtPLQZM1X57q
exkb6kPi2Q4XDRtQCowRe8JeFx/NjaQ8kk45CgBmtnRw9rM0nPpNgmm3PP31Hrdb
xWakg16PRIN3BDg/8tSNZlxbUXJpYGKhu+vrPQPBoNIeAxKqeW744sL8LX0YrM7o
fUNjkFBg7MsrGMk9gg2W0lcNItsRoaKGEDAb7/SQA/B7n9DcwDcOi70zWY0PG59Z
JIt0QeKVET/xD1J0cBiWQ3V7UblhbSfnSAJ4lFONvWqG+erdm1Ke39f8BFSK1a7L
bx2OIsB3PYEl0yabm8L7OZwC+gX07XORasuYXlkOptfqqeLtghSg9qxdA5tNIvmS
YqEVQjdo21Qz0ZDdHYhogP4Mr9MjO67j2pbjvL4/mLh4RKBVC30dWKuL80/ZeRZa
TdXpywNJj13iqEBHRmgbapux+wh2zvcHyMPMxU/1Df17EZTqPRlNEAw9hqBmrH2i
NmlOoMYmswRBF9WD6eB5mxCEaWHdFGO/nqGB61Q2oXEGq60i2EMuu24wt1kAMJvV
XbCSSGvenllQrfCgWwwjkq0m0qRC/kshX7LtUAf9JRaqhGG4c7kaSrm2WyDLQpv9
tlgAsDb1fYkj7J7u5CmJGHrGIXAJa2PCQdMuATFbKZHaYzfCtjl8NxK8o2yNN90/
sv0c0RhhIDT8Tnhum15zVGoW+9S0WDW8Uu3JaYag64NAhyibe/lMpwPA9gOHvttD
8rPRUMY38jUAdMfKkOQt0CrR3ws6OQkKPqAaqSQdryByMv0gYLUVv4TlONd1CgmK
+86bixPKg1Nku6YhO0JG7iuASZioDGmbNZ2oG4fKGevbE/inDTQ4EkSOmLoICIw6
6oyycuhVe4rF6+Q4JrwFjB0raVPnkMsRozHe6B8hR9kDem+BhJYqOYfkFYW9HCYr
miYXzaimCBD6VeUJD9C+ov6885x324BYvIc4q0gU+lnG8DAcJAIDEsyj5aI69iP8
/ziF63qiybYzw55bMs7T8gyBBVaL9VI+YXPDMtcnTVaOtbNvoDuvS895VR1VmQ7Q
sXyJGIvlepOz6JMzdweiy3rxe47gFCqCWVivcUkoMgn+npttoRe/sd7GHJKVqpLO
U3hT08fCh7Y/6u2Myvuaedh/khvxFzP+kDYMNJ+cCAwQ91VFdwnCfgTD3tTeNNpe
aEUv4PySwRemAazgFRXMSjSvpGdNjjDLK4npLr5i5lZ5hR+0dJk+AYf3NHdYgA7Y
Y6dVNzzX2lKF8eCVuGliHIq0UnNhK9Spe8bMVV4YHWqV0s1mfRsOexdyQidxvmIW
RRHkMU4Y4hEa/IC/xBcBRdwcSy0ylOQDuKyDhm5bbEg8k+Wc51ehL498YMDY92g+
1oZPGG6MbP5luFDfVAs+JxOuzcIoe61TrXFYDn3X2nnB2YT70URP5brU3/5EAbZ1
7Wsbkt4KV7B48iSI/BckPX5PDAmy+X2dfMqJ72SyjgiPsx3xpbpqXSGjSyzv99Kj
zHwr6qIl741p0CmokymrVtL6NlRmjW1NnXpvaO1PKP6gxsKcVbeUW9n//aWtUBBv
9Xin1CMCPVcDohjQyUADKGIW+a17TtZLq8hPz/GaYv0XMxTv/wAKgFoJZdER7S6R
QFnMFvjbLyWA07EBWMEVNXcCNIO7pcT/7rUOlhEDFzc2dEAOsbM6f5M36zKTcy9I
LnPKO7EvfEPie+cxuhAu58xLco3orYVsLAc/KZ3o2jN0OrdgEGOY8e6CvU+QeSE5
h8qVGRnl+SGl1QhczcVLKhx4UtXny0BFLmQVTVkfFuz685s3hnjXPYS2lKuKRjgP
2ptt8EQhkbfsg9mwia5N28Qbbvlce2IMZjX0hKT69Zb1bP9TR7WWiqiAji4UWG1+
XdgzTn2tsINDHF7eBTt9HXBiEFoDLHxe2U578Y7Y+iHcg8Fv2qHbHi23EP56vp7s
wzBb4cNBcpj6E7nmM318tSX533BpiIZYiHhzJ5rQ/EQxpDHnzM0mZohUh2vQIxBk
0aY0EI36LbTgK3iX3MYCxjq9t5q1cEjyD5Xyc8qYfTftoe8uGtLE30OrPdhTjnTc
TLOPG1hh8eoWXDSgN/Y8O89HWNM3OZHCrxPqR4qvJyKD8U01qKzda4U1DaThJ8Q9
GUaKhfFAp76UF/HdI7RFIpV4DriZ3Na56h6rmgUf+Lij78t2G47ucF9fY+4C00kC
shPjmYWfslycPxA+nLtiFpEx0rkvqpxSPYrFYj6/chpckxcsXbyRpJKFRTPjFjgH
KoaEhEudQ7pmnt5m6zEfSiQ9q6kVZ8wJuc5B5S3QMx0xyC30i5rXV+UkgEVME5bo
9lolKrtomQIdO4OFfyFIOBUKlzszLgfETMP9+a1QFY4HY1fGXv1oClkVPkQ5e0Ho
v+gqwX+Vd6QQWy90bIx0W5SAybgMtZtPZFLwpWLKje2kseGtDMpMlTjFRm/MmO8V
Dmt8XeaQIu1oUAMeWoLNIazZgf4ecw0pXy8hyJs2T5uzMS4TR53RAtbDtD8KL4Cx
JselAu5k/IIZfnqwpkt0aY8lHxsA8tiV0RjEQYZHau8neZYedKD6176kZmcsM7eS
CY3vdOX5Rsv0dLj2seDB5dP40QGay7OiZEtAGA/0qVosCvrZMHhU0FyhBLh0lTSW
xAQ8BiSLv4XqFWKcKU5TY3Ggq1sy+jXFurY9f6QRMTWstSEwDRLXN0S6MXqXv8/1
qhCfm34q3QfmLSPAey1zod1gEAhKkKUMHxvMDmEQuHM5eog2g8lJW/bRBR3AmfUJ
jkJs2H2ymzYfxo9IHgnM+8V3KNbI9iSnBjGTZEdJAl3Pzcr8UnBDRaxczm/VYVsn
CpQnZJMekz4nzjg2l4wYk7C+6VCY6FxdUb3oMIthXT482TRicuFno73bucdzREXB
YQEHnv0AFvZ/x3G5aSxaaEkjqw+3x643ESAUItLtI42d3j/Xt6RLSnZbNRQI64kC
+Qr6j+IwUHjchiuo975mxSdGMZT3U5OvPa3r0VQbv/+c688LFaAC/KFrWtosvoTX
7muyJQT/jQtpFNOOy1jRmlmPmP9HurB/AReJNeMn3tQ8GUFqedJ0GYhtFl0ur6d5
1GZmmNzHJ8MEG82OtedPtHVWLWM7H3heb2MlTkzQil9DJQZrOZmIaXLdxSTkPqsx
JwrKV043RJWczyC4haA+wSV/mPJqammswx+MSH3v7sA7sZalj7OeO0XOJgL7spSS
dAXGZvLhl71b1vchyaJuayfoqmh9lU7v/F5+rsiXJZ2vcIiSlLwucESV1gxYiqIV
lznE/mxmVO26sHOZNZp1CXKTGbItl6Ek2kydGkwb/oZ3AuQAbrKJo0M5KSawnBXO
L0Xj8imk7jws6SFsN2GbVrnkNDMLcQYy93X2TwKqa9YEgUX1B1lhNdf0uFshIG1s
nQeFnrgxM933aUh+6xsPEfGaP+Aq0Q0Qm2o7/PftCad/YNd6EkfWuj5iZUv/QJ4U
wV4nvQ1f0tATbWQSZO1uRTjECIrBixmcdg8ZtaRSFSVWMIVRzCHCr1CUR7+ZBC7W
/d+0iI75CP8lMs+Lvr9xW8UjSNOuBxsYOIrGzuwNOYhTzf+RJpTIoDPT5UFxcPnR
8ZDWGOp8ZXc2SG2bDnX2ofdS6vp5gM3i/7Iz5waJ/i42iYXGWthxtfbFbaiFS6SL
DaZ5uc1ao6E1kafnJCaULH/g1JfHkbP/2FnCYqhNjA5BWpzheaYkrCUsh+Q+rvRJ
YQ9FW4dNSYMpcTmWD10e36Xv6hRtaJ2UmlRrln/KrF1dkUN1EIrClmtpLEV5hX1f
K9H+3oY2X9YbbywCMLVRg8qgkpdx2ImbwHLUJeYRN8kehqh1WerkctVRDuqKKkfQ
rKjNO3pPDUsYG4BoB9w85dawAW42VxH6hFm2Q4r6WU7sg6/ogxmrNe/YcDeb8B3P
/dOR0F2REkdYS/NXw7R5k55jWntofYHGwTwKviQ46dzbK/1wErI4ym40yJU4EC2n
t7vxcpS83nHI6YUdKAIvilASCzJWpcG2OaV07K61geivvZmLZLqJ0LdHzVNJfGcP
5bYhxXCeXIKuF6GGDFsSelLHUK37KdEQva6wWlGRSGRVuDhAPhR8UaFsbvNADgi1
BPUtZ1gFDiiRQEevRyMGg8aJjw2A11amII3Pxd4Rra/epDVrUjzULKmjkbALONIg
EPjyv9CWj0Ue4t9JvmTaz7WMFyRF0gsvww9A+n1GRJa+0U7IwnMmjB1jqL6c9UUZ
X2iaGehSIgAP45TNx9DVMe64pG7AG489GdyOR1Rx6BCbvfH1AyZnXjRfGpmXVfCA
g/+eVIc6S5G/5cUX3WcJDS24ZLKjJRQniEZ6xyOZI9IXgsiNtUvWkSp2+AWab/Xx
9eGBGzqf8qBrBV4kFDJkn1l6+n/3ardPdFlFH4o7QLXr2g7lFUaq8jV8HDJ9WB2V
YVmy2t/siHFw4/Ij84PU/BScHQIM6H13t8NEqaGYJzGzqEhxGOIS7dI7P+Svj++h
Jpz5YUICmNoP9rALHKeZub/TDqAWeCQ7jA6aC/uSSTYORXPh7pzWENM+k4d1lABa
VV2AoEQ6DaVk4VEkAuEvfGIIl7dpNJOCdFWE02uySIfM45XG3Yd1XvMEmQWhAVp8
Ac18ehJb+X7BDFQGEkT13d1bG/vh/f4rp9JO5c55/XJ2nDvRtDIPPZbAqA44rk1d
mXbTIOE8UH4m/C0drPTAuMRFp5cz6yc6Urgb/UEaB7BpJAHAeqrBTSbbUYi127Ql
Xv5nzL8CEFsC2nzas1E74CAo4q+BRzIXG/nlri5mkRMJiuT+Rq1QWogdjERlKntF
MFuLwU9XYghE8wbeIY2YLXXMoXTNp3gzD2yXzUKodtgfDhLlFn+t/83Pb55M7Tda
35rtRWGhxXtZwdzvGz0FMfDIHyDjXF59h+MRPLflSW+tYmYklo72pnxhGTumLB6l
PdjdVCVfYqAast4DNevUnp2kFVkoSSBfi4d7mXfcVfYe5dOd8lOBreePN0WpHfAk
XL7qDCdUTKPQuaqjOFSIEgg2zQQe1TvBJOsDyj4fx4F+a6rsk97j53fQ0FfFIBFx
m+FA8IHRRlXWIk7UHLWBdgWgG9MB8Y0VnsYoiyCbkvZXZjk/9JSPodXoE21GW9Q3
951kV8cYL1BXFxS2BntmXiak4ofRMwwkiYe1l4cKgxuULYx3949zn0BceulgWi89
VkHZXZtp+f7W7LSGaCgoobbFd890/uv9xUj2G1QTsetRRnkS7v3CZ2xHSG2+mJsF
1MzaxmHto7IGhDeDcmjzgJBv2i7aNoytMVlS58nbXUQGqZkBKFPJSDpnwccTe996
O2Q/N91NiRLvAm7nrUXWuaE4J+PzqH1w6/gkoNnK+5yDuneM/uQmMOEfqPW4A/jk
Li3DxVe1tQexjvdAkBnOC98UIRin9oVm6+Sv4jTX/poGgekprxafJCtGsfsNrrfR
V63/P+++YPkagP9SwzRVBLfcf7XaKFx9KaBvUGhnj3XvLPG/BaNXsCZgaiCt8kva
4vf+ON2ECiV06r7MSFheGGBHM2uAGsnJG6bX3Tl52RKhiBtIltvtIQ+msDd0U4AN
0gb8XYfvjiitrnE6dj4n+t8blL99XwHIHIsgUv/2Tuov4NRa8AIzZk+EHn9tO/Lg
6Q/bi39px1GIJ6zwKmuJeCVfTknVyVJPJVWjJva4WpCsCVXRsq8UbFYyq+MTlYrC
bCOvlfiCcJeNENTe+7AZbg4h2NS9+i1zWh00B2n7EtnWNlbxjUYGJpSnOOozqru1
zyFe7MnXf9qapl/ouQmNVJ8Ab/VcRzCHW6puYnetXRva3hNRSzMz70hPE+Aaxp4F
kYLksQCZxNO2MzplApqRcD8eRe5uj/KDPpWxrMa4JwPeJ7Hla7+4x61SHtErVKeS
V9bWgWENn/ApOcv07+0WKda6ObGJCWCwgDcBupZfNFZa3veQDjCg0n1/NIYsE3cz
rrC+fJdG+tsQw+jBnyFqeGjCO56e6R2/TXiGfLKDO+RwbiTslO1tKi6IcXXctw6G
BS250Xaequx9C6V7ujiz5AI8s+J0Gy+Gy2wq0KfNnWwwGhlP1lVLTm6WXrpD6E7d
lZqtG8g+YYZw2RLeKOB4tzCM6GlVkBN1pQxZHm/UYReHtpIXYSg5avF2cvNGG2Zb
Wc625jjzwek2QjTidJwBs15X7xKXV5r4ems+OdExH7bI+w+mUR5SztBlZSr+RvMr
c7OnMBhfevguz/X0/z5cNIjol7Nb9nbfcX5v0m2MzrYWouxxD+LTz2/MeUeRQEOR
/UxIofCFCNUhr428qOrxSJTG2yZSu7AvwdVfXhvXKefRwEaRprEZvJ86zKjdASKu
QLwZ3wA6V6nWqI8B3IhvfQixSLUqkiXrsaTmcu2754mnv5LcjwLXq9a8BQMQWQro
NxjQThigIlio9r6xISlGmXc1TItljX9AZAJ7+5/Xosez1kf6+YgFZS6WlqaGEMF0
Lniss5qycQwTs+No2qlODEsIqqF7Q0W/FMjAgqe+YB+qbI9lF3IXFYFgKClyLfhL
9O8aMN+bV+86khjEn2RAkoY6anLMFgyLQQVkYTC4quyEr0s9q8f03QAkq0dLQ/C4
kVWJQCP2lO9SfL+5plYBYd2KG/yCO6Z8sHI2qWgjAR+NGBssVNZpYs//CfOuzFZs
do47xTFTwD73ekk8ZRUDBJUCmv8pw8GTQHXSX9EMyLEjCTfDQULShUBngatzA3+R
EY0kd8F+ia/bFuIuZVZjNFoDk2S7rIvm2sdguryR5zHhQ+hchdWzz9CJkzUajeoV
MP2Mo74O31k9igR6S0sFrqgcZcikSJ5irgnGfyEMYfotkuEw8J5yACy2UGp3VJXH
ouOgJ/v+jxpa0Y11lsoYgDFZZ+5WfoDJi8NE6zX+w8y0/iwLwUK7Djo+s0J9f1Uk
3JvNcwEoW3LRG7/ucclXA+a72l5z/jDkwyYn5AaRxW/VdbjG46zibgqI6kQzkqUR
jbAWXIxIOD42c4LX+fV9Qd3I+a7yzc2f5F41sqdYjhye/BbmpLJl9wHZNK4CL36G
ygH4Efja0nHdXOKFBSHQHftwgffsMJhcHB/03O8UL3YlU4OGJNiM/pt3f/ENhy8D
FYrKJTkYqu5O8hwQK+xPZXasS+Ose3Su08o6DwCCU4AhaYbQleQ0g0I+jCnNh5LY
kPC9xlb+XmAAPcnGrtNkmo6W5Hpkb/XAxvBJQ20p5u5GJvxW6S47zcFo98RPdvvP
CnGBHIaesqHy/09cNbTuQqQ1NUsWJpnrrKzGkfTHJGVAr+FlFK5vLeOac+QvSKPO
nRXL+V2UQ0bfz+DNYr+fHE58LN1kRDy06kwy7hf+4rm45AWUc3+lXbKQi4xqqQ9O
ygu1OQbR1cmSiuK3knacOCg0cXIwWIpY7PRfddLSB5elq9MDfIQEXTnOrITKs4gd
gIGff6w7dd+k1Qz+Apw0KjMT+huRBEoCXHGXG6oWhw61HuFWpW2O1L+7WjqLZ70j
Ni6SPWGDhZqOFRsUXjylAJwxR2rDy4zKQA02SGSvEqV+PAjfdfoR8aepftm2v8UF
VUWnP4kWfS5R0Y/JJLxTatzchyoo1yqtgzUNoUBUkv8/D8LgJB4QxWE4KDoYqMAk
MWC7azl2bjdw22r+Ll3ikv57pfold8LvixrVDBAUmMgfKGgwmWuNnLH8Ex79RPp1
9+BK5cpMKqIgV/xByO2hQpnqArtzy4HN2ATry34N+ySoGjhBTgkrKY16jkfL27Nq
Qt4RCosd8oY/JbX0LvxHjPdPeNxwW0dIdo82AfDfytfcD9TvqcgMFfe+8FuY+WXT
+xjLQ1jPFSmWqGeNExBol6OOKakx/qTbf6UQZXoHxPtWhlFdCkVl5YmUIZ3tx8HJ
rpQepdkSqXXIz0QcimggICmQWWX5slYgnU3sgCkPwo2GcZP3xqo5j4G5IzEZyHw0
0L3DHLnHkZl5J6QhF9EJ8G9eAKnU2dS0mj2HiHWbKRdeZgfoO8eeFb8cvAWGQLSu
cai8dJy/nYTrQizYlpABew1p8XA1v1WRoV028M+qfA1cu36C2AyKZ/ZMgf+ni4av
9S1qWABDcUcNRZ9IdEEXIs2EUu5TaY5FWETfDw46o7DVGAKSJYdgI/NwxStflLDI
cCdIvSf5pYdFaMObfTLqxVikyO3ah/koAX5s9g1GBY12HhPz7v1fVY4WD1GCLBlp
LWRuhoP/Hp7wzDF0gWFmH4VlEcu+UYW5HFWah5tfQbU7TszlHdnOte4pJ2G6ZE+i
S78TTkcm+rf14MjXS1yC/xzTByyXS5bC/mSxMbjDWRAmeXToezWd8KYI/VvlJbTE
R/gI/X8siFOpu95Yog9Ekjwj5aEd1ukQvW+iLZROOrOjFF+T644QxQLXEPy6dOHB
F9LsNcXJCCJFts0jrYec3bX7uIrGEE/JFX6xz50XIKU/QmbbGJl3yJXY4LJLG+pp
Za2BtLk3fil6k0B6+Dt3gTcVxkvSxtRfXlkL7GJcKGYElbBOwq1mWsCXMeoSpaHn
YztXlscuBWObIKN5AZbvK4grrD8+cybJHKWvv1TQ4oBfdfQLBaO03XKUkCL1Q4z8
sel7HZeybdIV88iieLt4iZS5oSOeDdG+BOobsF/gH3gaOru5/uwIb+1OZRACE1s1
nKfAlY3S9dNMAVjdk9tQstQmg53CYq2uwmygnRcVdQhQnwj2DHlbw5ClLGhlHyW4
KCxSyOsuy+gyNpFrC7Ce7Jpmpv9eDkHgMNJBWbLxlbQoZGovf7ChjMpueMZP0xQ7
Rr5qlSxa0Jj4G5s/fxBx2o4kadC47Oxa6gDz4GetAHT5/aq7SnTlyg/2F/jKpRKP
leR4wqbS3TruvCP7eIYjoCYNwUL9br33kxo72ynt8IHN407KRTGcuukfOLKvu3wW
WybpShv6rnVwm6+bNuvVmDddEtN8rPhOtSXczXJWDWtAQnX7xyZX1ssRxdt0BIva
pZPDsP/jPIs6ES6Uv/yUKYW0reElwe0cv4YgCOjjPfRco9u4I11w2EswuNapaoUQ
zNtnpMCrq5PdP+vExRyEGbKTE3LWcOo09bF7a5PxFX1zmo/AxRdRBbFraciPP+TS
k5+pZuTBnBKL1VSVfk1aS7euC6dxrM26zP99jVBd+YjJtodCYzwtVxLk9RtxwFzW
AUtkClP+HR49JkgLWt+PLaGYWHvunxZq+vY7l+gcEmLFQT/CxkknMglBbCyjBtBr
FjxlVNeTZqv+NSqAURq7Bu/rqbt/Lzb0z+YTFBLJ5DNRl4DItU6LtTnY6/l6aTWd
neZcyOrs604CQGW2YjzWRknNCN8nAFgM64OjDAmcxy3wXNfsKdSU5Ol8uxWNPFz+
TEZohZLkrIk9vA27nxSNb97n4nBIg3KZp4VmKB5DBXnvzznP3fbndreLGogP52Ve
NYkIgnuRCSy4WkS5lIem7WZb75Ogc3d7FNul/gvUrfOWXYiZwFlxq0ylQ1OQj05h
33hLDFI4BMJoaw/rISU079cObhmIsLwciVXQZ4FtUkjkQEtNChWdwFwMWtqBoEYp
+qLGNVrrBgYYkhKCX/P1mER/AbhwfhPpm3V/U2SePbaDhX8HlxpPCCLb8AsvBLKt
a+wtyZANNMlIWRAPWClaPLhtPiRA2KmAecylmLBfuEr82ZKRhDaMzrtbcN1foJ0b
JaFeiDNO+WHyoDMz08RkhLpcFRbpYMSxwS2phei7MYHVxP+Cw1VU+mvtlLn9Qkhh
+P6I6wN9oZMalk7pdViRAExRYmmFvnO6F35WCY6iicCF4azbzK3YVyLDK2CANci2
+syIoRciDF1N/t5NYeX/8Psg6Xj3gdS9lwJe5oEBoytbJ6KXQn7RiACbCIdJzfvS
1jwNcr5YnXpx4iqGV+GjvoG8JTSz7nsCIsGX+g7C8mEKEJ2SZolcIVtX1pvVlqvW
c8XsWLPEhHur9BieLtxyCYyaLhVgXepLc3h/apoCq8tWBwLSrgSCpq0dh9xO5PDM
UJ37j/2s5I8W5ZRvqZUh/n/oqzkIZ+Xt4ggxB73MLWDokMuuUeVfsTHuuHYfi/zm
D52XtRltrTxKs7PehkgVh6wxZUY42LXtKov3B1oZOPnOC1WEvsTUOgddJu7Y53gp
waqm8vP03iZeY5lZZadkR5wcTcYoLgqZ88UyVtkS4xd/TCehHVAaKoOEzDE5ds0h
pS1cquHLuH4BVlxLq2AI7U8o1E/cNfablAxwoSKje7vFrK7V8Ae9yc+7KIv8BAIL
LdYiw3jGcNWFEf9+D8ravotCwHNnL4SR7vlwPKV8aW9Q4sEwuLz5XgFgUD4CgpFA
5AuOVu61jawYlwP5RciODjE0v4THG+16rB9vBeq0nAtkJePMg9XhWBiULtdUOhQ4
zJYRS+jX0ushy7ksdWvGga1i8lUicl8jhK2vrAocSfO1yI5sqx1xRcLplwy9qHNF
cEDKHzMBOn5b62HkaKdq9v9z9MRe24H4j5xH6pRrIVtCOlTXS16JiAs0aWRk6Oey
xKhMjo1UvXXQPOHfBk1mcdOTaidj5/AqM7+HUPMIW3bKIYY0w8Ph1CQj1V7R9yne
RSDnF1+lDgLmC4bCf0CYzdi8vPBcCmXPH0b3GMiygn8lwCOY7tfeIydjTc8fro3n
vBYqqsBeE3J7qb06bNU2ZU8NMKfxUhl/B3qaizv2JwnZH9ZOkJbossh+OBW59r2k
UzkgcxUdIBovyr1F4pF6/NpQWcp2zPfJgRRvvSg7ehNGfw5F26AJSs7eWRQor+Vo
4GK1AndzR1CfbQ9abhDHFrxxtQFuMWGMYQpEXg/lvisveiMZWsO0D+csG7twbdhI
WUO5EkF8QeDKknVxMplv3MrfKfWM85Fs/TpvkbU0vRCAF1ekqdiqTOzUSiA6Gvwm
PiR+Pr9qun6Z+abSouk1e/56ex5xH3mdefiQ5h9Dc+5woOtMycDhnvP0N0v/PGPY
0kB6/2yBhhvvFXwqWKvxYcGXaIuAM5ZzT7wyJ3aT8G77ir2cPuhsDzO76pBL1YM1
hPhW2drer6lvsuAomTuAzGeY+A9+nfshHLfQdcqpto1X7MH3oyZLs361a65Wh04/
A2Bu6B7xWUzifbUyz5o68rDreEY3+cYV1W0hGpzXqOoYwLiICZo1FSxxeuEmZEr9
himmOTTpwG0uB3CxJOzeixPzw13BnQrRG0l+/Q8Twa/M1X7X7F9CwC0y79+stPgU
MnDHo7Q8a4TvwweZ4wZSL/e5EZ0vPSUWE5IJNieZZl49gO0wmHPFb8szQYdC8ryC
HmrUecsc7iFsa31JerSlBxtzOEmY7M4/f3YBYEU6KFx6yJwo0PVu/H1ogBMaEr8M
3Mz2LdSg78S69bSHDZLtCWXvXNFFcSvD6WAjI2BuLdXDkwpapUiphbVWLPpKYXjM
0ChXbScnBi9G6nncYQMpfeqkVW5GxP06ygvPSGvbsKQAuEAPTxVYofdD+qyA+t/V
DPaL/zpcLUcilqwqSxKP6gh5SjPvvq/MKX7VdRInCXJp8rRclFVczo9avL9c17Zp
JlVGNptq58YOsQynvw2j9L8KDBYJX4n3YoKhvhmvjyoXbpS2/XCYSKhVequTJIFa
XB9k05q6DEnpJl1HmgWiNj0AxurvY5bhb4FrxPoacruiC6qFNmPmvHb427pGkjig
DeK7iix3B8tZV9yfegZh83AxTComXi+gTsy3rO1r7pNdcAk6zRMYbHpCLlU3fbXX
ZT2/CmUwAbfYUF7F/Tg/EmMfiwS0Pxy6aUAiL1D0YZ4Pmw9uzhEadr1oYxyVoD1b
Cu+2UFRwcq2D9n9JKfo/j8dzcRVRwTYBt2iEQSu2/7zgjm/Imww3kjzvO3g06aaJ
Wk+w6s+QUyu77oWrAmjfIY8H+UKUvFVL2Pf33umwWoJvUcxJl8l6FoXUIgWXpcjH
iQju50uu1rESYtgIEaVQJRYx5oLJyDHbARlctUfR7oPQ4OPizcTd8qXtiRtXutoH
0e8D7q2xxnrixRYWtGkOZ2h81e1wt/7G8pqvr4iPFHOa1kkOKIXLlcazjMjsV6if
K+BN08AxBJSewktCBYKPbiIWKrC8w3StN8EpDPxLzr0ejxix2j/+z4yZfZYsmPCV
8xZubT+vZp99BOrxCueouF3K+ivdIUq3R99Lh1ewzRLF47dNxVOn045XE1w/CCM+
Yo+W6663KS4u+lAFH2pdfSa45Ueo0XQZKY54Zh2upou21nihxvxJOPIUiUtD7RpH
811QpPsn2WdAaCetPwaJRZonl0cZ/no7lq08AgfGzFlPNF1nH6uvW4zNInu6XFDe
BJj8K2eGW8P1nOvNcmcmPucxXE6T4bhGZMz4+oXVgUcbabkfUVot+oDfBDR/d+Fq
1Cmxl3oj7P/0zEsvkipBXELVOh2ApbmPvgB3NcOyAFCAxSfLlEam4yrdKgT6cNfN
/UdT22Ftu7+FMeJk4m5kqRMWja+1RANN6INXpWWj3r6i8sY0EIYYuErf2Y/UsPzs
g8PPesTOEqvDCGIWfZuLSHkBcer3kUsZD1ijLFwx0y5WzS4wmvkY8mxqJpr33Fh0
6r6CTIN2C97K8L6k5xoFoWL5bc+OvBj6FpfQb6zeW5UMQrlytyDTtd9LKYxC39jZ
VoPQ8akVCM72AyE/b2ueG/xZSDlYbXCaTUPWgOx4QY0GQHJTY1yB9aU1bmSIe2ID
6bjWtaYHFzpo9sBaW7FdugB3i5kPU5C1kIJhGtBvf8kPDOQPXFwtxy3AL0xLuJzG
NTdvs5CoA2WgvQucyP3CD9Zxz25twI7s7h2uSKNGmbTdfz0IVN5ZNdUrrejWHxr5
yAr5bYBRNmS4+FuwSgXCoCRC3alRkpNTPFY/6XrcYyD37hN3jXP6AJnxHOh7hFo+
0sI8scKJrTiGkXT/Kqy/U4sT9+ATzYnhgIKbBkMD8am5v1nwRYuOUh/ZnY2VrgYy
JgRjgnIxlHbuO7BkUXcjEHH7BY8rEehSGmhmy9SEOJeAvolK9HC7OAyfQJkz1Tu2
wj4X6VH0YY71kTQgH6mTy83DH2033vqADBI4GrkeC8PamTadtZ2HL4Ue+K7nF6tL
SxD8mKvKGwEEX/G1WSBOuLJBNC0Zzw2HqaI4TRfPbZ9vly1wMNmGGDGHzStOsEwS
ZbG1ztn4UQ4jbAT9a5sEEy9GjNPeZXguyBzwMj6CXqroRX6JkzGEsLQgkXX0zHeq
rXipYF0rk8XZXVo/ezNlUZkNGcgDpXuIhxj9oUGvGKWjEI0oCPgkgpnlfznp67eu
Lmwd7aPHJq1ExBhZ+wbG5K/KT/sJK45v7qK2FTs9U9EKgwsCDnx3eLg0ZBZ8SX9/
jdPBsp94ep80BzSnqSiqIDlul9xNyGzvVTynSw24+BZlUCIiButP6ApCjddIHHd1
7M0bscc9WCr0JfNL8Qf8Ms64mVJU7WHrqDie/D24C00ll5rTivvxy8ysOLWXIGrL
9JC/RkeuW1KGIEip/3bCqvyFaJKTbMmORbNvZiGSbKu7KFDE7dC8ZEL1b97Du97J
EOSdG4UgeZD3IlsBdqZKobO6afqRwMSvfvOCLN8hgTWRsCv4zjXxqWY5tWWvUmA4
spmhHKfjoE9m8YNHAnqkwm9JvBuAyxeuS+r6ms/DOCrkWdfkEgypzdygDstEcnVP
zzFmeyaNZW11x/XTyziLahnlij5HRdMCBlGGgXYoXVGnW94TNWTAnFOcCoguKpDR
yaO/TZehU/UdpVLSdfLFPuWO6TwuOwnglVhq4Q5t8tcfezpmbFGIrNCVTyWWXW0N
aUZmhxEe8FvQ6bdaubCPYbbbtJrUSw/+7pdLp2ioU23HwsQXt3QXakyJ+++NmJws
E8TOvjYPd0lM3AuOAwPKFvjC41E9cgLp64zaoKpsn1jMgdKjBYOAa3o0PVmEpZX4
oEx2BSHo0buzGZUxu2R+Nx+3k5LDdhJDtxU7TtVFSM8klDbHjzHYtDboZp/y3VhL
xQ+Po6I5eTzHlaE6VIVyvfoYe4LV4KxGrqy8XTQmppO4wXhpgbGddmAPgySrtlo9
ew6Yci6DackZBhCVYXjsr3+RcHfF03yJDttHeDacq1MH9+mkBG3IJJGBugDC6LPy
owGnwrt3hNX0i8AbeMDWefYcF/ymD8tVE6ZwClx9XSL49KTTYdrmMzw/A9krDOAl
RwkOvkbpP+aatviwmfZlitSCpHljuiKMic4ePokHHAUH+yXtxKmPD8e/CaZTOLke
MFVkPTYyuLyDqUyHCN0kGfJdPxmSIRm5ihDSrJBnVJvXwExG7vTj9cUeiEsfu4ag
MOq3dqIMM0HfK8l3nNPwAt0VkDd/CP4eWdf1esNvns4z776HRDM7ypdeMf+mhFpp
iSdvL9v6zbQSKW+HACcvXSPswRCmQ5c6Jyqou5opnujaxljP+lhK6d9L/dz89W8o
hlL2M5Rtiqhm7UiOhTPrXhXISK9QOSOycjZp47FnnQs8Gzlu30DdgvZu/NeEa0ba
NegEMivbjNiH2xVroGHChLPiagXVTHKNZK69l9uCGYj+P3blE49HrzHjXHLOQdLH
AUJVxYW2k1RcrnSIRZjMEp4S6lfxiB7PeTHz3bAZGyxHdoQL0x7vQG9Y8th9ewK6
8DTPsYgJ3oldW9+H9If8J0EY5f8RbnFbbeWvvFJwrwMYzzHQYcaqzWScPX4S9CHS
IAs6w8OP19pKbrQHqyoLdl2O3j/SLbn2s8PFNlYnLddYQRP/IN5u8J2Iqupn/Yrd
lci0PVrPaoFsfju0XWjYKHEsQph7wQLsgKEIvRopA8GhMQdSUGhYO7dc5xiEmTka
qge/zoJaxSMkJLAb82IzkHxzc9Mi0KNEiqbkKYJUwv1gIZ34mIUw2Y9F5rrCWS8b
f/KG62sYDeHZKFDQo9Y5y2juaSYTrUu9hvWUeNLQeKZwgT75QhWOzcFs6sRe4uBK
Eky1CQI+N/8bHxh0znXmnfZWv7rebs9c44vBuTYKrHViE5GLdrPjgCTb7hyXerpW
rzQ2lFtwrokvzhggMAGFdUn5WRT3Ir2g75peHy6gU6WHVTbaEeWSOcc/fDyT7pgM
Q/AKvhjDzddkE0h6Qm5oGXHVgxeYVcGy77GFEIdK0BCTgLzbD9ncP6dbYfWOn9Fk
czb3uZJw7E4hJPAA4pkB83WtvH0nkvLW8ThrwfW1D3N2wrzD64RZu0f0OYUIsmxG
13AJQqIkg81kLusY/io9DjyBb7ikAFFtBRqp+HLPjqoVv7Rc2UDTG6H3HGbhFy3L
NFwjSTNHi5pBDE4dGcw5WMfEss1eVAZtDTkMVALWgwiOr9KhgNgMrWBNTQnSwdPp
zxdzcIK7TNITlplzIfJ/Ntvf7aF5J2mI/W+S4Jen7qaPJFu7F5ZyW6CdQ5jkJzzI
a8kgmRWETRCorRTWG3FFzvs+DNQ81lnrljjyVZ+4liuKtWFqxZRTfbYIUn2VVdDz
o93yQZYsjb0FM7OyrzgXNYecFoAZMks7hdXTcAnCTT6E6E8o3cxiEWCD2csYHhee
GpJhc5KxmnYLkLHLgyEkWy2QtmuythEHDi/hWN+++tXv7XM9MIdcyvhYb+j25qRy
AiETAUujwxEqeSA4NOtNk1gIuZjw7+U5uEIcPp6h2QEKvTmoEuP4671TmavEXSiE
VrJuiSBXNLTs+ARowpwL/oP7rcygvxKVBtJl0OlsJXn2njdeJMDLNZQ3589/fNXi
vSnpTVoToWBtjbEgLfcPXRDsU/YAwsWkUKeBeOsJdIpmBJp28KCdLKWAOiNpZB5Q
Qrx0pgyxhzbsQd203u8dnA7Sc7mZ/aUgEFIJatg8PMpNd5Y1NQOQxTFA2tnzSoiu
9xK3ZBWopW3Wy+W0AfNswQtbyT0yoCenbMnmf074PVtXX1yRvesq7+P9lV3xh+3f
lGnMTHbrQ9s1EL3dOfrP3SB8I0YIwOXwUCJdu0x6+e3C/B/6R4+UR6X2v0Kcbrv4
8Twrm2c4/eexJbytWeDhAHUH9Egq0mGCsXgPOrdZdIcX/4Irl5cOJz6R6sI5WSAZ
xw2lPGNwVekQi7jml9EMsRz3y3z8eFVf3VduMKFanrr2pdi/W7IjtevAGlDLwg90
hurTQK23VE+vEwoRlgv7VDD6Z4BG0FMb4QpJRENBWcguIeMRA3CIPuJpeMUf/K4t
xOCf17PFIamMZDHT+Bo9/S9QNDH8CNuE4hIxxkVoX+WVmR5FiET6T4t2rl+Wwn3I
lmdYR8skSpC9tXGqEZfm0Rvtvz0wzx0YmzJ+nTPDJEUtYrAHPHdOWIG3e7VT6tQf
nlz4Y/x0Y9JnqFVmSt7a+CqWQ861VGLVpQaSirq9Z6ject7lJFfwRDhn+eqsXJfJ
y7f+13A8dBrqiX67tw3UzvIUWK0K74tpTJoR4i0bT7HGq9tWl6dD2riUQHdh+0zE
7gwecanPuWbdribfl/kw9zVLu6P/P6M+8iLUWMsPBA2InF/ierE1sbKGfRdLxQ/g
ByvLVyPDtxLFtjUzEW2MZKK5/KhNMRESoNFmXJ9THQOddJjsDEgstqfvnzTyVy8K
/eBGvBE0f2xlkFQvRUwSpdgf7GWInN1osJiDBmX7PYurJp5d0o/WAe9SN3FIY/IT
/6nqJVLRysrOnX/3gyovi6d/xXfMQEJYuKl1/1lJB9P2JEZNHM+sgQP7ieV9k4BQ
WdBkb68V01742p9ur+x3j60huP17dYbzstJK9pVtNeyDS95t78VeeGsv8dgS3QYy
PYiEcLruIuZvOfTlJz0vhTs5oWcbRunQ5zZ/30IUgwLXR2a4OL5tN37g5V0iq/q3
ds+Y+b88BUqRUb7FBCITuRdy6ANWhKLCiwNBT9xTeRjNX51qsdYSSeXupUhsEjdS
s/jvVkOcU3mTwwXjSb4l6i+FOwFJ+/+aszYYOr4jVC81QL2QC+Xv96uQXIIcs0AK
uyMhZbNhmGglJKQiMXZgfpwBFvuOzGHcTGqnitDD4kocANcEmOLuHG8zYSm4TrSm
eM0jR4VN3l6WzxQHO7O8gRm8QpmYf1/kXLGsAzJIyJpFKhRAC4NbZgWJ1E1Hl/O+
BNM/DXgfSrRwHB7/BYl1Em1fFsGviB6OkCNTyTMYcN3afv1ISciym5L/X74/QxA/
+3KBc42QOiGXhuKEJU0cBs+Stz4a9yyyIZiRyKB5zSPZAmtHWZtmRQ3cMVawszS7
A4sBv40XSZKY8/EyTO+BrMJkjZPulnf7nq6wwdIcdkvOOtXdKJDp7V4lJRvKbGib
pLw5Wr/zvhoVADSb5L+mtsvVpZjqxGWPhPyqAmghTjU2x0M1o8uCicNI7xsUKJ5+
jb+DqZaygtV/iuH7nlJ6yWS5hCBj8DhADAWdBTDAZ9KHN05yjtTO0CDa/KONHcEo
OlJwaNNlLW7HyOgEi380iFGDdDxRzzHXsYlyqrzajZGfwVAMKXJQsW93Lw/ETjEV
YfgY9THDN/l3AK30AZ31sexAj6NbtgsRfSAmtj7/VK04mTlLysRmla8WgweSn59h
5504CLPe5fD3eFIFtlUHOoPDPGt8naoQ/qFtmDW8tt6g/WG7iIcHf+BchfpGhfQJ
ORPFjlkvNjAuQJLW6xHeSB7Dn16mXNKOCNddngv0EcXLzrCofs2bUEQ3/FZ2pBM1
ZxRUaytnAHlSWr4fNzgjname3ahcu51+Kxw2KNk9/vTTerW7yHbDoXyqoD4quyI9
CpOHQhiFy7ggzGgo0EEpTsNHn6UrIV4T26HKIVUlqiWDIkkJstibh4LJoSuFCmFS
iFJHYPzsDW5nH/OPRkJyd3ClACAgXCKx1ilazwOjixmFfC+HZhG4ZcopKgjA5QEx
ahA0eaY6bYe74G2s1L5YsYfd6Al/MYebYSEBMmcXMzpBVF86ug0OkEfodd3GCLlx
cWAHM03TULY8YHcGIc9qrGa1OaCe887bLasUblgH/C+hxzzgr4tH8XNbw4VnEs39
ki9Fee6g0OLsLVLwu3d4qnJPhdaZ4wa+13tTNajJjECIJi94Wc+kJ2ww0Kc6mKis
DyBwU6n3pDOvX3bt9toXO6ja7RWai9K7v3ZRnXYjbpiXCoNA4GJ6e2oWOBu/nnwa
EZSrkbvFqQKQPvhhdOP8rDFEEB7VGY5QYq+vu3iG1d9j9XgkSoWJnMz6SaKb0mgn
vMf9oVjdz9cLuVLX4IMh2raRmvzqYcElZIL9R7tu/cGWO65EFgwoJpLGlsnL4aEu
AI4a1GMoL3GEFasBoiNE2T/t03rtlWRHcKL2LwN01GADhWrWwhTQG/vP30V0Iio1
GZFS2FIaEM/MwP0IxG1wV5Q52Ni+kZwnYewVhFuI/NffBwpVGkr82++xWVmtwBpc
4RVQ2xkOlxeYiER51rWnsCAdcjRoAQGKc80jd3Keqq2qCciGUesAKwCe98/dDVc0
YGKj/Ai4CqfK66QUsfTl3nzBWRjpffKzsV1guBrU6RWluJPxvBkLaQ13WJpKFXts
fuCv1sFioZypnyMK35eU7FxVZENDgjI8x2FgYdN4qtDgqnJT++AtsA1z0ydcql9h
XuJBkiGGfid8XLbgqJ36V/GKtLQAPhZsfqo+vtSZRMZzn299hZU5KcgiObUPLY6F
j+6JSMT3unoN559KszY5n0It1oWsE3xfmQKnTc5Rg+PEES6b7KHl+msSEOjGS08c
AD8wvFd9cQ+lkB7CTIhnLYKctGFxbjPOLibfhMY8gSJAAFDyJrqqwRHMjlvvieLt
pP4lOmAvqo0eTkzkyBbHo8fUnUncQA3PqDk7ltrsBqpwltp7GBn76TzkGt7SdOSh
mafsNG+lxnDZYWIMcoVLqstVmGReTddtqTyEDJa2bWoYEO2yE8symjT3IhIu95GE
0jOlHS6QxjX1HBY3Gf/X/phBfQudX2mfJakPYFiZh2hCIo6E0z1/rlcAtmQwhPsM
Ym9S/6K+c7B0u80gLiHC9XhdQ25WoJQ9+TRv0rNIxFtOpVN3aCLXml4vFnqChPb9
imKu/SBPNtGUMy0DK8FjSy3vKd/dLTcfLtk0+4hKBCm91+cpOZ/rsv9nu5nXgRYP
2z72HWtyv6lGH/8KsphjpPDE5XfW5wDyEaVPkwKfsf8OOCfoO/AMpMx1i8jSGbf+
+gzjh7rNDajqXk7pVJyoI9s/MXdAIwgbWyYAs+NlHqPtm7953tsLehYletFG9x/s
l+mGDIAapPI/5B/jx4EAoZE0bKakQDeRonsNzuAbq3IQ7kTaFik+kW1Ymvp9iIJ/
vQjqbf6cxjD+oa4g+o6Zge38plX1S2psGDc/LA21C6wxzatwKRy6e6GEKik2l93c
8/m4xKLYGjCIwWMdJYXul+wM5595fFS2H55AgpG3wWDSwGuW4r4aWDqscAdAuo+P
dSjgxzbHmnud2jGNUkItwqekKaieUgd5b5ebHxnt3/BjCO7HdcYP3WvkWVncU2jO
gxLTL4ZK7g6e64QAlI1hpdzC2qqRQaXSuQIaC6Cj5NaZTONooB6Ujc2xFszZ6HiI
2EQl04HeWIorP2fpKBxQK+KaNIAnQAVs0VbleL7jXXJM/HZ7f7S5yIw7e2I/0s8i
YKLlbAcGbcLxE97OO50ruJRsDJ0n8S9Gbn/W+iijqEkiJE9PbSZ2h/Lv4jkSJPWr
ZR4W+iR6Ea6gWPdSJkf+I8M6oqXisjTkvBh5QgG5hZayFKqGO/rVEpbHYtqtb+9C
ZTiOGwvzkc22QaXGtUhBTMonYzB0M6v1OPoKf6tQD1t4kvso3K0Nnt8reHrM13h3
96UDKasQtGSsMTwNhOeNx0nIoZyGswkAsM+K+dCCcT61Y9TVuVaTomyPD5RIbWUG
s777YGX2nohH1O0dvDjNLzDUc8kEHhojJ/VCUe8Ln6IOXm8CGPmAfaRLK+1lESRJ
i68Jguc1rTm/hVxMwztwWltV8+grKLPDmGd1Mlb+mhEuGa9AK/x25YnHoUNBr6Wk
YqVHqp7kVGyjZkrbxdVp9LE9kuYk8tcamuTRsL4WsoOd0NPD9PilanVPsKdHRZcQ
uo15Esw97+k7Am5F4mL0Q+d56/qoEvf1vJDSbn0dmG4AHo1c1KiJqABxoawx039t
PYmjHdwXtNYu5mYC4+HKmhfV61Z/iIxkusbBL8iNr7F9bgVA6Mh4tyPxZOf/NeRE
AOpRM6oWv9thEzk364DQxfNsuST7weJDydkRls74lJf0AQcwJhH21wK5KmRo1NiO
pxoHgWZzivXwU3AmYZsDx5vZ6HxMVeViA27wiZ+jzgRJcDbRycp9XItcS2KBbvhB
4bLMM9kuIV0aqtndnOwJ4qjJ2YVtpdB1+adpaZ0+VT1IffYNIfFl38Hw4899qDCW
mPIgWsPoDBKVU9HGuOd3Z7JNPmuThip7zhcP9YLLj3CSidM+OZk6YSRBZrehChVE
M9qJ8BpogS/FylQVrdtedwNcCy5H/jbP6j8IHe+cPxTi2lKpTN6qwvSjnKljwPg9
FxYOjcXDYj+oCMQC4orDAdE98NGVAwp185Cbb/0BgSIvYc5G3PhhSq5Pay5e+8DF
68Hxmh42DmCixM2rfEaeYl1Ln/gm2Ei/b6d6OuSe45hPJsgWnp/8emeou2FRjaWd
qolf7ApvNlQiPifc7gFdtIkAzoqyD9uF7qI6HzaA9bTOorbDZX/As/uLRTq574N5
UQyn6iGROX5C+BuXhFW3vNs4+j1+KQ1nrFhqwcBq3FfzHAUN2+Mw55UisPlvJxbH
sAUhy0Puz2L8KdWbb13I1RnY0F7v8f6VJ9Q2cSUhCG7yqGHbF41fAr/spsrx186o
pDUfP/Ne6UAhRwTdaJvI1k4tcKTUcxHvL219qFnLP2sD2ngbRD1h7Y56SdaZZRuZ
JAuo6xuTwUOUHg9cW/P3PIyNP0N1MRzITuBwbint8FehAa/a8HcBHRI9Mv123gNK
8XQ6ADd+O91rrQ9I14iehWbNZKvP6fwjmP9VRsnFwIcQHi6SBD0MA2tdwWTz2E3M
vdnLrfnJluS5tAZjNQ5YTqq7tW/2/y6gNR5zmgIji6ownkzco8WibGTv4wRjlPU2
al5dGuHUvyAUTE1HQo4rcofGXGMl6kqqn42gx4L4vaG5Vi1Z0FW6AcDKZt3d0EcR
7TDzJm/SATqC6uWb3s4EtKPUNX8PD3A6joGRtBYwEx4JhnU89gXLROyHZANgHVM1
aFhO57x6BAqJJs8VVhE0Bv1ssHv0mp9C36so1iSCH6Zx5IIX1q4QPV2H4xFyvp5O
PO8YTXKf3p3wb+wYYQnI1FR6G4T1fUeWoiboBL4vOgleDnGhTFQcb1gQ/kd//l24
5aiODgGQaHTN7l0j2ONNRGwQ2T+p3IARjQryD/22jKO+x6sZS+N2kPIfzGJKM9dL
vmROK5RU8vDya2g27Zfe85xitVxFuuctcCdrtgkd6pOHcZ9/182CeidTMiDRFAgT
uVmhUvSoHy3E+dqi4fcl1z/9Bu5+bmyhnqLZAyQtA+gJHyk50/NjVQIj2iNIAK3Q
917y+E8QCz3w1Ac9fMY13v3bZxRRbnfcWNoYUN70QxCRx4FYsNAFo40rMAvlZ13F
q1YPW8uXBbUqGVwjvAXWEbl+PtWFH1g+F2/8bZjdrzOkZoDZ0dVXud02MIz5C6ZF
L1CgQAZXkJq+K8IPSmrdFTc665X6aduRoRsvbeM9lCV814kKnbKTqT2NbLPo/nbp
yNedTBliIMjE+srQXf5bxYNJmHyb44V8m/DAQK/wWricwUx83LnBcIMIhqzAbANg
bCJQX+5zbE0Ck1/8S9pnX2oPkj7JmEF+0+YNaQUP+ilnBAJFAYq1Dc9cqlvDryBu
bi2qw5zj3c+oGILJoml91SFe2w0a7lxnufEEwIHs1jmj2WF61RPgKL0gHDAqHt42
cI5m+ywP24TBJlGtsNX9UZXjrtgTaE8VYI0naixLNKnwYcuCYsuZuMSjQzdptYS9
JhRE0l0Ly388hj6c/xz6pHtNAX9JQ6A4G8/aO368mFnF1YsdbZ7BFviKGbXCFTlQ
mSiQ5o++F/f6yY5k9HFk5PsMf+xkYaow+OpytV7FRK/3a+VyENlTnj5O9mk2hO/D
9hFq+n7v100FetUyem2ehbLNAxProcCfYuUvLNCHFn1r9xGZ7Duu2NlpVqZcGbYS
IluyAjC7h18StLh3GrhVOKUa7EXmvEfD0jhXqd9BKOd36/s7BWzZYHQhF6VCQFIC
j/eWNhdmiPE3F33sVpPiQ1z4MUBtgOT+s+pyCIcg6AQYbRsBEVeJGh8vYwBbCdyK
eMfKs4FTf7b+emtgLuFeLX8mW3kuU9Bkf/DcnbH/TDRjh9FoRWiL45O0TtH5foge
u3MShoiRHQMfmgU/lj5fUHvxvBJPM1yFk2xs5hZktwSCDyqdYayrjqg8Zi82f+rf
B6YXJfWH3CV9K1AwL8mnqIqVDmSkEbcpgro6XTZnsUsnbJ2mLGpXCOLRlmxsRF1G
9E9jSTfGbEMiNKgIMnw2GKodNa3k7PxeDV/sJnNlie/WRBZgg7J2A8sj2WvXLdaE
pLOApJak6CDduW9/y7iKqDsiUb3TBfV+glmLw4w42ZkLNyskDQkg5AI7EVBoqxYS
CA+YNgjwfRjtkrwAbY+sB7ADJcKlU6XVeimZnH+/GzfGCmjjCxtIK4wWWdetUh8Q
oHYodHOXmxpb27Uwqz0aJ2RBD1beC1YrW2lLVgNOXi+mlKL9INpizPNa/iamudty
PyUI519VmDS+C8aXsR7RmuonnT6BAvsv/E4Kv7VTz/QUf1nBR+GnqHDZwbeZlN4j
kCdQeaTY5QX+Duk956GZ4H/piAa3tRORRtjdp1VYIF+wfbnh1fyKiU1hQkCPChRA
UWSauJr52Z+fv+IFQyCYDlTqPJjW5C4ShQBDvfkurmS/TOw9MbPk1w4T6bOjySPr
vhrfkiymr1jriwQklzSchN4jp3YWer1U1027jgfDs8k3fkgRcBhJiieIlf4LVYW5
Slh0Fvl+bE9p/W7qe+PjI+dSsRC2VNnxKFC+9BG3MteWKE3tDFjmEB+10gQMSd75
F+rP+1qX8VObwvq/yujyzxxzSZele+x2ctHC1RRU+jn756cRKrK7X3DqPCau81Ap
jcHb4ppL9kUwqxA4HMN3x0CVnjvoEF7zquhIq1kzkO7NRD1wflIVNzUgejSnjz4m
jU5NAw9Uuh1HHFkIqxA0sJ8yAZF4ywl78Q1CzkuZf6UaWmrot5Z7mfCrLb6wBn4F
WIKSJM3cwzfeDUZ91pe6UXbk3UIlnqTjbfOFu1huw4DOCkHUC1/qDRUc/o7OhCas
CgO6y1cqon2Rl5lOO1MuT3j/6WpmqOaSPxoiDdwzo5YJOASHqStn0Pqy2a4wEcrv
hhU3vxrAiRat1Shz5xpZBRTbiCNkXvO82EnDAS04yJrUiulzvcBO7gDu2gz4sxWS
KUKuxJaIow0AOZMIyuJtktigoyaRnCXjYDyfOqV+iHs66Qv2wVpakR5eR3O5BoFT
5BYSwkClG3MOvLfxCjEFxVT6py97taeOtrWjI1o/5MK39D1Ui6BoZ8eQTkucDAoj
y7ayWJEiS5R03hv9MqMr4ftdfzBFX+mhqLSDWRF7hNJAn4tSLJVUR2WRyCxzts75
FLTKgFa/YAALqQa27l/4DM29XshFJKD+3kaUIc6D+1EY/UERDRVeb6Rm8lzjgLLo
QyWM27lDBXrkCv35BechChm5DfDaDqaBDiwHXHCYzJaXdHTcENC9QZsCKbpka3BE
kgGgtdlLiWYlLm5UQ1Fn4XXohk4AULH2KQDuFGsHqakWpmbyAocLqRLBdcGkEUzc
PISRNDL1Kcf0fb19Qsib6uzz7BxB5KkY24IIT2p3jRqB24hhTY6zB7THqQPvOWku
Sgt6jRFvnWohQC9KpFtG+f6r7edZQJCE9tlb/q5Sjs6/1WYP2QkstKBoG/dMfT0O
aXs6dMZP+9p4v0k/HGEZIzp+kR/McUQoihYaIjjemH9lip/BfZtMIujDjHtK8n5T
dmBw+mK/50wSyRm4l8tc740OEOJQ4nLpyryvumIZFZ7AWT6v0xZ5qpLKK6VGewo7
NMQkZuBhre3LX78EcKhMZowelnvqv1I7ZD/sSzJ5ScTVBwDlM4z1KyciYBUhdh/k
SwF9b0IrswiwmEtiGS7pEgZIIZAQks3nJCsRc9Zs5l2N/K8st82t7g1YtjOZFRme
jUwNKbsnCpXzQWUbo7BZBXW2V97Mjr5rwGO+VPnntXtuaPna/LRUMuj9WXOdynLR
sNikF7ZkL+1IXWOspN6Z9x0aq9UH+4rS92YhXBIy5nla3olKe/CkDXBJkjqn+8lq
gOdWYIFwToTLdOzzOPEE163RmnYNPFnDiOBjunvoe4YX2lF/quNft9TsNbB2Y2iG
DSHb7Wk34Y4Xq+tuq5PGfvvqvIeaNlFHpqxfAHe/bZqkaHaLkjWs2avJR0q/+6as
d1wU0FaiWKuDeZGEhE9hrKh9oEu26cAkIGJhcP92fYY/f9KMygrUQ+whNBXSKYWP
B2nmezPv44CvC7lWSRk6tGJZYepSzyIXHf6KWu7C55+qY/OfMbArTniKlxVGepRN
6FsvpQT0z9NsyQLHn9blwx7iB0ldNdmq60mZpOYSa2MzF0GrNskuJFqOYbzxfB+M
I7w2WFRTVC2ez6ypVZ5BpEllj9LG5hT3HLK+mVsmErmbS8FNZGsBMaFhd2CjgvzH
GZ/u7v6ih2UT8IkpuVF4+92j//+55hBmIsd+MELAsyhQ+XCBSN+Fk1a5XdVeG5wd
xkCn0SJLO6FE4W6/PT8cLDYLHJf1XU3kUhrYW/PAhyYK2pUTuPMva0fxzmCAcpJk
t957MAJKBPPn36ptb3Fx5rUmTB73RBP5K++aNu5En0szbQ+tZCyqmNeYSKJycrKY
RpGLFZBTRFWRgLNr9eeOBbbPnho7qb6d6m0C1wIls+d998A4pGT46BIl7FBVEWR6
foEVLFzWSxenjIy3GlkNzakm27G8WagBVCxRLU6yZFLX6soxCprarkMootjsoAix
n8naWoG3sQHIMT9sIrLgNG005YsCvLzfjC//+9tWWovnG5G3F6l+IMHrQ17++5oi
sQ2Gzytw7HWvIH6BhotPtlJrewFeTi9LaO/qQE8vUCbLqBy+CNvULT5/wuIaaRlM
m/glhTvB7hdcdsdmvqzYtkE5yOTceT+LS7ggoz+klPDrtFNxOVmZfk8YEec/c0CS
SnWdprRDfzKznwg+IriSyT6br1u++/zUal5J0AWagwqV50f+Ts7Dv0kIkVy/S/HX
PuCH23D/goJ9QfRtPw/nWIQYAXqclD7a8cxr3L7C31KwsPSpUBMdtGYYqRcVjGSD
E9EKWZoeOeWFu+YWVTT8X+isfE9MZ43U553vJzbItsceBwmByWXLL/JxPAYf9lZi
vGIOCerdfKcx6Riz/Y+HrTvOYxIl9FXbBgIsWQoEpb3HOMF/5rGQcyXgMp94uhOC
b6EJ8+aYOVOnEh0MZr4e3G+mEUwp1QxRQRntQXNXnpHOyh7jgC98okBxy2ZSJ+0E
lklTFWLCCfEl7OI2gPPkxfklatnkrZyRz7Z3LeuCTi40EeeXAdzkrZbIGIKro5dF
/bUH+DzftOLjcViiPoDr7ucvejwPYv2PGr4qEw+cB8Cvdc2j2jKleetNcdxq34nW
3sgRGaV7P/U+mpqTSekCokYyQ+YjlflkWth9IbfU4r7AGcuh66GD3lIP0etWX0oi
ar0HJpH2k15n9CzD5HltPOuG+h0eiGsz7NT6ugXE0LzgdkEa0LH5jqrT1LTAtpSE
1OrRkxywiwJ58oO2ShXc7ZnYYLjo3hy3kCmTj7xlfnz5OMYIR+PtUtkQKMx5Awi2
AocmqBSwCb64+mV9zrNFoHheNuAYhCaUnpvWA4jqpSl6do6LkLEAMOn2bHiRJHzc
Cy3YlRzMEEX4UWROtUlIxk5oJxFkTj7IeoMuXPbkPBZXPR1gUwcb9yKlm8HKz0TI
OYEpfDvSzQp6gUE9rtHtQ8+pKue+2eI0v0gdYfUrAMHrjFODlmDAz5FwAMo/6A3j
8bGlOQRb5eYP+Pt1JmbbFfM333PjoD+8l7SnbSHRT6R18jDkd/lp+1ZR+eqK30WE
91v1gzW1mNMCGPkWl/jGLQIMKSesP8QB8eZnvnNpbPZYXMKg6NUFmtFPAKEfuIcb
ddVv3e+LS80nY9uE52CwzrINEJCBMi5x85TZ5il8uNZ3oWcTv3WQ1Aeo52UfXUHy
5fBBoF0X2SasWXS0/+IbiI9khqoSNyam+P7YRG+0OR88HA1BHcKibj9H3epoRyY3
2XnP2GhHuKE3LVjRpYiD9zYsKwC9evLHpWS4rN2qIt2CimzNh+0/hcJLf8hVRskg
tPCn00r644IL1flzMbwUQfdBjGVupW5EQNq+vqDW6hcS63B47WyDJJbrHJqoKbM/
CCuZJ+YwFhHbudC+jRm/RXFKrdYPaPCq0UuyZnwoRXkZC8yKIYUpuIKv6okRn2hL
cDvQg1NWSC7l55xGWHJCjmgGi+wWgZPo6gkr/7M44FffJbWc1KfAsBzGvSqjyCfq
UJ+2RW3BGRRytNEe0dCxWMwRmsmAn4aCPmCv2vAirN76nrfBalolDXxf2q6GrJMd
kuJfsodAlX67nUh/lhwKm/HGNFh6Mh5IzsFoUHyEq8oqEmErdY9cMgKyT2ln0AIr
ZKop6Qt0ho9V7eO4lvYXtq88cyceb9nNPQjROA3fmavwZtXd1w09uR/+HPT5e5hO
Kl3X2SB4FLqk0dvmg550aGISM7sgX3CHwp3L2VRtWtvi3XMKV7UM7flZp01fzQUc
oovYjIHwIIr8E/4jx96lUU9dJyitEG5FgRSwhSU4cXXsDXYTb/LKETEgvucej1g6
T35hXhrwa9Jzhpxe+spcxe5lyW4YSPFs5Xqu1sf9t2gmMnuPdmSGi8VHC9ibFnNO
C3ivG1nhNGk1n84L22IhuXIn1AGjHqkkeWWMp8kIGnaAqFqGC9oyP5B8yzZ+SB1m
OaCgaZFM4rpBL8cyAve4BcGbPmWlRyq7pjj5vCA5BKQpd8rklvBj5MNz3rVvrH2n
9N2J77A6LG6GeJsZSMeS9fR5r4iF2ec04BsjuBHKcBQS6CFhrm0PukmyOEu9f/2X
67NJV7QqnNutl6t2d3Q5x9eiVlw5AegxSfdsabj6dmrFbt/yaGCp5O9H38bvf1B4
OCB1pnr+ryzoJ+pxi05bnHl3Ylkgtf124DnFKda7WU8tunayRHKMAfc6yCKxeFXI
3RbFodDdgBDSE9mg54J2pYS6BQELIaTHFUBQ9sKIuG35bD/wMRh/ohp17XLqB4O5
975eCzpV4Sc4SnG/O5ceuv8r+KodGLNPBMolS8fusphOh44S0c5m6Lf+uRYs2oVG
c4Xo8OnulCJx7of80oTSniQLO+vGgfUSSgKnvA8geissjIgMsxpOXTrhA5cuGSM5
1V6zlXOAwnya2mYmba8wSyCwMc56odgWbdi/D2yE3DLikSEWLaG4yyIaUH3t98OU
hgNejITRFv00i7rwWjxXi2BF+OALf78ZtWIu7LqCNWYIAqJQ9LBiHCNoig5FqZqu
JBxHq/oFWR0Aq8CNy+gTeIim+ih7TsfU3loN+Q63Wj0lVS1KzzF7+uvxMpelDCYW
ScWh8A1nzCY83/wWPHyHefHSh8FMqRv2R1mJtM0r7qS6YAI50jIeYEL65KIFo+vb
36b1yX4wrDwPUiCae5UrKthjq5Ftq2VbDuA7yRe0uaPiJMH8Swfsgt/ljIIjSNhS
hwptSV3vCBpxOjXzGaV9rnYmHaymECCBCq7//E5FPBqWTipGkzKhGGRk8sLBVv9G
4UOQdYGioxA427ewRrDgBjIBdNIa5yiPn47wYOPS2N2WjxS+e6OegwXcYCh9OIQB
NtTWCLj/nNmtodVMiANaIQkb3AJ8JJSZkYMnShy4s/I2HDFX+nqpQY9lZBq2Iexa
lZASSvrNGQsCDW5cyRO5hQP7ePGi/YPTwIS6Eh2WgJWoFgiuQkSS/7O5ot++fDYV
O1IK4VdtgxtDNYWp1gqKKtylYr3BfFqObDELrxqCDKu1PjiTOdWxQrS7GreeefCu
2S67CVa6B+3eZJXJi/8GzRrnyaml9FNsSqIHY/LMuXiGNPLAzf1lXfW5zdozkCSL
V2dw/aRFxSxCqVdFHeUyPMCsuInlNAiC3JA+tBjWzcOa7WLI6Q9447IH/OJVQNf+
uf2G8QEEweqeXQEOL1uWpsr0guRusi4NtDe/gN/+PVUhWz4WHsiS96uR9g+UKm7s
Zhg/6CucVYZJ1pdSK/rnKD6Tyhghm+SH4qeI17z7Dbq7NxfA4VWc1t4qSeunHAjC
KNyXwyCd2QbgLmi9kUNqD04PN3EE46fNIyT5U3BMpQKn2k2pjbZgTTvmC9USIl3W
6f3QrrrqR+xzqG1CaUUoxq2LGtu7OQ/cF3kF37pBXvZt7AgJm9Si/NL3J4BWmhAi
rDPaVgYwW0JZ84kXuiUXvk8c+B88rAcBWWqwcA5dM35TG4VduXEReLt5VXLthYAz
+VHwYg0QOhkX6GYo7NubPWUSbRODbPqdztPTfkGNlO+E+6T4khDc5qRVS5T8gdmi
RBZnoagB28JZQIxDAFLQ72mt+BQRdr9yszNxp5HsvGQh0PFcrBwLu/4T8Zh5IfdN
faX3Gfu5lZFp8NgKQLuVUyI9r6fYXzMAeY6Ksm1cQgmgLfzt1ihvNiYqYu8xPVqz
O6ShDODP2gy9rLoIc9gklaJbiBauwRMAvDupfo42idY8dIHZALqT5BcGUIr+yf3t
ZAVT40pyMwoHDUt7IibI86ZUWlm1ZyvCdqSjYsCckCbdjDCFyRiYiDiHqFu20ZAL
PYEhBTa46GifbN6EyNqvngNRx94iBeGaIpuOK8Ipop/YkO5nyZtBlSSvAnz6ORZy
S7gT30/B7ekDoQQ6UXE9eyDpBiG+97RfcrXttYZVrNJZ8+VRPV7Il79EbW6ReJyY
WTjWGKVNjK9f05f8hjE5+3UiPL0V1LEVZoXAX8QHBM+w6hoHJeRE9Usp1PEkyjS1
5ADP7EUnDjgt/CewM5kHB19/GoA0VXhUpSjoDGHtxJTVZ92TP33he1dxLYg13U9t
sft2NZ3bvGUzYN85ZpiKGCbl2TaI/DaTxEWf877ckOS05s44pxghH7iYD2NulWBB
6sRkbGXDpcTfyhdm3hYdRBL8wCV7ryPC5dr6gnDK1T5FrR+QkOiGrERtAuXHGsed
MI9i3wASQ+yc5XVFHSwwghc3nE4PN+08BE8E7gzqG3m/27oUivOiK99/s4el32dP
r2WQSQXXqplCAgoalaJjQ/OljfDCYT6qe+QId1ukteUKvpaKcef0PVJ1FX0t7p8B
6S4ox8LHpw0furKx+zB6sS8juBSpTCYm7LUItM3K904FyXbpK9dfq8jwswSMiwMe
Di+ZpJXdNrzZlxiILUsKiZuCnNTEzkoX3TK671R8l1EIOxG4nj5Q0eFmLlQATijv
LVfJJMt90++tuWRPPjM1XsthSsHjUHwhytpbnS+2bCVx4GdeG6qakJcXqXchg58L
0FWl7yCUtl2jzECvNivsBlyTIsVfofYd7KpiNS7gI3PCcziRsTRjYI9mpuS7J8f3
laGUSBZ80MZxK5C51h8SQ+WlllENXC0/ViMaAo6u5vhqQPuqk/kwyZSajtIVdP+7
IFxWo01JrCRYccNSmyN0N247HWUtU2pYxRPFX70K4bpGDpZl6iF5/zlFFLooNfxI
HC+SVAiDcFks54ES4v0BmUqn4M1i1zRZLDAwZvaM32jyxwRyNCIDqpZ1uXc0UgdC
RvqSTELj6+JkkyoH1WGHfQPoB1iY/0c5JqiP2XQStPTV9IzjqgT2BdXYEwKR6+i3
y9sbtdPEkDT78DZ1YajgWN6W8VB5RuF9UGDJ6KtRVc/ZSZHsI9VEbMfGbQdX3OyD
HMO1SgI/iq0SneoSI2uhsFvjh7iNa7QcwJ4vrKg+r7k8ioChNh8oa2tyRgX25b6U
NbDdaEgpS+hsVSshvI+keb8YNqk0tdiKfOmEdJZbToqXQBb1s1lUrYyyFk5FtcmF
8z1ndLA5Bag0+03/mtoQnuE2paPm3e/Oo2NwB3x7sZaQvTrMZqMyg274NpEoc/Py
00FZlsf3olL0y/o+fVB+kIYNlBLFDdh8AfvdwyEG2c9Ox+1Vmtw5fa18ENvG1v+r
3ptTIn8Stsn6ah4FuZ/M2CBic7OskhEiFBXYT7aHbLYpkfsiM6OosBpZKMBOEeCF
9pbU4TnOkY+XQbF8pxVLiipEC5FWvGp34kAEIWvGsbO+PVnoGnE9LfQ2f9OIvdLS
QsQw4XYblbaTUxboL7w2cw9Ea0oY+juq4T8rA+KIV4bIY4NRReAZ3Y4nmT6H5dmf
G+AlzwIrJ6JWAHMeNNAYKkiaytg5GUnqKr7gKA5icho7qWptWLOBthGhOaagQ8tY
glJLTDsFKglvbxPnAGZDHP1uNEtbv5g+q5VZjYYxHrEWMYSZUOJpXxUhjDLADmFu
C4TiFYnoD53/fuZqAx+Xzz2s/PH91oo1lj2BQh6U7Iqi5SUP8rAa+aq2fqUeQL8s
msNyjzHVrXFugrCGvX+hSNfh6zCmKIvT3yB5ZLevcGja4MSC3ELb/h1AwmLNNBzb
LqnSl7OrqtkvAQ/8z9I6PgtH6S04aEVBZV9oqRlz+Mg54yd8cUoQ+oQtgF0+NEOF
J/UmmQOFXkJrR3cOFtmBwaYqeJQXcYRuEosdejQ9lyKNDC7nRYbDbNPxU0hadlmz
978ZzaSf18zQUT3DgR5G8BA0b8M5YL9PqrOe4sF61y9rX/aer5N1Itaqk7C7kQkm
Hyyz/fHbByEW0d85Hqd9kn1b3OfKFWQ7zDk0w0r2wdNhJSco4wsWOOl0kvke6+A7
0zLZI9RXBQEn2gaVTT0wParCnRYi+jTrxJNlEh0DBT97X62i9OESWhcrV68ndgzz
4KxKMxAZwzK8z5bGTzH3erzja+fj4Vx6weSV5VHeVIGZhkNHmnXH2zkPkfagjVxk
47Uaq3UnWWvNwtCnE2SRt0MP5xKP+mecb4PYTIZ0aj41hwCwtn3FPMFL7xk2Yacs
qo6+HIJYNU1mDxnOICyKxuzNhXwQI7xC4sxiN3z4/6X+f7wjmlV0LXOY0mgWDkMB
AfMYA+11wG0vpjCKXbxuyN9/IVXGN0a2XiQ9m3IP6b/TniMlu+I0f8WkLh4sxWph
IVEHPwYVmtvF7dUc7F2TgE6j/Aa5/N+G0cDZYycDmj4FcoC+JIdkEQjtVIEMcfA6
cCEqma3PMHWO41RsxccSlLB3OJhwpcg8SFDWd8/L6Cwxv4FxGpAAJp6F7neo0nVs
mDeftylwlh2j1r3a3NU5AyEdsEIUAAE9P+2KPGkWnpRFlRKBax9o4w63HYJiQR5h
dQrseaajHxDl1pbyEILuiJ+Ksg4kJV3BIGzHX9Dm/o2HJrg1AyYZIjO0YCCygwIt
NM3AAUp1GdMV67a8AQGu+2Xas0MyLNEpAP9xZbg7N0ev+CHfQr9DlkUhVZ2+RPKB
1o2FWy92+8Xd05UO1uTj6rgMQizrS6N6nclxQPfqWfi6DLGC3v0VgA7HyldVQ2Rn
nUiNiJauesU50d2Q8TR3P7E0Fzw6lPDcRyljKWy7vkItJevk1/KO+nMoPfvY89tU
CsnbHqM6TTQlI+JsMQ3y7YR8kcXCXlEKr9PmrTWU6kEEkP6rS2Dfo1aOheG5yuuS
2xCOTHbk59Mt7IellfF9eQtPvtHn76w8uj0j5wufDcWOudLBGbV5DnlPyFvrpNKq
gijBdETrvG4EkQMfdo0SoXVevRNE9vosmH9t/wYK32XDkXQcOUIqwoWHTe4FZAsy
05D3vSond0vChux5wNd1keo7LAq08cFHw/N8+XOKpdWY5vHlFktmu+5oCjoQQelU
GexsIrz8zBCu17/o5BOTO9HSRx87y9ntqe+UmEdWazHQ1EkPGRgKSMV2WM8PEq+E
/VEQlE3pl11o7vdo9KEooDpxjp6zLUeIk75QhfcI9zxHRmU1ne6BuO49NI6ILei8
NADudoDBZXdMn0iibjH4RG4TcQ9DyZz5EYJU5w71Yki2EPbhB9LwvuKdCCz5gCks
t7a0DQgYU5PXLTS/ZX/almE0tzi6YFOAPRmf5UHNaCSH3daF0wNokng/b4FBKnqB
uxhPXzSzxnMmxmHsXIWUUPDYmrsKbylIl3OnKzwYSJK2I33gXgclfD5uh7iadP1Q
D2Epu1/LwvLAHcpcJ5YyiqDWofw5EfQ1t/giyx0WqzslQ1Y9ns61ji94McGVsChe
11T24ZPSXwCD6KukIaoxPhp79EfduNef80ZvePKbg56hhRQpEPOQUHGAR6nudIHz
nxGwfe7jvslwIYQhWVsZFqiZ2ntx9uom/Pbx47hTi9/YnuUbFDjKazMvtE5nxqfD
FND6je49UoQP5GLW9VY4GDKDEudutf16ClbQhTO4jd8owXKax0bef3M0KzoUkwZg
O/DdjF1lTK2qsgs2xGT9OmCZpyVdrMUcza9e1Qx53YbEZXsbmIZR8zPHpdujVayG
BxNnNXAUm0Kis0YJ37dUlYxhU/SdPuW6Oagcgm7BSvjnaYjDZrEeiL0JLvXDKTae
A3Y3/uo57wXDJntijs6d2ggTVTHyBRYywTzo8YV0vmAKESspMymW2KnuwXjfUE0W
du/jAtx9UdYfdgvUdgfULHPNxJf6gFEzvKMHRNzzDDQCdYyR6TNaNDq2O2dWQ8qc
MTm7cm4XGj+AjCzUKpHL37vm1SSUXY2NXXI9GR+la9eK3lE5hbH9ulx8l0Dt3Oew
hAy19DmvwbGcmqyO7irzDc89wbnK6uJwlLPyZOM4uVaBF7BVlQAcM7FwAl2ZoNWT
SsoCbyUFTAAGKGVHqTwYN6mr/FO20+QIiMIkTjJsvHMNpOdZ8HPgPnIbjzHyzUHc
Q2Gh5H3rclm5QTpZImSEVhcTkVtdMfOa7vHrceaoLZMpCUWwZN8x7ypKcjPvGjKH
OSk6p23YS+v1qmjmpOM6m7vQNNZDZt/Df49xjORG95gvf02dVKIGuKQ2EVMiE0ta
/k4uKnDS1dIOkIgb9E2KXTRHs2DGQ49Q8qoSEsNkYRQH6RgYarnnZ80336uMho+N
DWiMG2GHrakjpgvRhabYX/n2FOQz5vsvMktNEES1c6IcWpJCQC0A9f3LnF1yTQow
S81J0E0OnpBhClbJLyXTNhoNTS9Rr+yktkLXh+NXxFg1kf/p1rYMSwAk/aUVb2IK
j9bHdg+oUf9tCXnqkUgK/OSa1NnXKnvEJNY9rXxmFg8phgJmcAJAIW8vxvnEPgSY
unpeTfyXb3bUbxYyTBlt2Xcbr7U3j5zBUr6lfh6pWWOKcpH+s/gL0iJx5wRKAiIH
5uFHFo/iWw103G8RcCvBSiWBq8lrmqHpGZpz9Q7RkQKSzbH8Gq0HEkEVsnH+aJXZ
rxAinIRALK9Fp/B+N6GlUmiRpDfKeKJLcets98tXqdu5widg4r4Jaisut+wttDKu
wJeZNXLrCpm3/4CZCqzTlrJ3KTAt2vLsqkhpXv+yYxfovLus09e7Lm8ZvIduD2+g
kKtBcXZKCEsG8djJyFX3jFlz2WjJws7tKSex5K6WFARVA0NHnUtWNa6yB6RbEGWL
lhTlLgeltTGLJnexY7JNo87H48rL/1kxgsDO4Bx/1ewLpjVHpZmOD8j2dv8PiTtJ
2Brn4mJ1vHqOOnGUym74wL208pxtwFtbVqk/pjW2jRXDEGNvo2OFAstVP7z+ypsJ
bgJ8/aiQZB420qeMWlvI9gCbhUYRS1Mp7qL3ffEbXKKapCchfP/OITUhUw4Sq/Jy
cvEQZzb2DzpEvSCsvZwjhlw99pfRpWuW7aWilCRM57s707HKGgSjMdy9ZKBGbEP/
RvmoM4mU53apmZ3cekbMjOMp1UanJzvDqdDAc46HmZfuTPWB7dfEs47ALSgZ193k
31ki6U3i31VB7yBecN5jbMkB57lWVYTQ7vOmJrNONhknybc+MlDlK1DgQ5bqx1Z8
y02K96kusb0oRLuixXZ4LG5ix1hzcOcvfr4o3JYM0+FOwzQgNbULbsbGsiuIPZJQ
2FbXSLGNKCQnOrI+ObwYd8YicXuXaOxIVUif82A48Zlbod9XFw2vKiq1iopstnS0
IsA+Zl1qvsCyHHypg4iOUcnXND3zikFK39S1wcqp2G22D0lPdEz0pIJluTPhtRgG
6bGTV4YhZxmOSMBq55La7MqeXt/Ypo3aEOCXWQYf3EE1+Wy59LrUQHzZ9KwpGZRs
oqbefPyZXPDZhd7CZs6+X7MmSF5STGIrc54cABi2nP+VgLETtqEs0s2XbBBH17cQ
Ro4xs04IB9mKhyO1YVVGQ8ewjoMa/Q303hfKmuMmQOUV7upTNvSaTI3/ybNpJMZV
+FDiLnVBA3MUyLddAa2NcLAvWfBVa70YjpHrgVtuXZ8210FBlPHy9BRpjruBgsoI
H/IeWHAzMQYJmfi8nPFAcSb4Gn75swuayi1GprrXxODFCW8eD2x4sEtUi9T8w1A2
BPUvbAhEK0tTDVuTjySoPqUd06PIOIA9PIIw2tUrmoLLR3aEK5+bA2uDmfkUM9vf
Wh8hwYknfAzzLPAK4tUcHmEIhWbRMTYZnwEDPZyYyq7/y7S3Kc02CkRSBg8xjubE
oLH9+a93+VQmgY/0nGfS5wFsCBVvdQrWJaGNEledD9gK024pWVP7uM5LuMQPWRJ8
2PdsT+ClGfcWdFX7/5Cw27wONM/tD2YxnqKlJMKwn9nOuiE77GSWcxXPaY6+snWM
KXsDfJIBqy4mcg7GY17LaUoIf4vsstonr7Jy8PaAEw5lcf/zVcEmAJL9ytLnjQVB
a9jhkQlCKn9gAQT3GxAc4yg/0Y2B4WgcXlhLV+prYiXKgcwRrU6rX2s4jkId8sq+
jD8FsZ6TKq1MZbYai/8/2XyDKBzEenREu1eZ3DpZLKJfzxkQQnBruFRBpr3MiYYd
SZodr2hpai7d78VG/V66nmZ/HCzO7eys/wAzO3slm9y1UE19WAqQlfjcd5eyGhwl
gFJJSIJJP/UNuAQ+QhplZUEmU/W7bEIGzHFs7Vwlme+W+b318LrpLptTfqKmYbhU
NybxY+DlPIqKLoKaDmOYZ4As1IPzZ0O35RkyVz3bvSTYY50+JodgfmWhjaJ8B/5W
OzTDM2+KG4n2zVIezT1ZLS3lTlFiV+b4FGiNkSdjOMjcJGJSQD2ipkB4AMyu0HBR
4XczOYo7zict/6NZw5/8/QtUQmOUzP1kPwiP5Dl7bts0jNumGA1V24vVUgXgUDzL
MEM9togp4bncOVvQ0bVxWsWWo6Bvqi0WXFLCe8BVr1SFSmfDj4GVsm3dmkVyU6eH
iWJCmZ1oCtmf7WsCecTHGcPSmAy3dqFYFKyUGtIvuyiOq3jYbNwxVsvSzsmOX5wD
t9JAZy7flBoNtRwduRxtzRY1a9pbB2GFcgg28BpsGBLE6sumlIir2xJu3P8TS+Ru
5crv+7hVriaZtjVtVQZVH4lUILUPSob9uSSfSWGYuj0Bc3deb7fPHY92rA99IG10
Kf+hlfADwRkNWfdGwgU/JUI7dECHwHHWzx1fkgiRFjRwxAy5tAY0WjMgd794Hn5O
dMTxV9m4/3ooG3SKxq4Z7qVXyYl06cVDLguuSncVGhCRc3aJyu868RXmglL8qiwu
A/pf+5Jj8QtOmJMydJiLQbYcwuY/DNTzvhbeoMW+c3qNn5NfQK8sxtMnizQgf3Vo
k/3/0CtsKVIdY3sv8tTXy1QdAxl0NeEytdEGOORILyKnqEbXEgFSEw4ktAfvOHtB
nZmVcaN/YVIz6LCaRE627URQeBiwQ8W8ZqJFYUUPrTIKRPwOQ1dwcRkhg8vdUh4B
jkkJ3r96AChTjlEq2yVQIqfWbK/hDKeNOBO90n5etTc1VNxHSvYY/4kE+X+8JZsW
bO/ATkjuxjb4zzQRtOsKfWPgtU9vT46qOG2PFoJQOeTBN1spIZfSsu2xuW7AHGqB
rqN98FMFmUrZxK2R+n5kFQ5DWIW7DZQyfrAmuwbLNjtoIgdODY1DPCtm8FKP5AKT
JOUXpaKjj1imW0+UOGpGZnhWrquUFAIl7WdfVrdt1hv0NXE8RheWILHX8wrG0MCS
0Z+2nguDIYCi21U1yqS8I68aFSofS88nP10CQmlBwIpLcjzI2j1Wrp6xllrgDzWy
w0ySGcpNrTUW4eCThra8vcx5OdANOD5ZaaOtxlwa1HFjtfWoXLHDxa09XqDp1DP8
TSbxPsDvAloA8A/2iZaooW4GkFN7pRY5wkMQoGWaI2xtbcX5hgcZkcw1xz+owF89
dZSjJAxBUL6Orkv40Glj1Y19gOWOkNFw+M5h+kJ869gCL6ZYFUo2FVQO69qOtgrx
gJReZSUB8M9nfacxOGOxODtC1f/utdCBAXPj4He9cdPmorhOMhui3IVl3GqKR7S8
bhlsg/W+VOTJqGBboGCEN99YgpYmK5HbtTWkCi4pMCvX8gzvMgilx+8GMBA19ERn
ZGtszotnzu/36h0yc9Xot2fDRgvg3ZE/KenaYKuKKK4iuoK9YoBsqj5BO3Xp7TBl
1AvLWBaQzrkgGzLynHA4m1LbO8/DS1QI9jFBbOTjRUvYGwFDw7ps1sRCzmMoU6R6
qJ86Dy654mCqQbmJFtWnoEk12xRVz/5B53iULQuPUJIBLfODVEmLb7A9AFFHag5C
+BHBl956G02zDHbxl/qATyTiRT5luIXgFlzjGVQjmODu8Anio8n7f8tQoeCO2dvR
X/8n8xzQTxRR/ox9CqwQ/hi2WhJrkl6DFk1jDbgmD4pB+29VLdUnCHaDNXV5hcde
md1RnW5Lr41LEr/JM042hkhaMH7Rgeent8JTNE866I/fuj+B6vf6RTaWLZ9jNdif
N2bMAxg9za6o3C4rcpO5MgaFfERwYXcyTC5WiEws1PcIH9s1Htcax2QmYCJP4b2n
5HXkOYiOMCZTFCOcYjEXqbCxZ16JeIC3Frp9u8pIM29Q1LIMmn3gnvh1mj5nZ7aC
jkdfJVyiVVMZf3Q/na45mORohLUy445Dh3cSF+8PHcrcc4CwiaoCh94Sj7llpYww
gL63uUJuprj1ltUC/hVKAVR3nELFZeWbvJ7JWyz171yum6c4jTpWszV7wpKLOjth
wMmPCJNpxOzTqy26b4IQ6foZWs1Wrh2aYcJ7YRMmpgnOqjbRoqP343x/U7fQjbMF
1McmlFzPBVyPH1J60UHbj2kae3sl0khddK+zqKmSKEpneDcOSY9A4wi4iO5X35o5
YSULSPTcFplBPJKERPbV0AqVN2Z+1Z8jgvbIrjZeXswVfx6gvgjhfp5rLxPW7Ia/
KZpsG0O9KoO2hb53Jr5Dd1V6YbthHep6t/03rjy7US6WuZ/b4ounyzc9IvLd3le1
4o20YbyvbshFLMzJVrVrjM56AOgOSf11zsAtnwB6Q8wTzUtYxsGkaU0yMYuAPJ3J
qKD6a3bQ5yNVCqdRj9R5hQ1olITQ4hyTeBNVyU/KUtdf3DK/3W5M3YXDSCWEV9pE
Thhni/wR85wmO654YP9JE64T6u1q56usAKKgKI1ZeKuK21o8AwYknzPnrOlRXzjq
DHfkwBnwhdf/5iVRBe7Bqs74irAk0zpOkPoiuIEwSkEvwgbg4aP/Mfd57aZl8mPw
GCp7+sevTijgUWZy8ISYzfETs4Y2/jt6HQYN0xxUPcODAyG0JmtetWgLKRx85NUt
bYuVMfLGUkP4d05zo+tBm1cn95k06j6Tz8QF+To1XTOkrlAa8kJ8X1TmcGhI8/k0
ltQc+eKFK5IKOWUwdrNKgA30Lc2OIhtWYXKFHPH7bOz7yebRv+AU6tjqMLzr8epJ
/jKpIVw31BNPSoNnzRCpGYL7NKGJW7R3JqxNrYyV/sPBSiK7YMHGiX3Wuai8g4Bf
NhqCA81WXELNN4EM34emD5TWPOyOTbrWFjHLJ67YULRdgxBdO8l8IYuVTgRFJsHd
vvcrxUyPCCWX2G8TUSW+DKnB71rngyZ5Fy8h8u3YeAUQft0x92mrt78IaEn4fgUA
wlOAzl4bfIEU52f1GZBwTKkww/Era6dDpPjDwZE9DwGsMQ/5yRoGd/DGkWl70U/D
WEVXjfY2UYPFSS6gvPIkDZMeBCEI8/pXVu4IAKW+e3xWhzmBrE0BisyuLSZ8StvY
31GBSRCdvbVBzbKWOuToOvSATH5zsfu3NhtxKOpfaRtop92v0lUBce4VyNogqM4M
AJwIloINcl6CZqQx+XecNe/rTeJHsmW6MbKZMQQCNSOsealT+TwWqFMbFp6jaRc5
xxgC+Mz2gGPafgxzsUZKdgeHBSNLFDun0kLx7/Shh5iaT1HLjuaIH8L0+uhq+Agn
4ginOIyLDOn1rOqSgKbZ8+drII4WxMp/OW/q8uc+bu+tagQUIDRd56Imp/Q4cBjs
mkNFrqYD/MM3yjx3jCS/KSK/Fyz518+9xxknzpTb30TDH/AnRb+78IoaZPC7RArd
3txXplMw4DguehzfrsdzDLihKGzozHHFjzuqBGCSMP8YyEPwKxWTw1JdqjOA9cE/
9sihAM3QBvYT7WuKY9FV3Pz0scZwPFTYekZuzo0V6fp/4ld7t44dweB3QJ1812bD
0/I+5VxewE8rifUg6YFU51WOB/guEkngwX5DmaE4R9I+kGOKkZ2CJ7TVIT/TKzBf
FX/NG/DVS6W85CmUCFv9ADcf6mQAsvZ+GmirflU0TTGyGYk1WWq3x64R0dx+4Yne
ghCxb8f5c/Ep2uvke4Qreq22bfz4lekwreSWmdUefzT5glMMCG6qah8uFQPzop04
eP2F7nLN90SAavLemipVYa4catggPvP7oHXBLe/m7fxzWFgApVac7wB2XjzJE/5a
kuqHwKLVR4QRPWCAGM8YK7PTxsZNCF9hHTnMda7GyxFTwUeaisiIxC5n8wv3qA8m
cbAWwgqv/N/JN+WR2H85l1ZaMevH6PdAhsAOlTWvcvFCFeWWM/st4W6A6VHiCzaG
zV7Nv2/bVM20fc32fk/yItL6tvQXRrWJlqkrcACQ+P2omHr6gIyqBWwL43IN/8jd
RXbjHsZPDYSuyKHpEoiDIcfZ9ngf8t0FUopYpBHcld6F2IayI6heP5RFTeR+nDtT
N5xpO2HWEiZYAPzPD78bNzw0/YY/WKS8B9+C2+3vWdbBIEzC9ubFzLpnmhO7RitK
Ob1udIVW0VYxk7oJ0AfqXnPCY42x2Kga8sk8Cuf36RyRqVkeQaAEpu+ILg0yhcss
oF/aM4mqOIVdjd6IWkVk9JQIVkdIqmniwgUV9CWJDLK15dZWcr0lsxL96zBpf60W
NqhXLYrjIOrBUR47e2jdq9czyM7tO+3ePSHQ0MHv16RjzstEsI5SY5RYR+fCqT4p
H+t7Kb3L2+64MDrI9uoWHaPJzAH6S2vSJNt+UhXCniDcjUPsDgnrCEJYsZfx60Dk
38HKY3stL1FEg/yucpaRynKfTcIq/eZjc3R9E2qycVVAg/hYlaUCrqvKWRHCiBbl
tw5ULUPds52q6ALQVEkCQcIzsE+i6/9dRaFonVm6zkJvrrJpTgoiiua5ozoKQXP0
mQBasTlQAE0Ysn1UgG4Or/qWVlA/dQ44UWIBRjT8tSt+iOEgwovUKBqmhViXLhqE
u15xqALUA5bcrIlicFklhQkMofth7WvkYObjVN67gPgyhW6QzM6F1Tf3/uUKYUHw
hdM3zEgUXaoEyj2ihsvG6DdBXqFS2sM+kb2BYvNroPwIj4t/BIF5qgsFat4d9psU
yCjWPjdwpFJR28/BKt9Ch66TZRd5OKIx+NbGCL4eVkVm/GTGZwp24UX+JxHCbHYh
eEZzPB8ebTYcmj8HZKjlPLGTo8kL2Wp8yI0IKr0M9Z881fz6CS7etoqs+qL2BxMm
U8+a7HTgrZTkJFGvPnEMwQZz1aQxysN6XxRyJQB/4vZomYkhER+nibqfhUO+Zcng
CyDDr/6LvPliTPXBEQZq59TUiIDUaqhfazSKBFjUnDSovQeqqZ9ydaSRinMHdqro
tvjxeJjHTLD0uMTudV8vYDeF50jZuKAxtraSobkhvU4cWgzqYepdyQe/eAjrip+N
qtoSY1/WoVjIrYxKkyBK1PX9uWF2yF432tDGK7iwVt1QI/V1eIz1sBmnWLAacOYI
yvKMTnqJCNWkz2UpYFu2Jt66X9WGY/xUKHN44/amFBGtH2QT2WVVd6zaTbagos30
xTuwbY27obcxFDU6PWI2bks87TaPchh+VS4uMelTytEHDiEGiJ5JjRFDuu2/pfvm
Bsh32HEmjYEjvlAK7J1A3WGgdpdkGtScHRIhUHGF1LzSuaj0q9p6gTk5Qvf/UHms
ybs4aoH4TxL3M6yfxShByB1nrQSwTvjUq4t+wwCQVrfCNOQoLDbSLgQuDzSKuZdi
OgM5PMNiYyNWuwsFS3nnRWtG00zvAYKOY31Rd793UTgnLzjIG1KNFZoY/vu9Es1e
xDUWDFIHmyMwB09agF5vlDLiUQog6I3pl6sO3hIA21SWnyRhnNlQST89NOsYloiD
w8uBpoFeTMECoXpXO6DDIcLlVDb0PCCph+wYYkaNkg9LJlGK/lt5ngTLDExX3vXd
fDXOMpvyIHFgCy7B8D760nKLxiSKUqrUo2BZLzpuCyJzlw/BlbAHQPLgJh+mzH3E
N2pqj4lrW60qKU+QsElNK2qVF1YyV0p7bRXolS8LggMSM4zZMQiQ2glv6tNpce9T
6502iyldr+UQtbt0fJ4bZewWFv9DWm8zAnu4PFy0UgObDT1EWZ5a9ULgckbGrugt
Ie87ZPl9E+wPgWvM7QQb0tABpRmapvDfWcXwj8efMpwW7KApsXNlG8NWxiE4Qv6i
bMUpMmzvQ+4UQVRkKz3W3e703nI1z42xZ9QWS56r/DK0lSnPwhq6yAyLpoHSHUVN
7OHwNe2pazJnh6xLF6JR6x2QXuIBg5yPnqQCb2+clGm0xlP6ZrpAurDotND39PmF
F9dk1O8cOBTeSgULPtRrQ8uR+4+vAlbDLikSEazrtyLfBmTPnOU82UGl5hJS8EB4
tPM/lJwyUI2+4MBBbTU4DkOw0S9tFnqvJIzNhKOIlx46VjfUlFPZ2wn5Nb5d+31S
v1EQpxz3BVo9xt78v7X5PpEKsgfo8XxlCwnnwLRVp7aN8rTM9+NjxA/sHqgijAMW
7ppHzicgjwTi78p9CwvSfh/oIe0BmcHn+XMaE5eXk5u9hxWzYQa03R1MadFSeWnf
6zNcrTylHjiO7buBVSgLl4lz/oKrGYVn2+EV0/bLrIn6nW3AoQv+wBfajfZAKXc9
q7h/r5x39qZR9lhYMrnaZI9ulirF4ZOhOimIPRqllOOGqK5sPZOX52BNGkwDzyvq
cO8ttA2SB5foSqBXaAuZbUvdqXWJ45hxhsWYU8FPFcu/n4Lc5JSJ0cYSmzcIjJ8H
h8ZXQN7iQFZteC1i5U+0Hhrk6wpx9cdKACCfT+5YqQdzvWYtxTReN8KJLQNP+V/L
GiIFqCElOuX14zxKjDVCnw+rvyxQFqAdU2VZ7vI+itbXzooNZpibUSiA/O/dBixC
eOyjww/uDmT0BC6/IEP1qj66BJXN97y9PaQwUpPET8Zuti1xtrYVgagwV4P7sPPI
azwzZR389KhR7Fok1Ky28/+1Jv+QrDe9FV/86DrVdNVYlOK2Vzn4ItTn3Rbmz7kL
nZIkYqCu1CuKbTIIna57DD31lcW8bH6sqnJzRaejBoTfFIo6uvEwWmUT01bwzQSc
Qk1yH/FYUhlVQKyz+uJ8WCMWUJ2e1mAebeElNCoO0IDZOBySkmEIjLpABFejuWs7
T7jNCrhEJ2cE63CNC5uemb+9OQrqECNBwIzrlO3bTRQx5G2wglItkBxSTwu83usK
ZOhTEjqkTzfvIQsifLm9NTfJ0+d6YbV2djxvHV246RB+dm3wC+J9IiTipOy80yIS
PMRR97uqMNP4SzWm0APNIYQuVav2JapihzPPowbvZ7lp5Ab9qKSI/WwHgVmVgZcN
9rAfsbQlXwU3GI6QY2ZQG82XkJOEGX3FWd77ME42YNEOVt85bDBaSMrJ1lyAmXDL
Pf0urzunoeh8OVEUmGnXDTkydxkVNjIywmr7KY5esGhoBLz4jL9zAGC12FaCjcvJ
4h4yRiv2Y5ImgQjZK8/hzhhSci7dks0pw2dwzS6T5CZ1lLfk931sa38qS7esR76S
H7a//WQFvE8qZRot7gd4K1fyhAPQ2CiGvZNLzVo2lXl0paDu7Jd/kSld6bgF01rk
k1mhMZ0pMaPV0SBV80oaLhL00xujqnhYEDqU77/AyLctkDzavRXCDtzlON6Okj7U
SyCaGGHwcTsgpAjg335aN73B8jAgL1Gf6dQ15FB5RyAT+gy1uM0QIHJH6Kk3PYMZ
EDcqKg+g2I4LZb+kzETy660BIZwpFFISuzn4SYdhYbevUC4gI6gQfLfQLXHPrmbS
UHNLNFh+BtsnP66hzzuLzzA8blxTFHsWJAApJTjVelMKrxg3eDzt6sgxINIp7Qoq
jTjqdlg3WSfTL560loduP5+xGh9yPd1BFJ6MVd/rA24Qwkem7mSxPGelk59UVve6
j33cgJ+Ev7ktF9Tr3ZOSFPNEUrPgFZlGcZPPlOVztyY85AFNuJItPaBx25zqNSkQ
+6GdYXdkJz37JmmIB+jEo0TvSh75vpBshZ6yv6U3NouX7P/ldFgP+0KMSIwlp925
NpcmTWOhRqNlWlAgGlYoB8Xe+pxcq9ULuWsbhDSZGLqvkUk0ex3EZdycDVm8dWN4
2hWQCpqTgqw38b2Y/hXCOOiPIP6gjA95xX579db/z9vjB9s/13K45/5K1hfM2DRs
qC4207IonY2gc6bMo/zBZ/bnSmwWYZtCo6+gTMGsVRZfBbAn4FFW0reQUTksWM3n
hQpsxJqloGIPOCCbDd8o/9Agrmm8iFNIBfLR1lJ6wivcCp8w62MGNwjGpiWcfrYZ
YKEVbH7YhuBV7aQEBLp6VeLOI3BngfUJSL0Y35ZMLccT0KMYzwNvRBynM62e/D2d
VDiKGokVtdKZzYfVCVwn+VIDrK3dMinWPu6O2//EMv+58MCZu/UweT+xNaUkuU4w
cZrBnXI+8hbeZzjj7ygeQPAvH8j/XTsxBSCHxLn54XhqQ0vBJM57KWwNZIyXMu3L
XPBtG62O1ZHG3qH95IADcM9LbhzHin05ruCTZp8TNwEiIrIBBwvczyVNCUp1TQoH
g5j7okIKU46kBety8ffk4G2EDFuFtC0I4vsW2OaAFx5H0wJ3IKRhr7qkKckBhdtW
GCdXPd0/RNqIuxr4Emj/3fMfH8f0IIjsEiVAixzQ6hRLl8v965/pA1yDnLt+vThR
mUgfeUNoZJza9qGz5iXUBW6n4MzJ9kXzYQpr9GRGqzvbQbM8p+n+VZCrHB80rt79
9EYLDguOQTO1haOkyW66FvM4QURRZclJ+EZmSTH8GmFcS3sHHfeiwxKZpUeYznqZ
cJRgbrhEEOLcz8oIOrr71eXn4WLEqt3EClcpleA4YkxeWndEKF+sjb+ZQm40UbnQ
AlTQQKGe3fuziSVyC+k6RwBYhhTFzmW43AA0t3KJHOZaAn6uBaXA4oCvSC7W2gpK
fb7RMdrP/win2iZ19XXx0ufodU2OEeRfoSzq4QhEPu+PU2S3k/oZPQX2nljN8YJE
7jqz81Yl42WHcoT6lCMRWLkYfmq447Xo4uIwA9imKg7vBv4OfTHqRd7vjaQi0YKS
qb4ktzhmUnhShVZ/VDG0XVFsX5uuMvnK2IlrcpJULCtqmFIiWDRikbASaigibyW+
tKUeK5cvKqpK4h0pGChz/m0+VPK9ijSR546PEst4d6Fc3TEOrjjSqYALJCjox7Vf
+rS9wOHDyGyhCZM3vyyJ1BNI/FTkjNYjyQjh9WHrOviXwrWUVcnZwmhVxo/LaQel
9c4gV3K55QLY7TJzYWRVLY1lTLq6e2rpy52YI/J2NA8te4xH1OcSKwVB3flPMKT4
v2FUuGwzMhYha37yn7R+F8tWofY0Db2yGMENka7IP3h9s+TJe7Tn+IpaAG4nytv7
8qMJfIIKHbY9oxKCPTUAcTWR4xX0WnKk3USEvdZWK1R6AA5IydIh/oMkRS5RnuR3
ETBKEe2nGpmGupimRKCjVwdxbyIeKzOrw6qWSXEwWVgpb79z4p1wgfG9z0pNWjCz
EaVEWu54sHiEbf1+SCU9iBSTymVn41N9+PGGWD6OFZp3xa9RJ61e9XmtLRs1mTVR
dPdK0rt89nSKQOrXiaRy8eWDGMgYTHtfOAEn4ZJKiv6ZZzL2hOeImeRcMYzgBZAt
5RSgoyDW6AnSL/POvbSEANGPB0/YjTZVSXBfJECGxLF5DVWb58EoeTID7YVMU8/D
u76aW+RuOjxpmxkW+Nz9/MGWbTZa5Ia5VHuBU9akVr4+Ppnrhw3dqBc1AkNTmzRb
ONRyuS5HutGfJLRrqEnxap/LLamkKGoy0p6zQRkSE7RPNtnobO12N32uUW4Z8bsg
BSVQxVcviWx8D1sXuBv3btX/Ppad19+DDbzHv8Gn8cO4oQfbPlf3Dvl30904c8TW
ug3ffrROfc1BuTtNSlWaPN/4t1Tyz06QEf/gpGvZsbYkvIN/x7z71XqSPuSIOLAZ
udlnIsPVDGJhMkb8P8UgxekHZSlqp1mvA/K3NoAsrGqnv5ClVJGAEQjKXEN+xncW
6rMB6gC4wAKlUvn8bq17q5cG+0RlhCeXE0dCaLuNZ96et6E+Ys9+WkdcjnYThELj
GKLhObftLD5WWIBu+Ad6SPkwcasz+kkF97mGlgi7nRNk2bj9qv9a7gwmUw2HMCxL
Nqp6qejHNOEF/QCLqAkZHCbCXq8vJ+bIOOHVg2kr1/9d5lDRhsapLeZNRmwlOT3L
1hPJL04/wIf4ibp/OGDmBYaJgNDjom3bbN562OMj4tQbnbeWcDi0Wb2hfKjyQGXV
TGciMWMo+AvWEqDV2+0t4OgKf5mUYe7eQQN00x6wrxI/G2L6KTh89g6TgxKfWx7L
dXjX/5UVG/Mdi5kVLzI04Lg2ZxAyJQLQ54R+ByFqW/cPrNUYAeEzEvnlCIYJAQs6
ZRFMox7CgBGgQVSWpO5mAvcnZOUjhgvWDpso1d5T9PHcz6qVDEbnIjt7GBdv219Y
YiW+D7vzGWhTw2A7np5vsghQabHhGD1Cjld4oSQWTIfdPYZbpM4qfXr4GXUz0p0B
ApjHIX9QvT6MYFSG9WFpNWKDZ8GTKUMrhYVoV11aQC25e2zAFBWLVrnfKg9v/K7x
d752UZW52sBe1K83BqSIuT4ov+aLNtLwL4PJ8ipfh5Ofcf5BolMCYaGPpP4ibOZ8
yFGaE1Emam1IYFF19MsSsMcphI9VToNxLdxVHu6R1eCoAfKJllssVJLrKHMFpymy
McsfHFOftah4o3Mkcu8FYls9ouMjqA+Vjlwr+Nv+ek+R+9sbUsmveVEHPxr3SzCe
XZj/ZgXrNMfemIoLwjqbyuDvrXSxPCIaT9F0+axDWcyv+9a0KQUL/OeSAT2xTu5M
pGFs8WvFA+SYWludKpJtUrvnUkOl7kPEKZv1V2uTKOion+rQ1w7Jp/bjYx3Jdgm5
Rwig+8B/yZpVRCz0WStm1kSkpySSmeLLL/P7DZObGQtudoL5dvDL55VQgheVZKpz
p7UOV9a0VyvhksCTDqTAfuJs/OanUpubUS43tFG26FJnmclFq22UxeOmVTNKp4ux
GZ7DFtRWAx1sSiFmwP6epg2o8k4fI5GSE8wbV0FH2YU8azQLiBOyTUD6ziet8eZN
/CczVnJvzZhsiMYCYvqqZvPlObXM0Su+yIKCVpNoGMMdvxnhKcVIRMp4rlligZLr
ch0UJdEke0tpqmaMHmyR8sRNmtkVtCK1TG7R5U6U3+kzJHB0GSDmlU3J758URZOg
CCy0HvKHlFX4/whyg9YW+UKLvs/5Z4UvkaDQPApyGBD1H7IeeVTELhcK5KJ3W8g7
fBwgYFT80YQQiVF7pbh+doeyxEt2zRB4qBxhfkwAWrMeFynHgHAz68oEyVd6VAkY
61wl12cVBBRadTl+ImQWamqs7r3WaRawlJgH293XLTsPOCOtOyjbv5JFg+lDSH+D
ph6TWQtbIEoiHPJwmfuptIPXYZbHHM096pwf2GmOPxmGklgYB0CG49+MTOoRTlW9
2wNolPgJikMIjuKj84KTWFUx6wnYEcRhxqkw+xhpFVthI/K4Z3T1oiMeRTTDlZeY
1kxUihbI8TVBCIl6obEDT7htoMw8jKgWnEFWtcr4z0zbSMHhh8W0ONDsafX4GUzH
HOuLOyZPZNIe9Sg4RyaUJGNDemRpzaQmMsCksmOgZErWbvnZwEB5GMsJBe6f3y/l
5shLjAzASejOSDaNsYsnoFEegfvZwkARoCa/ToAAko7LS/ORWUVo0jXlqczkuTjY
YZbkdzoIP4i3WoIGN2Kb271mN0EoQ16GiOz6w22l4g60xTzy7EdtKTxJzb5H1RX7
63phWBjjLav1IrE6y0ZyfyBXN5OvgsLLqYL9sBIofsO516oYXhQnDRt4W7Mtfpr1
8oXc2PmrepIhTJ7ba+BrAUdPuTDAAppsOOaQkgLFT83Nn4Irrfvr3BSfM6+K+9Oj
N6SvCAXfIVGXKW53G06RSUN3Qy7CsusY8NXPJW+R72Wv65hkgcDnpdvp383sDVm7
OAQrQPo3ex0LM8Ux4FwTGVEau5CDCIK4vxYN3K3nzaREG1a+mr8wYxtsLUvgPQjK
4x1A3mf+E6BRcoqu9S3y52gWD8WoofqEGqX8xjiPtJ16XaeWXACIHi+Y96yo4DJJ
3sz1gQlKpUq+MT5MJDht4UFUeM1nQ274Rc73Ud3IyIj5siindqp6zcqbt2yDtAjO
jdYQ8leto5Y4XhSaIScYoDBjX11K5woUxtiLYRv3oLqOWe+M7uPjI1JbFExEjHnH
YdVALvNhzhN+cC+ssDFtcMhrL8PG/yIqm2uuSvj9A3Rqp4PBwqPe2YgtDNDVswWu
hGJG4bhKUAvMaUJOXPLJlSCafBLA2xSrSlsdhgjvhb5P1O2tLQX9T1MWBzRExUw/
w9VfiJqRz8cBAfOF4+CliPR59rZWiMMrtIhMs7Bq8p7w7NSzExXsdttC44jKCkvp
P849fDYJnzBaGchQFTiQ6cK5hA4eWvoGANi8W37i1dfIlQC7n0X2kwAsR/Qy6iDJ
KSFqQYSACTjPyPdNjbTwHiu9v6f2ClA1A3jkd+SQMIk8gg7ZCD98t95vcALNEbxE
n5TKXz/XohT3AL7l2XIgka0yOku+0Msimi07k2rTs/N1ipSe78WBgPmapIAm2oFT
1yxYp55mfztnO/r51IJbTP9UcP/cq/JZxVU1KiTAnbBv4Eos4ORD3NZdybFJhgZT
bVFrahnuf0LtRNX4tSZRJ7pEEXelU1quDeHJpJOtsBROio4X3lF3AsvZQsvYa1+w
55bZBmjuGEuw2QOD8poAKkaX0wWrFAYBHz07za4qtqC/YD/Y3objVZL0G9HEwSyR
f09Fmvo4u6+tprv+uR4lLjb5ZrqmKZ6jhbpuIyCvhvQTqDpH8RbVjT+WZipjkcjA
1aHy3vC4k/8BdJLkCmKNPmZmHrv4O2X3wFogyBwL9tDi5WMGjCmovM6qGgVudf4V
iijhQEkkmkRWYEfNy1H6gaqcy/xcQcCpAU8PhaDJmlVNR9/rwcMyspT/SE/EXiYr
pvZ5K3JDoaf1CpgCi03KH+CuLxJ6Om7KFJyZxnbSCc8CuZn82TQ1ugJgPQXgRGfr
pdQgJkQSgRmocXabIfcW+RXUjd0E6Rh/eTxPvaGIAGxI7q8o05QtpEtkTujJuvg1
6Z0KCcoTGJwSmu9wmZE7OVtYSig4wXq8rjEGvSOOsEJ2EAhZtITrBfkezuvsOpjt
glPK+EjsLlSYtTxrYQWblXQ7qZW6z9uE65kCj32Zxonyih9QT0GnkDmhFX6dS2YP
Q+c5oeglbhn8D0Jw1b0pE8an4ZIxMN222/TfFje0+sNWbH6cpSemIfsPw6S0s9AO
ai2FPq9R2XaO5i3AFIwEA3LrLRYDIIjzCYWeNMKkPOXNM/aJ0YVgkqWmnHFJ8TNy
x5w5l8h0G9EHDm0gfc6J3427rzAJ0yGuhEQDqNC6nte3O5xSZYx8gLmpwgKX+70+
HM/XbZ9l4cQHkK5oymbIP5/UFiZG5ieDXMtAEh3RaN33c9M1rGKzc9v/VFfRiKoE
6TE21CqlKz/uwWzIqjt0FuS/y2WL7wcWMrFFF2bCvLWfTb700GjDXc5WSvFHvZBS
UBPElT/xPQIVRSN36LGcYLmQgZFHXPX0CgLQD/ng2z5UJ2Uj+rpEOE/K4ewL3Y6K
LiYAhIhoaEwAnGqCJYD8pwj4tG1loqAgtrS6N65PBpYZY6s2im1ettqvlC39+VY3
pO1Hm0NFImb97YjRKIcyDi107RGE59Eub9RX4uZ3Hescwmj8gpd1dqZvjJm7mDAP
J5EMtcoCrVaJORpNzgEQKTZ5y248ybELrVOl6JY5XXBdXJ4SnSNYNxwRHRvXLJ2u
vs4pCKpyxU9CU5VOrsohcZn3DkzzlouSNRfIvS4yPSRgn5Vby2xZhiWEkC5YiRA+
iBTfu7UObDMAor9iiNX6F6E6U67DaJw27drEmkzYcsjRFexRwSVYCNQvEFCfCs5c
hqNXEmsh2BbmDeM1k3NWpCEaPPDCV7e8jzSMUeZ56PheYeL92StVZlzeoJBvpi77
NWT8QQINS+wgqjabWofRgbfjInd5m0/w8f8uvszvT+ye0c9vXLhlwdMDR69L0zIZ
cVyAM2q51wF+2SskOR4RN/14q8zHZrrOk6hOXcBQ4X+kq4kGqiN3Yhkl9ycsuofD
Kds4B5eFRTt5GtxF/88sAMqB+ecTu74xdFGGwz7tKabNsr6HVg5pvsok5lDWmrUF
l6hPLFC652yMvENXzswJhq08OurHgalaMwYNLD/96jXjRIMrw+iQPDDaA0uE/AJC
kA02porzlp6xl+L56YXOMlAoKIg/llVx8Rt3xblLwHTcTTK52v3tYoU3AGUxX0aX
iB9Pjl835IfbEJKoa51AQ2NMzLKx+EHDJR4tOZ6EKhetSjq1dorLj92pbNUGiuG6
z59g+9xULF4C10okGE803X7I2sMIp2f8tkbvnwAKfa7NOJq6Z9ceUF2Q4u9i8Cb+
3QcQK0En9PT8tEhqLtBY63Q5QRiTsZ5lJmedpMVphyvzLGqPbiLTVISqCnoD+8Mo
ACV9pWG4My294/LgN1Pz2PfB2DGbHk620k1yZfvACKSLSidIogTThs+fDhfsVrks
5BSsW/SSvjgiBSvxE5EkK803IEGkyOACR4VecVjw6hhHD716e26+qxl68iGMkUVd
5i2mnHmKw2W5lIBeo4gMJdFdVHmotwCIlSZfeEF4MyJ9XkVgnr6+QKt7F1fUrqTt
es7J6KeWvp0mo07vTbugZ0aL6LNfoaSChrYEtiAdSUOIhe8A296rnFdRidLCUtIu
D1C5Ovk3NInlPZU7ZJ94w1ApkbLD6GMXL6jTLZDE+oOFmlmDppOBrfmPhpsTihDP
Jt8XYxl2Px4Tu+OlRDJh/qbcxYqzln7wi/LnM6UdkzmohmfVFrZehoz5UjT1u7WU
B/3mYkQr/vdQWdEW9ufyKW94SEHnuZYYEdKysAPUpqHCOyAOkAN4LW7paXWj+t8k
9enQEzvjzma0dG9szLgeDrW/3bnt8a112Z9Z1X1cR8lWRWjzEtZZBc6dRCQ95RnF
891sZZ3AjORZXyksXdHOjn52ssH7VadDLQPzmaqXrkIt1PL2Dg+DGPUfclTnoecH
Zum0HOn69/sz56khjTsA/aPbCoYnpowqehncZOSf+u1C2JqhxfciSKOuxM5Ru0YG
IDkzlWtSFNptUfU414xmVIdJS/aOeFVAEwWu51GE2YwUPOKvu1pK5MjCUEOvsooC
Wg6d4DcrQz7LfmPEzHq2TGR12H8k0a6WTnJSMovpaRiUoTyF1wQfEG8WtmdrYs+z
KxDnqK7b0o7l/Pl4hqSB0vxnXhSD/6rAF3UJM2lyYdI2SRzwdwlZBGAaAWJi9Nsa
pSQCJg4B1GWhQ+vgT1U2GKK44hM9Z1LOXa1ihWBPGNnnhPMvlvsy1QWl5lSeFcD7
mf/f+zDI+El7UgW8VBkYrIzoAqKjLpR4u4hQeiiqJZ939URKAk6PF3I91GU15ANw
ZzbGualGJQ7/wsQkUrmiZDhsev/PrpF8TmEJe3uW4HatYxiDD0Y3dll+eGhYb6vl
Y7RSA4UN4kOihui/MCnizD6o4cGb9kUFn5zoy2vM9jEkBEVBqEVmASF8vZr4ushs
ejD2PA8NzuKQ14uDqJWVno5l2C9qrSAiTpiwML4fXx0R3yzyavDosvskepXm7ZXr
qOXcjf9RJGXnVXmWH3SGqJMeFXDLHkYCT03MgzWC3ZmTxWPCJXimZJ+bqt/e3RIS
N14oU8QjNaxiXGWXDjhm0tXqTxOuUahl8zycRB5tCbFXXCLIiW+7zoFDb425K3j7
9UCqJRLMYNOXwNNZPU0ixAasFUP5vPWV7IXzTpGog/vCsGDvq8GZRj1aiH35WyA4
ESJyHakhoxK3LSjLNfDZvbvoK/cfhBuT0mGsUfuo7YlsiueNPehQzTqgkQvwlupc
So1A1GpLaTL6DUvLhVohcf0nx3dMy4ibqByn1j6htUrvioq+SUhHW8Z8E0uC6lSH
lG7U9xqA4jT3sZM2p8NY/MCHu2jRhMnB0ash+CrSeFElIw2iUpA3id3LDnq2gPUw
by/MOzkyLDr6/J3iiegF5GFLCK/nDRfNYzMbeQ5wDnzmX/SI0VUormbNECbm0IOR
+96KDmRiYTNNIxzxgweuaypSsaXhsp3fDNTWrfvzj2fYM/VQmA5l5pq4bc5bVerU
Aa+1WcixcWlQCuuNMZwo+AxLKkOV4Op65SjMzD0nJW1ewe6ixpB8royJ+F22Af8C
+tzhvfvlCpC3P9GF2lD7KO7ybSdvaS+mmj3mNDEfJkyFzKhykhLMsNLsxg9kDZtG
hoLJSrXTFrZ506VegB9HR1kxHg0j2tMNpGT/f6BPVx9f0tWS7rdlF+vOaF8zjFyf
jKUaynAkUtixwRALL9HeILvOR8Mgj6NWyKtxVxLiuHwY8YcutR5Zf8+e/YCQMakF
YJvwPcM95ByaZADHs7eWx4TbSzPio7kLZpZ5KIqdUNEG9R3115Si4QnDKNOZ71mB
+unhI2WK8FMWSzflJhTSMZnXN9lxiCorw9D79Sl0y1GpHLPlmzx1WYKVKOMRVSZd
BMXZKH15WPvchST3qGxnOBcPFq1XKhxSPkl+D9q4jhXASUIgeyjYZLG3dHSNrdMC
wCWTva+efy7EoqPk1a/KRtMrMTw9OC8YwS1hmakYp6OIoqrpAlORe7DN1B1ELPlQ
d/ayxaOT8gTJWxZH4+rGfH32UI4ujXj7yyG0GMnk3g+YbEik4e1Iaf4TYln6yhJA
l6t2dR7dxhfNvGfStuA795LHf6V9/8GzwT+SXob4OMcUyubDYPBv+elo/3aNVTPC
K+WSGfau0PvTStmwhSv6jfqpwpQGDh3aDR05epILuv1oc2F9cscx13pc9sni1/yK
jv/FKxx5jbexg0m4sYx5+7DTGF/1hf/EP8dqfiT5xzcuTXA0CclWrPNmWXiF7heI
BLSjsSfPDOrdkACtwjxssQYM7s+GD60RNOchKujM7wtZiuLeRa2obFg7Oy19ZSJl
s6EXMdJLsj0CHMXpgp6ri5RjDMaJUGKdO9WCU6HVXiQE3FFy9V8Ac00loprfgoDW
gf8sZ0e9BvXm9FHph8hf7MZ09rW1kzOrwVBLRh92d0nyiyCm8bXvu3Tu2gvvvodl
VZmgxLvb9juFIXC3NMNirOiAkWeTO21pmGLsds8XU0sjNlxX0Hn6eYrFVOka4+72
tiCY/2UnlJ5DzO+XRe9fONiFhvJTn6T8EPXCvCaErw6OnEGJ5wG+eNR3VehfJMOt
ve4lmEnaqatEMW6exMENrNWfy/u1V0M7owRasFrZyO4IR1cjJd/ANcpug5mbpC98
liFhtxxDh/KwOHydodlLbmH+fWIhvz7r0J7h/jotdVHoX3WCzWtpQGzccSm3EcGD
On7J4XTAELmuerDAG6GFfxW8pzcDfro10T1HsBm7XNsXw3OKiVxjwV3a+KifNkxC
1kosQiVPV2s1bJxwDm4hWeI031TP+Yc9kGtSkGAfHP4GMD4Uy8AJbOpZQUgqJyNo
MR2QQMEhikDJIf3hJ5ZSor6D4c1PUvZ/c4EDmyXb3Tb/yJGTCuB+65FW0hy83u0T
TAkjtmFGQ2xKbZpWbBY7LXLplX4mDxPa+QjShOK3b1ln/Csubwrppl19FDIL4V/o
/eUcyhXNWIWE5tU5WeD+68cptBIfc9b07eTLzHqTJPe6mUa8lfpYSFMCW14TZC2a
gfA05qLDQyH1s7ppwdcDN4AE2morf9jMkAIrPCqDzuEOf++iIN+4TwRODXxxnGcd
F0YfqQ742PiTCOE7ED5aj3+/2X/EuaCeP/awIyVb/d57+PaAmeboBTrpNkupXyAD
pVd8Br4Uxs+z6yKpH5VUhOjwHiS4I3QQ8vdo9mXXxfndpWR+4syhhvAiXGbsS2GY
RgOklvKjP5D4HuQOi1ZdY5AE1PA8tojzYreFlXUQY0eiLyNC7ByL+JbKsjINa2/K
4KdCAsEiI6cMgDtoVTG6dgPDWvteur+sXkB90QlbD4pxamn6yYXW/qPqaBYsKnx9
esls+mj4E+Z0RHTSHdWDSCKaFrxDb4mM7ZuWqhgDdNhM83r48raYPXAE4xWYWTH3
szFdPtheoYcB1MqcaMp+2kDqTSDn/cz/kWFhXlsbc3sWOtfjAw5qesa4+Jx/nMQY
ZiCwhCFp7FS7dDsImbgGL5ql1hwmn7BcUvMQ33qkgboKfdkkiA0yKZUQ+ju7VSK4
xVYpIg8eQIrSlRH4Lp6385a0242Gd9y7dLwGQAdKdsExzZRyqOXqeSe6XHD5IfrI
bGD25viibML3akbDtS9uQxbeGyLTloyEpSSpZC682/wdns7SUAQwR8/55sAD94xm
4rzbaRS/+NVsxZLml6OFIXsnvOROQgtUn9Kvdgc7x3cEtS9e9w6sWDjbXvuWdZhe
tcjN0rCwAs07CyENivzNxlo/B2U5V9tnaYksKLDlGh5NdV/mFU6cxE1ECMVF35/t
Jfx7/icX1l5w+aZeq5tgxdPadqt+SBPDfCYahXt7kfCOXPV0QpaaWxanHqxl5yRW
lwQjTMUbFD7BHhY0M0IkgXcPEYOOlEMteb45daFmmg9bZ/SXoIKdQnx6txKndhCX
WqnlfEvR+woQQ3wvcj+1aDipbdEFMukyYjYIgp7F0EMaWoyKn7hZ8ZmLa8NJ9LtT
OMMSrAb8XK3Fa++GmqKo7PpaLCC9FwK7e4p0cNmr6ltJzhthJcJvTiaiuNdWrsW6
E4JbOTDDrKV/WPtMcwSLH9t6T/ehCZlrZW0o61tvIgn0yq4VUhpHZXVKYqideMQV
sqoq9p5mromUpWqnHLeMcLaerAcgs4jlop7tL2fZ88gGkKrq0GB+MalsO6YVUrZH
096UL07iVDwM1WdXHHzqvPFog5t0A+lB8mMl1B7T0Afr7/aSYVNO/TV/MqJTJfAm
oaNRHYRFTctV4NX5WyfhOXVA0VIGJy6PbNW8iEIyAmuZY4gETYsdTvGt0ghmmU7Y
JydViwVACalTTGPd96msBOG6uU4blnrNuS/wLIRLUbU0gWdhvufqy/CfYdazVqdP
4bOV/yTaRw3PQechOT5fAINvTIy664qTLORsuMChOLDB7hjyLt+F2ETCpF53U5AR
MQEvLkVfeX8x7McqyP+pjW2BRYHJ7Cv3lIvLY1Uzl8QIotTEBHKEaid0RQ0YRd4z
T3jCLhan0F/ZnBnYBNFrRVWysQQVdgC0I0v58SQUUaq2y3P7wKgwBbghgNZXDaqM
iagS8953m/KWvbTw2t4ovCNMLuxxbPbesOvFyJhlk/o6O13ZysCn+cPUMRcPbKLQ
SaRGV+UYGo/9QmOgcLILgQM5W5VsIzijZJMHE2X2WDtKnRXG51gbMquoFf2NnZID
89jCC8udQDTj2WuLWfVXt54ZAuxAkWNwg7279ev8lTuwm+F9fuASqnrkYkwMrBU+
kNTr0t4njEhrQ4LjNO/GLAaCxy8GePiDbqJ4NkvguYpNyBstaEQsMc5B34vhy2Xb
jIk4SisR21SR3q8Gp3g2kxWmb0dTadvddBdRDMBy/DkEq6DcjqG9UQQd9P4/7cFk
o5AzE9YFsriIcMg70xzh84D/Ld18xY/KTy+ebLKRdrmMpzGg9wgjdxv7I/zi0ZFK
UQJepO/1/GUhwHdJ9OYb+MaxtEi/hK6KU4/MRivjEX7vtLMzc6THkChX2BtDsy02
KvHsGkgK6XK8Y+uM57yq9dRMUozRJNnzqQLMmzOTcznGMWGUvbmblt/U0yfgFDIU
wkk/ohgrXqLsvaCeQk68O4zZgBJyntOoPB71iu4aOAOwNreh8VXnWzAQphEKd30o
xhjxS7Y8vEX09vlsdWQZv+qrV4B8nZWaTYRrAMtRuEsG225Z/7bmQItbFjoN4ZHY
UyLbBLRNaZSD8qgsySa58qCvk6rK+TP8BYDqmFknCtRirnF8Cm1L6MMr8m/kZxGQ
e5fwXa1slolDCotTA63Wr6xbKOqNROYAjP9AYGBZLEObi7rgQ4Svkm4pN6NjgpyH
cZPwFxoSO0bcLc81OKFyJ9aTn//gSWpWA4PpPjD8OCWE3vLwxjs+VlGAC4FKmpaM
G/Fp26ROrkNBqSBiFw0QAnDaOF7PzI39nVoQmzpkjVv2KEnywicqkAfeeoxGLC+l
M9dW2YM9/hTmtn12KMKw0T9r+y18mHdn4WFD93W/F1ValdlgKy8KtR7BDRmThqV+
jKJghp89mYuHWTEQu0fhLFfgyIGjQpNuQ12vNdocOFY2yz56LZjfctq2qFrPs5XB
oX65FI+iIJCsVN09jdDz/3EZsTmYQBX3vIenHki9klwcBhRjDQ3n2Ds3KG+002V8
epBRsJL9b2uP0mH6Myoq9dBkeRK0FWH35ktUVmeG2dXFoIdq0tWBeGUv1UZxQ6wE
hFKyFcFwl7WQ0qwIQ+MrDkey5eRiGBJG6znVhBFU04HzlRs1FaHLb2jdHZulMtzH
SuLXiZ0E9QK5KJRnA6ckgUzvGDjSfUezc8QTu1E2lhb6AM9lecJYkc3EJ6aHTM5u
/AtVW3CRX/1ASf54XIaCHwl2ORIImck6i7dUEkQx1MQF234LFxDsnbb0XmAKyYOa
eGRCYBDI0DdMg+FJ9jqTY8IgSJJ+gYlM4WsIQHJ02X47apOuUcru4rSd7vNmUaCS
CD4XgNhDiPHrHUnHKhhbnzjnzijUNCOHDxuzxa26l81NjGm1253HDktiJWRTsRvw
EVTp/SnVMjdoaqwZ8Ah3LS2xjOQAlNNVidcE6UMFOrcxhrL4sitJeBmqq4542NTT
MIFt9T48npVEL6LRRuYBvyYuWB+a/Yd1Mn1cXU1Y3zvzakRvj+EpQ88V6sRoJSQ8
RUJxFEBJ61sXoeyXGgShD7iygKQwIa/inA/iY1FKadc1j0eSXskTPQGm59/BMliJ
zeMtRBPj+CeqHZWAxFaFBYCr83+EH04RXnBF9zKBQQ2amlSeXoo+V85ZIxXOevEd
bQqIIdc+o33iP4TndkBBEzPfJ/WPgbRwG1tSNNXGfqv718EoYzwgalzsHHa7geJy
ghvO/CAoTDM8fYO20hE0lO11G50z85flHvXB6YXphJKsYZiQvyXVQUo9KmwNOPUP
UadE5iPcwkDRoLRKo6al8cax8BmdIXkBITBILE5rG3zwbtKokDHkz1Bjeda5n10F
L+dN9ci4BtKfdO7wuOcDhwFg8kFPsAPlRLCukYiboeqk1bAPlu3LWkzxkSa+CGlb
E1uJyYpT5tztGgwFdRcpsQRj/C8lU8vetX2fZxZGGvy+vmY0uW/GWIFnc86SOaUy
w3Fvf6yAnrC+0IaOZRMTKWu83tXUdTVTii1Xx0gE0E1GgpGA5GRKUpFwJEf9USV4
uvkWieMMRIcjeBGdO2ZuP4yEDTdtM5lAt8k3+34ucNVQmNf0p6mJtXAHMvX85Ot0
MnTHJnDc64NHektjJPrgVSLZ5VkqLNRzmVbJks4mSHaLdBq8ntsh6ub1+WQ2um3Z
toeF9l7N6hxd1Jd5wfTUS4btD79kMGrH0lF+FR9Ym3qhSVC1eFx1xRK+GmlVCMp7
SNhEcJ4d7uihysktqSc9aMbC+i3gt6sriqskLexr3wvf720S8MLcmIkqljtCRTaT
MS9X1KvyCoHbZ0e/BJ1HnfMpIJGqg+RZ2ym/snC5ehowI281upbWGBpLh6funvcq
V3gqvz9fKWEYRD+1RSFUfaQh6blRcxqRYxSR7EmOkBsm+cX49EJVnh0mbg0Kk5vL
8eunden4mSllMFGO5pJ0KSsSLuTww2ZWcEY1JUJZVIJR0stJrvlxc9Dl04redqAK
AWnZoqtvfudCi2HgVGV8kn2fgh59jOcSbVxd5EgM+rsw+13xkIfrMyBD4YHoS+CL
ZeUag5KOYGRq2Wy9s653XJeecj+mFZDcyMzclTHLjXuZ5c5Kjgu8IA0hcncGDPGr
R//S93AdOHI3lRSpxj1RC6IfytNpZmwfbK+BQqJBGT/T5M3pYtg3PGTaGogBYYiQ
55ziF81rv6L6qbP6nKrmrXFOtdN9HZhFZ007ipaXem/yGAvgb46cKItnjxn1xGHw
aeQR73TVk5OIRNEMgy86JexTQC96FPYwP8oiRyV4Mtkdi8aXeVAc/RftFCMWGnz8
2ICgEruNFnzugTlXcnwsJ6cm1BQWAE+1kf7vfbRLbg0x4O2Hm1/YOd+l8fq9EvGQ
jWZY5kKfN2CmoDIEHT92F3HRAZgB41ld4sfR8BOniwSSaJPizx+m8xFGYW4kAjkn
TW4nGwVTi69rq3WFm6t6Op+8J4emTP6rQ9W/eRSTCMGHxt4z+vg+GSv2NIMLLD1r
wvQFPrzSknVQ8d0+Qz+pSQhqanFYjNnFHYkJc34wZpEr+Y2g5jfskDE+xARZAuQx
gocPk2uxr73jTblV0GETrH8WgRxTvG25HiqRoPjndIn599yQcWZFtTkrPlbV82YS
Ljz2+xsQwtTW7I4X4z18pqfEZkOVvIr45bC6aEiSbcV2moMjmG3g6s7saeAbR8YX
nHmIjOy7DzpYYjJTxfXFkP5C3YD7VvUgRyWBoammTlw8ymOS8AOX+qduN8okyS3n
+PaiXjoXJAyiZ9hacIQ9aJDGT77E6wR+gXN45yYa5GO9uoFbXmHlCXYFls/+PWV7
cJYi5CpMoVllh6ZQBGTlU4m56PJ33UAZbzTfuDjySTFTvsv/CmBSe5TuMox8F6lV
/AzOJhKLg+9gjrypQTcZmSJkJzHqBhF09EMsLTbx6GzoStnoYyKZddfGiyAE3+aw
rXRZIimmNErjEemod0K+pvUXuEfNLE9/pgO6TWpBI+zuCkJqHidm9x22PIBIknoA
II2hjgjRdpuMFgbi1CcORuu4wg8JrCDKWVVecOvCBYXpqr3DGH0CeIo5FI0QvodG
1Vo37ZtQGz6CNxdGy0NhhgoybHicGaHUMAawP+umxel3p/tqxKzNr1Ke/UCrJx9J
Dnk4U3MeCBJBJ9B7QwyNpwjDr7WGn8eqA5fmS8X1HfOYhRiGGvy1WuBZSeSSe5lP
lrJ9mmRElxvsFp6fNnDsOW1fyG98aQ+sOoS24FUqvxB1ytWzlHAJNdk1uBQrWb1u
1UZxBm+bHj3JJ2AI0sQzJkX1ahKAdBTgztnvg6KWorhJ2VGOf4baZKzlLS+U8ykg
wfbtcNOY/4CDJN+sU+/rLRl96hlK6HUXtdQQxe+MHLBDXDbTdrl7YO8XtIoA6KS2
k6nx/85ndEEe1CCOscB5uy1gcHykQh5hTYuQ4+nuAngf7EpV8EAooh61ntIBXB0y
rtUWZBSCs8caEVAMu4ThCi0u2kLzTqMKx+jTk/kMktRkDe0rYG5S5uOq7wkC71sQ
DX+vw3RZG0QYypRX6dMofmVd0vdvRjPtfQTHdnuAO7MLJj3IMfwapMuDLGEswUd1
Vbr1l/32yRDgpTsNsh1a6EZLHY0NFcdpbbYKZIa96OkONYbH7KDDTZRUebVVCzpK
gUvYT3+SDts5bhHNBKy9vq0g626/rMZQdJ3MHELAhLfYLUbv5ryR96L1lW2gpMdv
R2X0afssBlcE/0I1U8ilPbY21HCwuaRQVbbuxTCS5UMJ8STJ+xJWZ4TD73Lg0nvm
qD0c6lvuarC1iVVx/r9UY7Zq9spRdqRGzmjjmCz2PMgxzCJa2LmZ82KoWWr9rWH5
Tdnr3/7R7okZsAlGdpQK0yIyS1eDYycxvIoR8qLrFm8YPKt2X2EstZdGbv8NleQ4
eslKUAHBZgIAoVRCiTxrsjOjARmiUSiXA5LafVbdXT87hnm61og+TI5UA6AtsLq0
l/JmS73zpB+ugPP30qPlh6wn2a4zFCJ0OayYZKFKSM840cJhTlaPBTpXZkJ0FO6P
Za953lPeDQEdstlDN2VB9W3JBWE7dt47uMEW9GWXRirAFxx4MsNylSZSnbedcFLH
ABBVdFGaUwxaeVuoUH518icRTAkRgFBT4IXo8UB3FisyDU9lssViYgon7+L+pZmf
IQS4W3Os/xrVBROH6VEskpza/8bZxskGca3+PAvRT4n/ireLAq4A1PF4jNmBG6gj
Ai/8xYGFzyTa1fe97bpUvjyRs2Pk8Dayt+4xc7GW9BrVeZWtoOh7SlFy8S3NqKmR
eK4i/7Ptm2dwoU+o4asQC2QPeXG8VViiwbbOwHpMVs4Gwmq4+oqR4bQ2EeYCFq3V
lEKGsnipJgINwELXyWBNwaNo//2cUHgwTkQNQa6SneLpbHOJpyc7+acmSml6VI+z
mi8phqYdGkTgM51x2UqzPaPW67LhK4mxNSrXP5aCKNBhK+njhXMjBfMmqfTsq8H4
VakGhuID64uMZEaEbB0YizozzMg3JUO+Yo7deKXO+gRp989g0p9/lkpEd9P7JGlU
x25dLGv7FttBUYMG5supesY3l41+sZncAMfIwgVlslf3crluDmS/FU01gfha9Ask
JlmywXDuwYBTua/TDO/ZU5G8loBkg5KNtp9tHFYiCBswwGYyrgOdwRAiLlpT/8zK
Y/vBPk5MPSU5qBawMy3KuXU4+l7ZdRjtvxeBkjwd+/ieu4qUDf9a6hCGYogRSY6Y
sX5ig3bAT1ey30M9zuCxs7z0wk2R/b/glQmI+TlEc0S2ok7lZGmnxhORJbFrbFCp
MyCvCRCy8SVJW76jsPXl0IrKPzvHPzQ1lFMPGUKy2AWfqn1lCnE6as0mlPNKP84q
5z4nTKwjz4dtFmkoFmhRVFzV3kfaKF6VqiZZA7EebBq5qAKUCfuUjmoEqAWtnSl6
Fc63uqkA7hBJQ7k+mOaCYrAVACYYl2XPepWT2j0FINwS2k+qc474anwA/oUQuY9T
LSgmH5y1JdZnEk/GVp3Wt26PDHKODPiw6KOTRawjkQwlUdE19P1q13FieTuTyH3b
MYgICoKBWBZl0ko7+2N8XSo64XLvUN0R0qe3x4BHHaudKLi1nHyF6KoRZu22b0nO
DSFRH0SPmYpeKcz3n9Dl9mFWBJ6sPjr+QGADLl4Kw50dHsGdj1Cs0jtr0MtGj22m
17uLdx3Vreqb9J0MXgav0TNaSzEU5XrzQ+KB5+DJf2OC75Rq3VwgJRR7oW4szw2T
znPEbJU61HJRelplGEZP8y97ArDI4Zr/Y+5m4AdjWztNyQ8XtXsFk95MDP1sxUVt
e47gknFlw1w5bpAXaVQU9J7gHwnb2rYKuaQMF82+F7jB/mYNAyYn+Yf24+5ViqEA
/YujcT/ksGq+RNVdNs0RhVu8xwhikHqsTQroUBScCB8peIOHtzAu2XDkjk5VP8qm
Yy6ISdZiYLc3TUhC37uzQB5ADQ9FUzNRm0U9+cW5SqZZ35okAzU058VMWKwcKQyB
GAy3DEhLu6CxgPx0tjLqthSuhKS55iqgcPb2EJGzCD0g7k/tS/um3L69KyLH3YFD
Q0sM8zsQVVOqit4hOkllFGQKlNo5Hyo2P2dGkKIsRap0zwTzvGlGiyVC+Q7/oOkP
UM4s0tdTCoeSlRnCicghYAza2/lzSoq20ccakzHva+ofJw5TXOtnSczVOlnEZis8
N7SoTItZqVwkc6LX85NBrfQ3xsZ9lAInR0DogIcjPwGxXG3ZJmEkdb8nJwNKCrl4
bpRkEGzv/usLKs6A3fWoIFBwNFxzVj+COy2wl47n3GmSohPLYGMS7DRsKyhBg4lP
D2MMwj3ET/37DGeIuSVnydgxL02rleyu/0tn0RRCUEX6aNAbZJQzIUWALCU9wDr3
c52TXpMDm/Nb60DCGkf5WYv2WrQJy+TQw5URFFNkkS9Qr8uQitOy5VcbuwgGjaz9
YiMkmkfLPV4qN2wL1sjTg3hdCOjp36YICSdtod8r3FFMapgSL67aeJGp3MYk2Gb2
ZG62sLiCYOLzjGMr+TMLFs+7jIphaY3Nt4GXOBNSvGJkbXwQ5Wqm0eEp1oMMpXvq
XWQoaCxL0ovvbtQPaHFX/bH6LYl2kV20iLxJBWef5rFc3bFp/UZJsTd1Elcbn3Sw
z9uUjhDEPInO06//8QztOD9bxX7eMRarvmRArnBe3rttOGvXyh/Caf6dbKLiSH81
vGINMYmeLsgFn4lOeUGSu5CpVzPFmcRQiUvys+OSivDGYGjsRJCCNWcdXt9AxfG5
/HCRsjeNsPFQNGrBFEVJF3/hfYG1mRoyn84JY0BU3YvEA0nhdrp39fNgYvbwLwJp
vgwJScCPt6dOTvjlbtqzNXSjJiXXWRzz/Dsrzjb1aVoLedXs75M+I5t9QQZ63EKA
80eoVQ2j12or5/vPPhmqPV9AXdU9HxvxnLMB3cN9PQjOguHvWBTahjqrVHv9ziOY
bqqZB52g3FJGom+jWVMHITxCy3hixOKInIjVMb9NyWhnbvTWNy6+ZxBvVyqgJSjy
GmVZaP24Qf0TT5lKSPj+8f/QD5VHc6i0Lc+eqVpCvUNKyUdnz/m3SIvmikHsm1sH
D6b37YNI4e/v9h2xrCh7zfU8DygZ3yDFk8Hq33VfWFlhuzHhRneuEPoEk1c99nr7
VBn/pjpZrNN6EsL54y1rorAU4DtYt71FAIOOnbIhRG/HVU0xs2uJqUAXht8/jybT
ywsjhuKK/OqGb6AEf8Fn1jniWmhLZ7i2kYpwAmRFHttpNEFbmHOQ/ULOi8UZ5dkf
cOcGnBsrf8l77CRgpyH6Z6yVjZ8QZmCzqBj64JXzdoaP1yot2YkmeeGx5qIIm04Y
Z7xv+DpN4w3JM6wOYk0Yx/AHxgxzH3vuIAbSN2Shn48oBjZijXXHg3vcm8cyiV45
cTsztRKrO7LkdoHwKVCtG+Q8wRr7bjdC/B5GOrhuMI927vhJOM6ZX8SxiiwILdD/
ohjA2CYdZi9WWx8uKbw0l/L0p1X5yOf5fMX4I9AX5sNC8RBkNeLsHdj1IbNwJevw
ZnucruLgDjg61nFV33ei4NUwv5jeD1BtyirpC71hNlSlmIQAUNRcZfSUir4tcKCz
R5qwQ/xKFAtITAYUoibYUv0/d80aa+a6qv+YAoFZhyN7tjHr9AxT1qqwlqrnBJcz
i2YDVVqmCE0MYh4O1xAa+66Rl4Rs0HBAW0WXZlzpt5pyw56Ek8THVIVHRlsFZ934
ckZfKTxsxlcvDNarP49lNB2A1wDTE3x1ps4nr1J9LG0jRvBBOo8E8Xzl9oupYeac
UCU7YUjed2qa53IunfTkH9Sw8CUh7ZPPhQa2fcnw/EFjY26EmhyxT/TGZn/06CMe
NsSsJnC4XZikEhLWgfadu5a9QsT1GsUorlhee8euE8XBhUAw01IRMk1KOPS/obgO
12mbzj/DVcydLB7emGmBcZMHVnSJr0/ePUi9RaAbvTkPl5ZdmvYJZTBkGRtfA0jc
AWit4Ru5fqwiNoZX+2enCGJnDrx22HbHW2DK+PyE4RRlNcxZSQquE7P9s3q7ecOW
0tHz/JgALIwyDjVUj32FGGP4o5c/nI56XDXb+N1Llij7UwkFyl2iMZQ0N5QnW9u2
F+QGDvYgmQmUADVp0dPjwK2g5TK5tPqOnNnCbopeuZbpyOl0gW2UXLk/8Dl+hjL6
aWI1CzJjGXRYOSfVhUDAes1XODOQtYNX4RyN7oTLAi/cZPcPmYTlvf9/dIz8rXDL
ftZvg3m1wjHX2rYBnKZs2FPXTcr2KvYSWiHzQiOVoF3R25ZF7kSP52UEmRcVUaVB
mNy2iSerb9SnvhJ+IzvhQpDztLkXSrx3VUsxkS3CUk24iPSew3dOSbJ9XO/qzCNW
ViBE+O3Y3FJRaRGUKu3eEoUniLQ4hq1oD64fG/B9730uzgfqrMczeaUCVVZpfzRY
BhO6c2LxU8bJYP3Cv6Dx7lYkzP/oPJlcfjll6ncryCIYUuUVNUqrSG0amlpNUM5w
P8WZo8VbySuBUe1A8NE84OOvkBjtU6aHJMuNGDeILnO86g0KAS4Dr7bopN6cSHvZ
pX27Vkm1kb4uOk9dhL4c/avRd1ylLh68RDmT9pRnM/r2yDgbFN9upHELQdSah10S
TuiJUIEPyCvRGGVMKe7O4nUA5CuRt9Ni+YEoayMyD+L4YMYEavYToVsOu4OI/3Hs
kG20+mxWuxkf4/+Mf6ZVS+k+l7QfHQGqzjdRCrLFrW2dLAcQ3bpsRPAFTJ6I5Jag
aE9HdROBkdiMYQh6KzkWT32sGiHoKyWVTHuOamJf+B8PHbamM5yXHXAB8IaSYOmG
KACBbLgUltq0ncMZ8wYdjNO0Yi9LIVlCCwyfB8fMyOQtTHX19t6rfiE8RFeza/8V
FbFj0ASo+Vx0cAOkWOnR0PMGGfAwiCWidzZQ/rGIyAicW27S6a5lkHzC/RJX1bgK
peLFSjqTNsQfiUcTdaKQ87wcWTi/q+JjAdtIGzRR+G9Y222cVyHXtZYFkEG6JtCl
Ilgv6qTbWH8nQTXoJT2kHFKMZMrzFESwQce0OpP+3Xve8rs2ydIyBzOiMB8bV9Ah
DRnovIZwKF97H6xYkkG3jT9CGyTO1mdiaw6XLH7XJ0pYgVYTiX0gGzSaze52P149
DCqhexB8z1594YQIGLVgNnZwl/M/thhc+042ftYtg1j/m8Yarf8IKXIcWIwmBbv4
PgNSdvm9MleartIQWf0r3n3N/4mOgjIzlD1jCGp0ljYUK5kkHOqYIB2v2UKNTRnN
MfTbIKf9mRBv8o119luxrrRwfFsKvJeZzjUe7JoL7P+njB9bMos1YlOClPqkC4rt
dlA3caM+bAjI2Jw2o2QcKiDVz2WWyAIiXtxpzxoMDDk0e8V1xNPtlSKjem9S9JH1
7mSoyY/r/X7MMOEsYg09vig649iWogNlOdecFusWhq/AbWLV60yrvgOALV9pcsTM
BpUusoHFQ7l7EevCilwqPSn6ztCrNjbDIb+LekVfvozFI/P9IWaIZkmlCVL0Owjz
XXXUKbcyqVAqH+gi+jU8vhkXHiHOxpu7KL06OadsYs+yQq+oLFv1/HKckVqD77g8
N0GqkulGzki/zY+G1vnFcrGrtRGxmWZAWGlzD0LBQeO+fSFK3UCOs3WIJ4mUAglP
N18gU9uv720eYSOavG73vWpgBygvx2+PK/tlXHew2flP0ieFovoVqBXTpbCPKcXI
EN9RZ4BtGMpRvA8yy6bTJ2rbb54H2eU5Vo+Fwikz1oco/MAJjN5/jZh9VQwMiFqP
Pqo6gpqjRZABuaijQB3D5rF+qQsKtO7NCMEA4ydcwL5GMunMNaetSl6Fj9q6SXtg
kLPMuGKyHw+uSIQ4odPXYzU5R5/i0WIcBvrl/+Ua862EncawbnGLGK9EntRs5Qqn
zt9d/An/NnvuJYCnKVRZ35yV+l4B8AzIhzBNwDbl+0MXCX+5SCNFYdlUA6osNyNS
uz78boCt9VYwVandso3aJtg8BOQGUFKzsKUUzVhdmF3Yug/9s6J3mVTqeYRI4ffU
w/GwoL11NcpWM7d//mAwUk8N68uMatrFCULalZQkC+obO6hVqtkeeSVVLdIAg6tZ
xigq9KP9+/Yt28xxaHSEDETMpibyyXj0DOTAfUNdCpnGs1qateiA/BJ/qghUvW21
bXGjtWPtX1+nVl7vxCrmaK3eX97M0N4ma0bo2Yo3UYmuq1eeh1ubgOpz0JLTidMY
4BIWA3WHXFOU+sQ53VH1kgxdK0xvylvQ8YaHp8z2MkJZDk31sF1nnOhTjXZICTNz
+pfBR/2xZInZb4wrF18zbwyrM+6isjmjYB/vqSNKzEcW+QUSJ7aaSiAAg8sUzggD
z9nM+09p+pGcDW5H3QplfO/iFRkUJqqnPx9BY1bBEj6ODRt7flrpb8TKq1yzNs0I
0BEXzoFNJsGol9f11CY1SejMREMfSP5sKh9ppmtbUXOs8lJHfyk992Yy8NX/LwuG
FuuqAdvka8r7BZKkToXE85ObJXkfbXJ/IpqE6YbrXyf90372m0W18qPM/fcxD7lB
hXXNqJfufhAgrpEn94FjSDcGsIsjbjR5yFJyIQfDPbjEJ7BDNFdPHSWL8jSFn5VL
uM6CoAzOji3tHxA1UDaX/Gkz5F1t56xlAVu40xG571SgC1OZUsW3OFSZFb4rK4lE
u7BcKLQ0NopEWA4t04C3MSMzG91Rl0t8WGlDb1xC1380xa4iSovPhRB3RrmIjgpf
p5NM6XHbmO0dQPfJ+6nIAzfG/xHE4nwaRyU5KhDECTu9++y221zwpaqkr+q9mYvs
S1dGSO3t/WmC3twzuZvT90yDLrej0g59UC+lm3HunK/vieIX5/ERWs55DX2zcdRT
MR/caVvUnaMbwMY1U6Q2/XR1IFOK+tMpFo95jJ2b/Eg25j0EhimV2pPK37x93r1b
oFtHeu1Ehh42lYQVguPv8Cvh+4n+2uS7axM4Is3rSHo/0htlVxMOxIX2y8JgqW3B
/cL1X6CohuCTnechtfUX8bGtz/XE8G85owOC9PEUFTSqJAZmPNvHbjgwnXQAtVAW
VMx2jm5EgvQzlV1P77bPyz/JbxYk69YqjCyd72JOB1IMDWz+dB8+xMsjBYGyyAwO
UkUkig6YIBCQyx44a49C2Y4R/7dMad1NkeC5TmXk/5jJo71NU+o9H/C0ZRtv0G0y
ajuu9pzSJHtJhYP7XMjps4tI/WUsdyWiln9wmZAtpjP08OCb4Ii8VB2h42Hlb/ai
P8a37YK/HeiOI6JYqIGRVOPNh95uxdnfQgQ28y/0J0cXaZRu89NdRYXUXP7luX9L
RimoP8WUm8upEnmPQbIiwPBvJ7L+Y8ebh4IYdYvhrBpTWM13Fa9hDfZjoWwsQFvW
Avl5rsp+UdD9EHcfphdxsCU0dgZwas+Ll96vmsPEeGiKAL/Zrkue3CyBrw7giMhf
rm/6CsbSx0jYhAkbn+ShjXs3RGMQ7u8gtq2RYnsOH9Uobehb7P8zwRyEAi0eixxy
jbHmRWfe8qZ6PdwBKuErPPKpsc6NLrsbv0U5w6p0iaZE5Zu5g9Tb/waN4r9OXDuL
pAjqi+GhCeO7tHhJiHN0uuM5jxN2Cx/i6+6gotaKduHegKsiUPuG3jLcjk1giP5v
yQNS0xCv2AVUswi4IT+OicalYNQx/3Wc2JoNHUGjhwdjuBV3J37eYq0lfHXpbslg
7SHuweDreJGCmQanWtTaIEnm/kh6I5IBHezxK7VFOQymncL6VlLjFvwCshJQeT9V
DHZQfmQ40IepaghFW1RGUmqLPKyFErDhK3eyYan0UdtmHhdeCkYzb6EyLVB3fce/
97WVSXI2qzLLeCnmo0XURL82KD7qwSMVNPJ6eqF+4+aYikE/U1cV7/+RToJH2roY
mW1HTHrhdONKrt9IaK59K4mzmYupuGnBl5tNO2ctkQdjYayRW4UoeTuVpcEwfTp7
BL6Fsw2ADEUymAFO7wKD+tYD7KZLG3J/iGugaUIfJpiuJ57BzQXB8KEaYQcX7X0v
VM8IsxBiB/LCKOjA7mBuGMgH91fjWIMyQcJa53B0VwR5PPGOQWdOjAWZA1I7c8LF
cW20f65LrdEtmgWLLfUkqWL/QwLiesRzF46+Q0OpVb6j+Oqepsx7+Kp10r00HFnK
PWCcC9nQcbh9Agj/ppZurJgfZNrbFRho/0ZsdV0OjyyldLA2zQB1S10FHSgXXj/y
f0k9QzxSWWZbdQM7jlgg7BAChfStPsvx3QCc7i3NPnuPF3WWc4ggJZt1Dgkw43Wh
CLoKaSx6ksm1x2FiAsmZC4pgGvzkJFGGUKhY7reZVRlv+oDiJORZ0UasaIoeCxL6
zNv8cpzMf5cOXuMNqvky7WY26auM9/sKC/G4mI9mMY7jV251kb7dEc/QoiN4+jkv
M15IzLGL1s39NP357ouVNXXpekLmD62I1Xi700luBP8fedwZ/Z1tAWsjbJzDoanA
3QKpgEYTMgUDL5gcyfQNGzT+8aARZwbpzry60PSa9+2MPwU6wm8y9pH31jZipq3b
7xoRgHzIcGdg26MBYan33q4JlU7SxkzGYivwDIj5ORfIwR/+VF3F5ys2iriIw12K
Vtb2igIp896BnbEwebD/Hl17dLgxT1PViWzpr0sxsqAfLsMygLXSSDhJ4yjKU9hX
+x6cTdLiXZeDCX5tc8puRRrGCS8E7Vq8jE3K1JAqqQZNgILOGj1AtEv3wAMsljF/
ddcSgjid3jT1e+q6JF3Ye5wA1OPwqZ43TV/tDVNfUukLDVmwcLl9DQ5jA12oDHBk
NWyQKDksiLKtnc0NRQvvagjFGhjT08xYK+qTuCxxZmoy1VDZjzwr1i6YXl/a1htn
Pn3XqxMZhowD3vVA0fagoAoTA33zbP5QTBqJ3lybG3OplLwRaPb7OzDxWDp4s9YI
LY/t0NIZnO+tl9Of/NmpU0FyLC4KkHyg381Fu4kcEfW7eDZtpKrCK/NYmJyc7EcV
y20TqkGKRjVbcms3vJc2Z0F4ovCT2vzAJnVZ4wIesJpifHg66noBqRbXEUX32D5Y
kJZTWmU2S2r0js7Q9J08RaJAp/KYyWOqrUIxAE3VmFBXEVCgeR1q+1oCnqHMeW33
l9/DBxqpfspnNhEErtog5RDUJCMwUPfmJXWS7LrCJHNd8YrN0xX2BUGTYd0d6+7R
KXJ/SbUGvhfi7mOev1waX/s/UePm1SuzR53tiIO4BWdLjgqJAaZtE2jufuWarKV+
yfxaPr/1XI1pmOEF5kyZkKQ6wrvBLLbltmVek07tKBsiJE1m4MUlj8KlGheTFWBy
zb1VJrUKxRw/snULjss5VVcGPi6PkloRv/Koltp1OLFVzQqnh9KxsGLDuQZ327YW
fzqXUZvLD+S/M3spt/fdwmessNUsQGzyPtZ/Ew2zfkDo3Zp6dOGTbCo6igmRE7LC
um9S8nLZnLJqRp/Q0afSMsHjAmvfFnsSap7Iz+9ogWGgeY9KU7JMgGrD7mcOdTl6
f3bPEytIgVWMihCg6ET3RaM8LvffoJpUf60oce9Lg9daB75h21rAJeo08Hw6GnSY
BkHGV13blk0t+hw/ATatrF/luStwwyXRQvJw6CSFeWNasc07jNCIvLRHbcyvtazc
da2qftW7WJn6+vpO8LseOa+XAnC9sJ7Xox/K7sh0OLF9rVhOJJFjFfBegrHgFYbS
r7pFifenN75BuKdL5wjKa80c1MiAV3zpyZpTzto4yQGvZOvcfBdSX2yU70r0OTGb
0xD3a5CylLNXfj+PfxSY1CTMCKx+7z4itrqiuK7Yr/Is98fIZ5vVhmtWKxFZH/EA
WZoiweE10G+ho4b2+BZek4nfLtoU7p6Mm38irMWYfOLlG0KEORXiq1dqvkWR/fHB
s7dIHYN0xEYAOtAZTZ09hEckmdfyTJPBZLv//KRb7v+bL/m/wFhPsLSfrsrzVUhD
3wPsZX44wAAo3KLtSVb7PIbs9LdQ2DL03XBFFtyA8uGe4q+DakGwGeoT2a1YOeQ5
O2JQ04d2rufUYg5Uwn5yOGKkd3RV0o0lwRHj/G8D+5jzpOIjqs7xjIX5HJSWNuVH
BuR+aKCBJOww1Qo4JTEB9S/1J/UHWQe2LOjkbQNI5bx0qlXbO2Um1u7V1pxXp9hH
8Hp5Kqv/maSM39GtgrRjnd2K0RCkusZvpK7FXnDFb0cQfsOp5cdNvxF0kBSXYp/7
EIzzYHEGSuDmrDxhKPAKqt4PiBO9jvb5XywiUXUHEi1E8k/nbbAXNXU4+qHUpnvV
Ji1idWE9oHHZ6uZCg5hRs98W0uxS+clKC7GU6XnjKDAVv4NnB2V3uKN3oCHkliDM
x/9PguNRjLo1jIkaCEkDtf3vnyG63QGuYa3Hk5i4Vii2yKaEALw21G4stf+EqgL8
OALWKc41ipCmCd2AaXj9L+4H1me9wbxQmX2q0Fv16/kSjdMraSKAlTqjB1gkxtOF
nJSzSnoGvMHVDB0bXBNq07PdVdRiWKdKq1MOj9y87bQwHHZcnZSI9JK7qjn+mtIx
BdGY2qyYJhNEXKzrO3kYO+aozEDQC7UxeMg0i5jZDFnB3K7WuJ288gjSvcloSJli
wGtuanx/Yme8Nc1SdvcswgW+R+2Ggp4Bsafxzl3DPZTFuBkCptIhAJNDIqc4sj+7
cFYG4/TfZVoPPeNioNjnUgFkxc0NLtSrQQdakU5ky3kiMrFgeVq5ha8AqJEayGKY
mCKVxmR1SKNenQQYohXVtOyjuEEZQj3WneDTYYO2RZL+wiGUSS5LsZ86bCKWkBtp
FjiwzeCjZybQQc68ayQoD1osWJQA3JHPHTIeMl1MtYD3xsXoaOhrUHnv2uKDZLjI
9KlivRT/lf6cMJC2W3j+IcdTucq1zyU+gudtrvS+Gg4vWpEwpAG8V6yDmj4oxP1t
bJXUt3SNuV1MEFN6QkdAbg6nKKf5rI5gLzfzD6W9b7X1NM4NKvjHUGItOtI4f6gb
72ns2EyanWXrKsJwjKGQ7RllZn3O2O5AfyB0C9YcFGR3wJqRZQAjXzE43SDKHNVh
RUNOvOHkTHu2KJvod+KFBvamZl4JbyO8bexyV34s3fzfxayc0gTvIo2CS5a7EP1C
kp1Yl9YzmtsAPWvRp9oyZtNVYlawltG28WxTucE3yfyXYgT1SbUOhScjIAFupUdm
HUTrTrvi5oWI1vIX1ivP52uOJW3Q4+0w3em+9yUYLFN9BXqPGyG/jVDPkRkkOi7W
RDOblnvPGQzMxYCtDjNXty6hx5tNCue8NdgfrD1A1mYguIWwOVJLGgpn7/rLkkNu
RadnrmaTDCKF101w+RqIdLPc/6VWrQiVls6TTJpFiZ/+hHGrAGl12i9P+QHlT+4p
xPG+cKefqIX+Sm0o7tweZXqLh8f/6dYHnKwG8G3/K0XzvLfvXD5t0Al9QddzzG8s
jY8LtcT3OrpnUXhY7V7yRQ42Ba34pegoX4R8DTd6NX0gpTI68IQ6XjDupky+tivS
sjozaDtruY391mU4aRzrL/hZ1OqOtPIzM0PdPhGBBnkELB6CodlYGaRckxsiQM2z
kfr3oGdAMkUa6BeXSi+Lr+NAfFxHeKA+wgkxh2729XmJ/HCOMZQ/mM7DS2kjKnl9
Yp72RM2Gsl7fZDKenRYMcPoc+C89rx34tgBlk+IuuIM34D2b90KlFk6lVmPbFKe8
bqQCVJMMEqdxAf6tEoAkp+8SmJ3SZBBk64xDWYtZTNMZ+UDp8cWRSHo0SWGdif8S
xgEEjFnrsq6f6ifvVJLmV9PJRXEPFhczwxE/eJLLlZJjA52sk2FA6+X2G7dvvW+G
XnPauHU9VIBYOthG2akDgI2fG+hwpmHbixILVgpdmo+th5S/vX86UOHT09ItxJ5E
KuScXQ+c2Wo9Fgj1qrWzvwak0heG1QywVjNeFmBWYgM8eNT2rW4Kf1GSqSlWQco/
cqIOfLHjgRv0z5+Powzzi36Ww7Fe/QJqIibLSJRMK5IEaXZi5JkhTg31nxj5xmBG
hcUv3gzkvyExCvEUp/jS2MsqT0tGg18zH3zPtBAx/sFqJoHCTTP1FSuQtwt0Oy5l
v+oHJqYvQV8LTLwm5mC/aSGkdDNR3Ft4qWZE2dKRu1OTr400Ncffdq5NO2mMKDvp
0KFHGkCrIX63cx81fbGNSSFymUkg2thLcd8rGm7zJZgYO58ibdCZsv6PhFLDoThW
uxS8Qt2ypjyJuGWlYmgK4gKfcsZnc4jOuG4yP2522YxOqbYxTixXEBGvMZSp41tU
6Sa2qwjmNp77kArrRZ9xd3YvWFWkRe3NA1GhfFCIgKI5IGFCjZVTP86Ycva4fSef
KViHycT9uJSq4xNime2yMVvFGC7gnJe3kQCCab1/IoDSak2tc4KiJeg/xIpWgwWj
PMgcc0aWzE3K7dMDJ75lERZ0mcjeJmGEONOfQif15RLDjc4SHlMo43lnikaqLaFA
/oGtDynXi9bdC8po6gDFFZ3NIHapWeoSYJhdo0o2WseVUVOGdgsCTh+l412vvOBB
e0U9AFwAoxdmvJMyELzOYKyl8fJ1WPHpvSAgUlqsIWz3+3VkvLqXLR71stOsERST
HxaApbd8Ssr6BFimFE+XRjYbtjrT9HsQA29G8sfE1sFjkRGk7KlvD2C158XqYLSJ
r9XVXTjD3+LLxBqg7Bua9mHMwzyYryhFVLTQq2skPKjxJlHUwaOA/c5YEOUkHmsW
Crfdm+88RN1R6FX+x1MhNWGBgdksQ3uJta4TaB5QjDrkRM4lGVmZuLelm5YIZahc
CruJUxx/T8/TRP1HUMiMbp8G4lkF0Xd9QHg27bW9sffDlfeR+2Pzg+PPhdrNcd+M
v7gxr6ATiHSPTaQYqwtSa5qmk8//DFbEpBBIXlW4Kpa7/EBECxEuslCxxaRn0dvR
foyrKM6z4Lx998z1toyNWxL0Yw+mQXZ+PqdbM3NsjZCn5MlQmUYr8oBQM2rhr3vh
w7MdHpyC049tIEO3M0DYsviN6JNaIYb8Evgrnuf0dy03vSBsXlNlxGNd4guD536a
Nlqb81A6Nqmx8OTqCCkmTn8zpILqXn/nkeAk518S8pFuKwbeMbRfC3bwSbKGOyBN
nve+XBmbWDHjVMWdtUc5GDA149pBq1nISBsou0RHgJtTv2iStgyAuTadd34M2Q1q
zocBRDddJcPi4Dh4HnCFxeb8Z8N21+Y0dzj19vhtV7n+Z2dWhYI6I3XlBm+Ls3Kh
ZrZ1WAL4i+iUA8NQ+ePcLY8ZA/0k8V24jowI4EmTnmcikJSwm/DSY78jlUJTdyRc
Ew7K0zSMKNesAtHGMc3miWI7uZTIVnNd6FPb1wmOjekH3oifkmBP5JfhMHxy3GOO
jBt704cx5pSy/TKf6IOCwfP75ffRSH3GdRHluxCtPQydrs2/z4nWP4Q8JWrafAxD
7zfgvBOgRC+R2HTOrnSl4uNxj5nliyE4Mk7MWpHfCrPWxghiR0Ob6+syYS2EioQ3
aY/lU6nYfIuJswvBETMmKo828LI2TSpKNNsFDoGbWZ0fejuiTFRjqzvrI9dNzqUv
ueGKf8oS1Rg22wDQyMAZbWalQ+evCC/CZ4Y/xb0E5KQE1D1ijDdFm/hXHpeT0v7W
7yvubDxGYtOLS4GN3X0Pi+IY2y3oOu3pZ1Vqe6IKgXSezD4YfYDzQKZW786aDeaP
f5FYcHlCxf4PYgQLbJtwtKt1S1g41v3uuPFGF4TshdRfR7LCNR5iZJycD18hkqfu
+0BQVgJmB0YTOqnPhcTTh7cfl+eovgjHZqZKkJIn5xwfnawlyea5PdFvRf2yEJwF
21ZJNeAbYefyowLlfdktDxzTf51eKFbmBY5M5f7CUEqITuivYSYb3hf4lNNDeqIK
FZP86IyJiXv9GUx9MXBHsOAs5ut/NU9ee/vByeoeYAg1KG+WHSHpx+QUCE4ob5UW
k62dLasa2fjVtQ1ytiDag8M78l8V/kCQgfPxyv3kH6gOOxrQ7CKSbuy9FiVzZv5e
oEfxlmreZsyZXCT3jD2nlF35GiUMCNetAqDf7Le3TG/br8FrqwbiHOsyDwtZPGwZ
c8z7jcCOpnlKJsiR53P1vlXpr+pnoZ5WecCOOCejs+Pb7bFRHDfo7MfCk6gY+NJq
ty0gc9tt/IjpBYCGdjMkZt2VCtmyNzJaJKWwthvYV4iG7zjP0HbZJ8QckJ4EzN37
YBjbuor3/nnJyMYbW79X3gzpm6VLOYOuXo36+tBJuw8mXHv1meM3LG9SWOjeJJ7S
dkrMum0mTwi+1z9bBL07IzAD5SfGZGp+dTDB10ZHi2Tf2EP1gBIHR8OQ6NntNwIL
bxSsWwrSyHFjOt/l3pSbV9mrRBAwsovGE50p7DhnNXD/CxvnhL0AjyNzPmBRYV6y
BNN4QLYrKVQztub2TmuaDrMuyprW+iHkleCSRW+7gMMQxRT7mNMXUwCfK4pFdcQ7
vXjzUo7rtbd39HVQyaYqH6BNG0Ge0BgTkZscGXoBLHz2/7qQXZB37FU0b6T6FoJa
GkH6r8j3rjPzxNEwk3E9hSJfIEmAy2xv1lsSYKyla3kceczXl+lzyJnWmEUxXJce
FlneeoI8+yirh9VlqJUN+vMY3zLNfruUGjMsQGBRh/ibpcJChpTna5bWAQlEsepz
5cvRTy1m5K1dqnWqRQmd9U+8aaur065EaW7ZP/86LmUPd2NuGMxVCUHA2ZzqGEvI
SWWTwG6lAFJXT4b+X+p1abv93kqfLkrYlGNvh/Jcqh/jkaGgoPUTyMiwy4ezLOVG
3xyVq2Xln1V6PSZtIAeFpVYjZrBZu2YZbwjzhN7LkUd28nMFvaYAjVWF+fukO506
yy9iGLb7HF+3x/CStlCH3TQnCF8+1XMvTqLz5zhRIucs85D7YETuSOtabLKODP/I
nOsQW0egTbPZHlPxZf+5Atba/n6KTwO6n2g8i7jMTXhFL5TCIlU7WUbS3bTstzRH
KftsZnKhOEYtLusA1DSeF/egXzJqgKXMwZyyRu6tuvahreUHgaAfgjCmh0CyEbd+
9BeqF+g6WlX7cEHWNAIbKbgm5QVN2inaJ25sc1xHv21B27E15Zz2HXrvq5QoywN6
fYIKFMOWHKkYc5e4iMQ2s45cNvj9GjLLQ+O+h8Dz9hglTw2pSiqM3+xO/f3LUDIv
2YFvaTQojG0gdwS8eM9YoFz+wTp/DRYNpQQ6NqXiRyACuCu2Ih9W6IbsynAl5piW
PuNFXoj1TPHiIQhmMtieJPGRVLpmCfNQ9GJl9NIjg4p+7K9Zt6EVNZOK/kbu3mb8
v1Sr1ZkdeZ12ZWtAqMdNzHLQmgTYyPWv554d5ln/2nguYbF+xmwpyLySmyZYrbGX
LF6Me75IV8eUf5ro3i2ph0XtGfTELt7qmeOktb6P+fs23zbkUwjzOccqbHUyGJWc
m25pWcywFY/mFRA73n1230kK15/zwAaKr1LXNCstNXN45FmsMLotRMFBDL5eElOb
3rPK4bHos+eIwMQAgCIMgaol3r+oKmrgdwtXhAB/AMzu11S0OcwcVs6ub+P42QD7
WblsHMagf1i86q1nvpcvEixX0HM9LdKBerQB13b/+xZpM3+IfVpNbhOFKAOvD1ZK
aE1eyHATTBLI30IsUu1ulsF6+xLYwc5ADTBxciM/mjpQ02uuiWXU8bF2C8uw9RNz
slhECllSKoBinLbKvDzaB+NCUsHWZLZqTuTM5dax1R+y5DLECMgMAbA7PyRIGxE8
TkTYWclBcxyuRc03o5N07MqzOdiyUG6k+J8o1FebQoliAqbyDAqEPbB8j0HvYeWo
HfD3INFlahlby2lBLO3oZDtpQNr/1/jeaCZgd2sJT0Tf1BzqiOjiYHJ2Uq6LZ5Hl
HSjyZ84K1QQUghR72ce3meHVSJ/CX0mpS92YUAd08LmXrfgiPjBLeKbC5aGmoKX2
awky5i6qZ0YMu/fvuy8mWsMO0Uznn6rzp0LE0zXhKUZ1fqQuFfAadSoYFt4Ul3KY
eGmO1M3Kt/RGaSyqMtDKE8N+WAxLZFrmowh6yfz8Dabd236Eo+6SDvnyLtqMFrYV
Jxico9SswCwWR25llV+5X14pvSZTwe/nQI+5cNHohNz8RurXfjPzsCsstUbMhxB6
OKb1X5mQj8u7C6lgZi0DSE9iRgqfa3eLYUeGPhBvD//KALWgzNNIuv42CFMiS0uA
S2br+gFj6c+o0MbqxXpDKfBN/e1F/Z6YIyiE6eANyMLLMFTpsOW1+RykuxRNxZ6Q
Q28f8VUN20/G5BmsMEQAjy6Qg5ZCLKP2Ben8iYNOfUZzR504oEAkt0hAp0FrGS+K
zT8Zy/BaGgHHDBAYLTYV//PCMsNUGCWMFit7jtBhFYqTfIglq3eMdrgVLKAv2BmW
EiSxHnB/nmZ2Z49ZmeOcoz/iCDV+UPkrmrWWQU8kAWDmSGueWZBieYapVezSWgms
sf6rKx9yBFgm4+S8n4KDv2fHScftnPN1pwtaBVmUcK28Vo5FGR+P0PchkfI7sVbk
fDLFPKN9YVmOTxxZDdSeN8cb0OaO0Mpkb646u7FGHMFQe9FmIKgAAggpV4h6PRxK
oPaDFwFeSonKVMbejKw88CjjE+h4aFx+yJJGv3SMUV0gd+bzP+HgB6sOQ4j5DyaG
7kiVibeZ9bWQkdzvXgJAr0CMSevCkLf9xPcJeDeK+0cmkoM4n6pdLnI5bZfgP5WR
9xFCXmqvChu08jMwmA6ASLV1Du5WdMI4BjPvWrZ9AlWfuj3IQ6JyZvcaCydZFyTX
lEXZQDyI3MM0l9dvPYwk5sveSv6oWYRCQbF7geKvV+nElSkv9YUZxjjIRkuh6u9N
c+jNcH7ZhoRUxTjO4GP0sO9MWwdhUQ0xrynA2dLqj5Z1sipPCXOTUNGXkJgL5bKA
abOE6XQnN7xua9AexHPg9Exh1RZu6lo7afKCL/P46qzZJtI/+gS+RdQ1YxS+xxip
FLVzujNMT3fRhjMNmrgUSLNgS5KwyA1GQS7rkKb8QwxOa0qNZNmYOAXMQnNTM3CH
msLImyv2gZ84IKol0HYtXEQCvL5CrisYGb+tRTogapO2gGLoOi4X8Or0dHPrHqR3
fAcQsgWGWkZP9f2JErdBGebHtaxvGDDZi9wG0U9UY60yJ6fw4SlhqAJBzchkTmPp
fYoWLmpZBgKIgZimCx1WyHlLzIjCCnLvxHzCk8f4T0JVhZNEdi1iGLon/+9It2Wy
Z/B4L46kAEgVH9R8zpY33DTnX3VzBKyOHMeLKINkVZqB5bN/lede35OhIXWYEx5F
Od96cAoFIjCM4pjxXtwIo/d7IxJdsh6gTsjmGHE06pod7T6lUAv4Rn+vtTRwrxDx
oagZ1FbqeB4oCcSLVDmeuyK/8V6UznBK1JoYBmJpaJROuS3E4q0+AFNJShB1CNww
CsfS3rtI+CUAQ54lDoPLRCPemjqVwJtMkDyuCyj+2lHeT1sozVdEyUZ/4YjyrTtM
zSKIV1qzbPtEiSEjfnVMXc6ObxT2kMbbZc1+oBujWarHSvjc1/ztR3tiTdD5vNJP
FzbUSHMHyovV/l+5uAx8p9vNFLMbU9pMEdpsu9fId5TH8Wjj57cueILX4JK8e57L
UAB5Q6kg2lmnat2/JqigFEdaHka/JGn6+pnjE5AbBuOSq6SVEYvKnHknKIa2MmbV
Oy6bdptlZll3ZgSVUFYXpdJmySdyq7L6zZHIttgeDZ7CZprfTAhDLkL2/9Zh/0Ui
KI5tUkhWb+tVggoibfnYqrhrW7T8NPLpGq7z2djbn/rRwB2Zl/lLtRRT2wX1B4yf
uOmv9vMCWkDsnYB0zkGGtcvLrFrZXiFhthGHFUbNtkWU5DS+8qQ62ZOIAInblY42
i1VhenFAhQoXJ8y0NU4ii6we646ELzhUbyTI6lChCrsHS2IS7FZE7XU33kH6wzct
OkUMMTsdwGg2UcBeSv5wQU8iJDVfkBVFoVswUB8wCwD9Xg2LIJcG7MxKylnXm+Gs
McAzUE/1ZFZ3Ygjh5bqtm/xJOVGG0GUmkx4g3uPnG9+jrtlBbJa2eStzq2xJTIjm
HI5UE0DJoMd10EEDlKeu6iUIknSnfSNo41rfmHo3ckt84is2yNaxkNjEQzNBYvGg
Ca28ewvqqxgLovumhT4dQdYY46xDRfLtg8rNJVMUxbNlxZ12GahK6vgQ0Yqe99/D
WGaIAT5B0UMhh9z6hl+zFIXnAl4H3xWRL+QmXXTO0IOnw++wIYBT2A6GOU0DKHXx
iHVMwOGRRb+mNcfD2xwsbZk5KMG+NVYUcXEGt8U96v3h/ZGn+OG1ixPxpAWbcPQ5
qbxST2n2phdDYoCPoW6fZShv8W9ZG403wTp4eVTMJ3YkJGeiEp4LCMkCzyFMGQ+6
PjLwzwH33D0hkcOyi7fxHN1YVsoYqYyPwDlsQqB9FyvaQ42QLKa12vPtZstwGVeJ
+7giw2Yk0sST0tKG+u+jveQ74LnMwocETBRYSdNEy8APs+BM+VtqNXKuw71/5kta
1I+jKEJkBBbr4ev5yIoQcZYKYgcJNMLh+9vF0Pe9tgaRwzw2CL/QUlcf8CeuHnle
bIUkS5TBjbo87Gi0qTY/vz6sbRlBaZLaPK6wtyCEdmB7wbsdkf9AIoC+IyNxGrYy
l2OrNh8xvQ6txD7X2M+wdFc69rLa6zpzAwpEALoL0EuBDYEV4A2D+65YOnvXneDH
NsmsI0+n7auoeZOyA0mOcknyYQil+RBZRSL/3lCkB8VQIGGnJYcWiAk0ffNLSrST
qK1Gckt0D/+p2wQ4d8UpzWYV928tPRNvKCoHFr+D6GI6bxyiAd3YnFFzC4LR9b1T
H4jp/0LGeBtHg/BLu9wSHHFL5JbuQEMWMLC2XHdk3K0Hva55RYDeXpX1lIT4GFUX
q51N5ECFPWYs/YBFEYTGV3VQfw98Au04HBvPSm8yrkIdl6dN2IB3KfIuJX8xkIz9
IfwMIo1mSiP+SGpqgCXnLsJUOUAyXCqTlErfU0HYnw2FDQbkxn+rw9bbYacDKObD
kbe4MzEGs7z4ttLyfRir9um9jbuL8XPetQ0bq8nDog6HK4D4LvnWleuvyijlxzmx
QUwJC7ZFXmsTyuGuUOXuYBuJ2BcRMW+rd58tilmcORAhdEBwCZiksxPcXNbywkDK
vE9sd4lwnNxiu2lC6iQaGJeH2iTDUg8KFcfjxpvdTT2DIKZ7Ofg0wJ5feNWg3a7H
TnIO65JydcBL2IpHqyB21jPsnnrypE74EWfFeP1Rl5ZAxc6f/b3rdt0LdDKpaINU
pSUv5SKP9F/HNeD4L3xwc1TQEtaColQ6xHqFzhCdHjZnDxnEvVxYlblp2vhuLp3s
Fx9ujqJCYdjso31IxB+LCN+dDgQx1aUWhQ+jQGAi6SF0a7wKBCiEtYnO241I3pUM
ptnrWckq12I9/O001RTgEF0Bq7ANHncZqp5bg1vEd+PNs3ZSxMMfkB6ThDNqTarH
dAMPN9KhVpzbtjajxwgkY58rz2AM+NXSFFgpWRoFtMJZdvkS5oDwOrkNYtRVR7gg
LVUJOrXysTSV0yk8NqP4GIylqj7k3G8N/L6zhSw8vDbuLs+6Os7LGI9L0S6mfu15
KZ0vyku5aL8WI/Wd3SWZ+xD78AoENHo2NvFbyroqnRZDMPPRLRa/27rFYCGfZITh
uXUv/ztGz44NADUfYYUoVXVEKB1CtGuNurnJtYuZBtNJ1exJ7ElJVOY7ZDjaDDIE
EcNn4kT8vzKaUTK37pK8K/U3kro+AWlHuVf22bRQJ3O0cPcyXW/6Xcv0nySYqkCw
CPL5kC/Ao+jwjg0/o+P7bJMHAxEcjohBLLR0ym4vlUnG5vxG7oftu5uRTqpLBUUA
a98rsf0ji34Vmsu45kyhDHP3QvDmfcGvirtlVgqXkHdmTehfi2qPitn9pgM06U2d
QmGbboiUc3WP4REEX8G9xMFf9ZHwnVuhhjWnKSGiqzenbnA9k6Lep8xJudWtcYUj
sqwrAOo+BujCQ5neW+4EZmLa0OWBmDKmYPUd1lY6wgYMD8bth3FNv+s1qrAT370U
fK7iIMKAB6Rn4BRjyuFEHrTi4vCyXzE2z1qERYtE6rTQfrd7cO8U2qBWeRE6ezik
m6tbxHnd5sBVuKBuPpo/GaRBYbifOjbNEGub5vfoj7LCnQFBXhnuYmUo1jxRi6nK
WFwWigSXqnEEhSrBnqy675Gjqwy4hyevyNaunEBNobuucWSSahn0mU7bMr2ZaD74
LttMT9qiZOzcx+3TKCbjw7lQQYl5zl9lvANxISK492BjWH9GI2j+DiUbQm6fUxX1
LOilrz3U+a5PZDz3BTW+K2V+IX0wNXU/bwx82NCHq0SeWoBjv0tbIA/aBulglLkL
DDX5w1gRyrZcEqmlD8g3QpX2C2NX9FCXQVwK3h22RtCAfWR8URwoz4JVKvcmeYW1
/o2SSWGAKmePGJqGUJ8557Ra9cWFqvfmG5uK0uQ9tQ5UWp2uCo+PTeH1RIaj3xU8
x/Cr2eo7x2majSw7X65aaIAJViPaGxt9S7nr+o9fP+s6RF3xUnfrB3MpfVRh6Soa
FU9JN2ynPv4RDmB5zS1iC/5KfdOsDIfgtMIRL2SqwXfmXApJA/PIY6uZNB7EbWVc
HbB3/GknBrS/0xhZQl3oDvZuYgn1xaoyvwb1o2kQCh1Au53i4u0skKTup+YSnBHh
GgR93E7gJ2mcCRzaP1iwFsGUjpxAkK6ydVxHITWGjPKLqqFNXpXNYHLneq+buIje
mUZiMFFfExWrNtfRw3+6uD5w/12vMd7bDhbQQblE3jY3pvRuSVTbemZFilJQ5YQ2
arQc1+FJPOFjvUya02pD7rGl/e7PghbxR/0b5kK333Ca9zwvTbpiO2AuIU900vDg
yfTSC/CRXffeELfcVsiZjYkDeZfiF9MJOj8jMF6lkTaSlGVwD3117rgn0JyXvKle
3LqM0CRoje8qbQc3iuno60r/Un19IgNUSY3jR7SDuZ4OTojhBcbzbAMIFzMzjkK/
IoxWTa9hVOJW+JE9tNI/sBC/F30I2vgmnMgOIXltg0Y4JcbvhOhOseqCJkT4rcCe
GQlx/6GZd7/hyqvX5cT+M7t8p+pfeGOvWYoaE1ojogo4PHkPh+NXOifayeO5qQh1
VKW7Tof4bu3kzmHPhp3B13ocHBKPdNmnCtXASvyEtScswJTt6JE1VFuHjRJZE3Go
RssxRxQ4aQlWYlFrAC0b/N55gFqeqDOWnyFQzYymtu+ovO0mu9Ylha7+wJcqpO05
tbaSAxm8oP0tWsYMYXrPVaipnuZT3NEViGqe7GMGW8xIoeoZbWwe8KM1lDQCTmLw
chvf0MmRUXZwlvPCppLuqq3Sfe1L7ijtpF8N9G6+sTvbRwypGmxeX8Eb2C4Gd5Rr
DbrHqatkn0CAywraMtQvA1KA39+Mk8g8G9RCk+22uC1EGtmwvR0en6T76XOEYllz
DMGSnxIyqnJDaB17yu4zUr2oYgjjguNig8NYTew9/K+0aulL58QSSZTBlqtv8nQ6
yvpz22KgDTTrfNC+HZUW2Pl5BhToQOaItGcLCNaXIJFS0pGamVxnCenvfx+whaYn
hR/wSIKvhr7aTwuo8iyH1MHIjxNRVB3nYs7q12qv1z0FJIQBuSVCuKxhHA6xLFdS
tecqZTPY+wiJWUl+qWILDYRCuip5jK+MFh+oZ43etL9C3e5N08tbM+PJmfttcHox
N7ml1FrQq9YTcZD0V5eHuQe6mWJzo2j1wv5uawJkScihIgfO50KV+LcxtY1aR2Fy
KA6Y1hhh7Al7iyXKbRVxyOe/jaQ0R2xlPTNKCRFnefl6hYkun5J3fu+o2P/zoyVx
hFrCLSZy3xAbEFzdUdYbSdwAriJB5vAmUI5MLq7KWRRQRoh26Xqa49jOe5qVV08a
UPDik/9sHC4eyYmoh6DwlOZN0Les3irehcu0sfAvU/mqf92dfumkCBk9HsvrPFRg
OcQnD2jYHENZS1yM3SNYJHNLRFOXATIytfijtaeLkR3fdHXAabpj0GvwpBYygtPE
r9TS7O8FG+4TsSptscZ4ehG4orIgfAXEFzqHtd1qTqziKsEphBFEQKcm82Hl54lJ
233iBgAAe3MdgXJt4Mb0MdvPJGMt8ix/7HaQ6qwBS6aLfpPBf19DLV9NitywCpFg
7m7H+5GvvaYR/CTnz3PgOdlV2UB/Mg8SH7jThbFTO3gcOpADb/i7jP8xa5imp068
eqr9h0Nm/yO4TjgPvENyQ7EpSGzVvHpm2B7uwRNV2BJRmgTTO6rn88tw7aPaQCiO
mUUdGq7whAQjtdXGtfvjLtGVH3Nl11tn09oR53MSOSLYolemnV2FOVoJpLWj6XeK
z66RhTyeYGSUC09x9x47x1YiUpSEQrLowZof6bi2JjcK9JqzTtbPbprbBH5Xo4KP
uZec3Xfar6APgzRU3vKjT3phZP2LedzHlksfQ8v0bkU493vyyi5Z4FFdKcCcyzmb
o6X31h3hJMZRblUEPtv7oUw+Fe1AoTGtnaPduSZsJUBUG+0tC2oP5kR+RBR4+vmc
6iPIR0MyWsRgQ1YGIE57LBqGdg6jfNRRBOVq+eGsLcuQfxBCE9eJjVZ8kwxz2hYw
pJWYMfJZGlcZs84MtSH24eZOrCpAqNTvvG/+8qQYgBVQO+MoreMK7bvoESwSazFp
k2mDS/C095j13DBJeD8maONqaVF2Z9Ugw+497mAXiZpSj4N2FXtKBzNcIhVmZ27M
ES/n/oULAREjYAD8i3Mmb5JLldBs9CXxbZXDr92DmtcBpo4VaxZoviPSrXw2mEkx
f4BcVGc5xbkFPA0VqdQsFBqHe3vcEehDA+6aHMkdtxKLbF0nXch274hIiDZntTUH
1XZJLkhKmMfzKi/Ug6NU0fBxMZUMtPn48FnaSi+nl6FE8jS0LX8Sv0fYwTEnAyka
TBEhLb05ZsMOANmZNq+qLOeuHLMAn9qC95uYup30j5+I4xIXc3pBCnbGHuWSi8UG
uJ//g8a/WQ2GCqvjbxOnVbcvq4zcrbVxab6wr4DR7AGFxX9dBdIJdL8TcyBGXBfh
5aJE/ID8zXJWy3HztzWo3+bw9gqeXLI2Qoms6UoT1P3t9qeIEYJZXDUnhyiunZpo
nuYyqPSEnPWY0R+Xuctiv0LHZwbu7tY5htdtP3D4HBe7PepHrO31lmttcz2J1Q34
Qau3tzVSsmM4POyTozEgWUQokQ72tJnmzl0GSMbMiD80lU06+Sjds3ZVp0N6V3/G
FjnrhIchCKsI3auXD8UFt/EVtXSvXBPBwOsbuus7Y58lZbsS2h4UW27NOAVslAN8
whzWeqT7IMkVblwkUFoYP6MN6k6P+dC59eE5F6pUBhTl+KXgePsmeojDl8awLsU6
MMWXWLxb2XaQb2JhDzqJyV0Yr7tLYcRe96fCWvyEptJ14kz9pKgiMJFc/XUhaiyP
Efg93e/xH7ert9tOtpGEwIL6aI306PwUZZu7PtEBW7/NdQv5m7ASyWchdKLJfze5
6NwJ78LwLuzqxlVmFHJ4YyqPdTc7aaUFhe+8PuLOeDslPBto8Wfi/kk409Y2VFDe
QyUXikEa5I/ThieCruUgxeUk7HaIEdyLNoYj9Z0Auooh7qY9y2eg9hv3FBOi1fNa
9GM5gK+rM3QOEv4/zccLtG8b8RkKpxQLQqdXhnScsV5K71cGP9EQMLIoRBdPyHa0
JMm+5Ny4u1qgbnj7RZHUowvvMkSgJsAanFYhk1E1f/dASr8uhzGBwqrf/saARJQc
1dA1VXQ/QInuYXQ+uV+FgKDtm32GDeeG5ar4qqDIupc3lOem6GkTVgNapJ+BJo7/
ogVKOw3G1f00poVz/C3STOcv6ATaLEUVCEu+dmQLqjnsZA6y0HrWB6prLYPDZGQr
R0YngxNnHTDyzvR9DnOWCY8wZ9uX7rzoYRqBYvMkEqKpPtmQF6uGi23NETaymoXu
JVZA86Vo/edCEP9ruKTxd71tmIhcvCAocnq97utrbV3/kd9MfK2okK6jXIbDZYfh
sbrm95TG/9r0lZgVm213E/3ZvpXkLMwGOhBRHYrPEFDm5yRRn04BJV6Pu00WsF1C
k5F5WQKiOVHw6K3acqvsiyh9123ib7CtQWiQ0QJMj2ePnd97LrLUvLNb2DNwEuLE
3NZxqX535S8CuxqAaT/w5GgnGFbshEoNrKUQhDeziSpDp0LIApN19zHtVcGazybI
1sb1ze1QbU2yGHZNoLa32qSbsGiyOHvodLfeUXivsNr4g2kPy+ZOW23cOWHmXi4m
/ItyYt7oVVx2m/HBmVni4jfWJxIP8gSarMJEagddnc3VaL5fNjJB+pnxdsLp4Dss
t22unHIH47wtxwLH7u8kdec9o5I0g35DykT9Bn5tBRoe7PLTHPENTSeSkbJ9QrcT
OQvB0yQ1EnVe8SFW3qdK3FOOC9gAVP39K56W7KYK02JH6AvEAbMwb+69QZ9ITmT3
AmpVb7/2eJX8JjwUOS/Ia3GQOgCG5wwQXmaLZ4zoX4shXHIXiy4IsYncfqiNwuN3
iyn59u7OE9JwGu1Ks/XySw97rgSx5KK+9Qs8kZEgvkyyYFaGsirFqkhd5CtsRI6q
NYsDCh+Cw3wUmIjWpKi1R98QEXv3NBHRm4Tpado7hGjz72jjIRHFW08kK4UdttHw
B2xE+emm9vuz+GTrv3si5ov9MsfToFYTn25msJ0viZsmJ9lqV8xsJE7c/jnoXsoR
1mpMSgfCeJZawXp+f9au6zG+k0YpYhvrL3el+bWOm0Pz1Py+4lwtG/fUAM9v43gn
TcTlpjnpZ56FNXYZmWWujIB7VTOIAtOUfNvn26EDwocNZLJikGMSyCsdQSNAL8hQ
Sh7uXMdM0DNI3JHzQs1f/ojZZ402Ff1USqaKU3dqTJFFhbAe7o682CNQkxanNSNq
jhR5I+aHQQ3KLXBTNgEqWdh9bQ+jmLLZLY3Lq1wKkpi0Ep0/k84Zla562UtFDRgr
b4gwyJn5NkZhWZS6KJj3MVZmcPqzQFNevLWYq9+PWFWMIu6nGpaDp1c5iw26cp3l
T5LdhNpQjLG9qd4k8naR/VNubC2DrgG4Ky8r3lHqS9cbQZwbdDCPGWBj7AD1z9Q5
23QWdWg2K2S4f/KmFkACM+dWVecLWWCkDV2L36pagxiPWBP27PofV/zpVcJYHlZE
WcsNOXiofuZTS3/TJTyfyXBZB0SrXjdNGqOqRcVlf2ul6mvE+hfGKCCg0c8XtxrT
jepnnjVwPzfisrDbhbhrAkPtGyShzFKyCuOh9zqHSW68Fx7a5xCggVYz3ZbY7u6s
CjLBrnk98DNDMsA8q6R+lIA8Y+Bxb9A+M8Au90hDHEaww0SuhZhNdE5NZjRp42Gm
EAUMGwog0JYTpIY2XJ6rlWd2hk1JlkO9ExZPDu1wj+eL1ErGZCbncc6kTGjVkyai
4wHYceV8lN8ghIgwAh3C9xnBWXRn69gMcQrxROv9Y0sU8aq2ponvaXTsrruci4xU
zAiVibSe6A63RRDMg+RwHHJV5ubTSDZ6pT+ezNqGvX5b5BOnKqLLfdH5E8oWOmhm
pD6yU1G1x3d1+FT8/raAhZvbke7lSWcuh/15TE9eHBemW376DaB0Hxr0vbhAaJMU
0MeXwsyBk3a7z4D8xLTfgEIpwnh2JlOqpSbN6oiCb0vAGBFfhNq71rXvvOhJUqRo
esYk1mFvSVQSllxmB7jXrUkESNMar0jM7jDFywZ6i6fXJpUGwMpIpKBnDly14aeZ
xeIDjmuJ5cQJ18+S1wCLfZy7a8fKoYFfizRy7bb5e6osQZYUCLIyfIHPdNRgMxr0
yz2q1P4CSfJ5vOPJnatNbhbnvjaFuqBjXblVVk02ZxgzWBfCg/HO9AMfuO4f5Ena
s60sDQtZWANrB1ZDlrjqga++aV3+E3Ha2sgRbUf7ZdadsRnnlHuorg+gRYIuZB+4
PHZkRfn6IcY0syT53rRApk6DcQp2teC/AYgeR4jmPLoCZ6lJADtZvxBIVnh66VX/
OPlzw05CxEk6DafMU3NK0hZqjUZrLW1YweEqTYjWpvhQlUdF3wbqb2Lx9IfPd2ny
Q9LOeE0/vBH4434xuHaSpvB7VfJiUfWxL6x2dVYc/F+Hb2xATfuSoQuiMXYH9yn8
ODmDtZQfdePuHaaaKOVU7HIHc0NKUBovYiQHaJnFg5cn2lULB8Qabhj5w5jibXzC
mM3jJ4lRAaVNifDRc0DW1L7KzcaOZNa8t0TC2NBscezWT2HCn1E0YAejjGpe1PTv
zwxVRDRqI/kh7cSYHUhIxozceW5YV4l9UcdrJsyv3yB5hzunhuKP2pcdUtN7nhNK
7KKz9mBf/kfw06bGdu3XWej5NPcc6YPbQlMC+BXYvMbUINbwv68QOqdCGkML0iNa
06YQyMPA5fyMAXWYiOhPcl/cSkKw/dA82bk/I7IrmMW1Q5DanIp7kWmjapMYF2xJ
50nIre+Q3frwWA/2bY6LfoTAYbwap5qznvuU7BNdUbKFTPD4BZIhLvlFFBgDYz83
MS6U5EOPmsbn9nvq/M2MjgNaWTTuH7hVJ5wt2FKW6LplSSPpRrRJSIvB+/6oe+gd
+BnEmt5pcw0iAa99kn2nxfoT5TKOMoHPBof7TeGEERgMOHHmPfTUVr2EuhOt71Ua
4/h3uVFZ0WRZSJ7vHfmhLovfFBFxbtr5v4Pi/bfrPaduOzBIosMwTe1rRpFD8ggH
dW/sjxjJr0cQCzplL1qJviEFfCf4lr/Ymovg8zoUhw6/G4d5PcdwjgUWrCKt52Qm
4nhClnhaujMaYiHOqE4EEqjdZQO0wn6BYGrzHMasV9rtMnbnNGjmeB4s9Si9Nh3E
npcNNY56QOMMD5isGV24LmRDXZx9IDE/a5+B7lJ0mIRMw/lM/k1J411AG0doi8yX
p5rZA4znmNhiayqHDNgQqxfK7WodTZ1k8Rk1OKBbRv37i/Cyyxa8HDddxW7HJNnN
V+ljd0yKgrydQZY1OgLsj0LGk+i4t+RW8wEiub9Vnh4ocgG6kb/iJRH1QqJuoTtO
eTL/tNCA7kcOrJShiNW5uhcdlB8TE9S8kr0QgTakoPt8kMVTmaVOJ7R/EhGZBuoR
/5AaR5i6hqPKxLHohQY4C0a4dAU/CJQfdng1cvFyP/C+k95zTxpjat44zhICRj8f
AMQSanMNEuru5CXpdn3mrPDYCQeyGTzICWmYRfmhmwVwqJ04nXaMxURAiT6pOBkS
SszWH9GVbUiD3MzHxPO1I+Fz8JJ0cfJqQKaJKt5uI/M8RmXZG26wq0gssqFt6k7C
CgfG0e0pmMmnq+vLyqTDG48EBwzFwC1/hwlPBfXIXhti6LJEqRlef/GWGBMI2v/m
9ibKw4fqSRfcmuoNzFooICBSn9xelTFXmpI6GWNuNIesnYREI1uhN9EaEkxjIuR5
vuPd4KhLLZN6j9hkteIDdNbNzJEif5oL0yAdjvoywUU/YUZOVmJgtXxy8cdBM4wv
/FNaOYp6G9osG+rrcSXcTRvnNUEAWvjO1K1me5UMR2RxlA27e8xP4VwdrHscic3p
eSpz98E8PHmvSkS8eXA8BgNcXB/zTtEKx1xJ1o7PzJxPxXQHMR7dpA0qkraEyLg+
AY02ZOdU9N73/i8Y5v//lGyG+YF62QsbpI4DOIPWzSIQD9ioDIpWpgfXXbiU9Bhd
yKQSKmNLNHvB6LeeqKWvVLvMT1GyLdqpwWtUe1UN+gV0NaEbUg6XnCb+Hh9g0a64
1DTcFVcx08g8DZDjAKMHAsYxQGzIXYBziKx4UvRxxI5CZFuJTonTl4erbYM0+pzf
IaX8ZOqktqtmqvGTSsadbZgHd4DJ7t9A3eP2DmoCNSAvj8J6okrx3IGJWIugPnWQ
CdEtn/s9DUgeouIMxdiLENo0jsWwWF3x/EfdzR+klu0iVzEC1FIQeGoORB+iBRGA
rAgrhuR/UhC/e8KtlUKMritGltFYBMokRuUqmy66xmgzFcGamlUTylHhBzXc+FMf
MYRC97i/l2IAlPcHH3g+ifGoSlhzOruShSBAitMBu90SGmBZJ727hA0I9eivERnR
ay7xrqmNgeTCzVpKvKN6xin+b63nDJhG2JoT7+oUgsjiTmLoxBsJ1QrRZh7Bkriv
aVMenvj+HQUh2IRzYBU1ZbJ1WbcSiX9Epryhzqw6NIRJCo4YY58MIj9hSyeYLxpw
kkOK6Ygf2xmvYLqWv5GiMm1YhMGwIR0s8489Dv9ldG/fuSckwYKxAZ8c4qHTrcLE
q9DxMA4NfmRh1i/cbqS9HFJ6lI2uhDazbB+REogSlcAgpbC+9mcJojBhI3L8Wowa
MNT7yWRUxGPHeZ+zY2Gqpr1C21kZna/t/3su8uu4GYoWJZ+z1b9GSVwdv3gLgbWe
Gw6qwJKyX5dMN8RAPtU18qvwONUDWLGlJT0/fMKAY158BUr95wezrOlUReBLBnOj
7RGla0dr93s3qlfngkDksjGtPN7CEBsGeEkq9oGHGhAKOp4A/wYKqL/ITQ0oL3jY
zMDni6rfCdza9A0Y2Fea3JUpak9CLztGdvtlClXOgujDYR+6khjfXUVcSv2OyKdK
18nTZupOqQHqMu9+wailYw2FbG4rlaus1FFry1vtSLEAnWqHLPx4fNLw6siACwwi
NdZilvhA6TCqy8Uk5S2I8vsZEwIqX8fl5AJ/xlXxmqUn2YjcQzs4H1KvycF2n/NL
Wh9zVFCVgEMQSF3FYONUSathYre7vQhWlw22832fdDdSnh1Ntau5z+4t3T4BgX9w
TCl5QVXfh6y2PH78X78AIk03uDs7AfjK3LZgPQPCC++FPCHYmcDhoPxNe+eikt10
CG+aBqk4UJnJnwZY5ry6T9q7tjdFGOwCkSdJD40a2+P96PqVcSEm1eLx5kIdoFmD
4Y6yFI3Q6/wOrbG9i3hxdUEsRtCi6N8USQbktIJWhKvqZsJ6BicANPgpRa6YrBP4
A0f33x3tBvnAYmyxZVxXO4bCI630VjEnLdHEob9avb4XaCK/BGVUV2anNmqnyVI0
r4C4Vh6zV//cwthWPHlDR8lj5XbEJrzHTAKTu6TRHdQmdHjFP4TPLIDLeD0bJYD/
3t2z0u/cB1LogTBvXeucHEjbTNJe69khLxOwfJ8n36rddIdmyPixQn2xr0BrVNJJ
u9nNRU2xYjckMREla2iaIz0ekJCZWef3aOurL9cgCWA3VE7ZyYEMx8uUbBzKuSLb
metxLsle4pIvQzNWkWWMyrdtjiVpgC/UehvYV1iJ4qTnJwZNEwI0ZPV1bKqbru6A
xA30gi9c0vmvkKb+yWR73pcomTblmG9YjaPpwPLwjsNksm6zOII6PDfjI9RyKJ98
1x7VmxR/Iw2x/rwUSU3WRdtBDR3Adhprq6p5A7dHxsRwPsK7oI7Xpm33fRcw6Ji5
RntMRJPrIWfdC27gi7T9HJEzuy+C8r54OT9NeScPtVGezEACeo6XiGeKnHTk6hWj
tBUYZQLSwKsTHscMjeE1hqTHOa11AMrLaDbqC+cw08BSzIYvnTLG7pxotn7GWDxr
RfLZtXDgcc87jXsmgfWp+bvygOQTybW0HHrpImXka5ErM7jF/bxsZP9SY4LgsAGX
OmKNkZ3CQ2cEoWm7nD7rroB8aWz798h40OLmJQNeEZBqaaC7qxf04/kfTx+Cbk7H
k71FtDSG0441SCQjIPc0KQHWkWzjvVCkJgXcwpiBg6TIHawf9FaJnsGGudV83js6
dKt04waPIRDbWL70IdTbBVz+kf14DzHf7tPh3vhWpNoitLREJzINUB4lSaHPD8ws
pJ0kJCpxSfNs1OF9Zp3hbExx1d4Gu2yBEF6VLyJ1u/OuBJqBeSBr2OOqGKbhlLHO
xoEek+qybDz2GHGjt5mntblmIgG04LsLnTLYsaS9Pu4+VuRPieVh02eLZ1Lkv7qk
iGPURyBy6fWWxD2k9xrlJhITrWk5s/Atbq9YdKCUWGNbWygXp/xZ9pEne28EVDm2
rsBNomsbEScR/Y0WvPsJwSvQ+BRE/n8i6LhYW6iQ9jbW+cwaBXzrImU4BDCLPQ/f
GfeLZNXMSFPcAWcfY+2YIOqiVYMo5qeCdcw4BhQKWe1TQabtl/YRsOsXizXSpNSd
IjSyTqDe1Ey3ZmY8k+tz+McJF9OvIHNzVScI1maBUZhhLMxF64oH0YXZi/v8IzQu
X4v9nafz8lW7vZN6X5Sk/tb8i0qqerVH7jcdYgRZNgdta43mmppadTjR6zMTxFqi
WJpaFFOsIQW2rnZ5/OhHxo7j5z4xFz1Dt7MAOnOZjHjfLadJYea+qFc801XGwt1n
WvOho0tIY9ErUvCYEGwnkTK4T/VATHFdV0EtDWQGaKkxn2x4pVnF9Q3NKfNbKBRT
h29WOkdWPNSRUUUfXP7QUNvVIHSQApQODjBVbp6l7JsCfa9Kc5uFIUeomDaX2hAZ
vHUy4eDf/+sGmcJe2HHh62tjzqcxHHW4oTtovstEmCMrOr+Ij1TCY0RcRXy3RKsP
ZMLIzlNIZWZGcfauq8RBWRT61YoSvNulCO/pPwPHdUOcHhiBNd1En02zLUME8E1W
9hMqYNkDET4pTEtlRLzr4Ow6tRwZbBXFbDuiWIyVuK6YSLCxI8xf4Xcuk5jw5hJY
NLXfijpZGlteKY+kLK4WGdsMxqz5Pq0Mgz3Zjr8IQGrjhljoVPy1XP04QyA3jACt
ltNpi9T/w9U7aqZ80Lr/Je9TXy6se/vxbqr3YjNFTGgQXq6JVCH6glLyTbtzkNuH
Sc9lXSV9bNv0zk5mTvZaW4NkKZ2Arp/0EodUWMRvipBtdkmdMPdcAOcSr0VbkZuJ
9I54IAXQ9p2p2ndTkIuWNTrvg0itpjCh904HzClkdngRu59aiRzL9I7Bz9zwQX20
hxsJ380B1nQJVdI8hvZRPT7IUPmpNbOgvsmxFelitRzH/hT4aZQ6F3b/KMJgEGcL
pek1/HOs+osJ3sQAznha0ZROWU+vQPEfSDi/6ewWQy281NqKfGBseelyEIh7lfVB
55GtORjtzICQGif4jlYV2v7bW7mfYd4a8mU1VRVHAcJ5WPCCDKqjRWRH1Jky0+QL
s0205HnfqLRx6tn8sxFnb6s2x/gYAkB8ObuEHZMIACKWBxR3TxU+h/B1VDAqLl7i
ObDQQHGgS19fKJOoaB0nAEBcs6SIFyHlFj4T63sR7IOi11k1K+8DklR5qhsrcyUQ
5XubBgoahNtsHIWao76eTxqNo3jvrcbFLze/ACffJzlbBZJ/tcIjNfAQjRbmswTG
48ncXGjtWttLTIkPRv07pn57g8/oFsaWWND+1KSQAasoUd8Y6Eqk/at0OFzIwK7k
TaRDI/mj55z+yuNEMcomMoXCrSdIvKjdzq65mggOPRlzDUnt+D/YyAPvey61f79s
mA1PgvA0lzLhR0gtKVQc+nmgYPpbqBaCjDJIW4LYIBggmUBE7oCIuaATTXeKSm1d
IqM9LZ3LV7nKLKlWhjyi/sEWl/YkZGD6kDYM9XS11ZvcAkQTGSHwIYlHy/NmyO/V
wV16zwoEHSQqNsUn+JsCA1T6KGbn15RBG9MXzz2X7yj8DkvytcsWR+kwEOLqte9c
ZKgWfvGPYKSQ+aJl8wbwRFV5BQrbHfV8hWIyVJFaRploXK08x9XxdR+MSEaTh51o
YoTJ0gHHgTYklDu9KNnqgCdLEojqoAgc2A/zgXJwyqbEzAu6pfOLNyg1+512lcOu
uJwRodfBxLckkmcDPWjOGNDfOxhVh51MgT9NmnwTYBt0jzGVzhae+n5x8kYtQVX8
IJGK1F0SJp2NdfUYebD1KjTQ+1DY9EpOYtyewukrOa2XTkr+T9ImOvRpZcFf9RyV
tXCEsGfwZg4/xIyTAqLjmNnOju2JZOHsKFBGxbqqt0+wj3+abiaz/Eli/iMapZ8r
c5pfx4LEstDwmfCLdDXMj/VNNKUrskLB6de1OfFCfMdWpnUR3fWYZN1X6akG4b+6
OrsNp1wopWAGWWWl/M6opSjsiFCMnA/MwhAirvJ5t2GpxXvqxSw3ZluCt4+CNH97
U1QfG5Yo4xXBH0P1KZPPbwaWiIcjRpGWHZsS9sGBk0iSVUBfsifKKFfY6URAslh2
2vV0W8tyw7wzc04CbHXxHwh+yAwL7XZGVyPI5d7uzRwfPO1LOemHKsNvwQG3enpU
Qxzr74k6WhmUI3PkRXttmI1EsypDhRgYNZ+2itrPN0EU2NcJndyntPbZrhnRJNzm
Z41izJwbUqM5dAbJXyuQ1Q9ZguwezxbtjX7dl3592vOFx8bofe00GAqcERdaTum3
FRfe2LdAWCUeKZgkYjqX8hEWKp6fN7Tycsth0WpEwiJ2YLP+yKRGq2j5lGZAfJ0Z
SoufSDULVX8xJqWNHOrgqCDHTVnR8yAvX06l0piQC/yMEEQBoIJHNE1GjrfFRZ7y
EIkxf+cxKzlowi5Pi8mH/DWhI6nLQ8AtNtNxDyMxj9Q5QBanoXD8HGPbwVpKGr3F
PIRKGck1Nk0XFhl0SDAhD1tn77f514p2Tdx1bkmw7E50t+luzGtrxnZ/AiCR5tDH
+8m62Lofz56Zmzq3Ld2SqlPEYu0f/HljnXrNn1vMJtxCJk706h4bt9SN5YO3rNdS
HLJQdo/9flMxTkjmkGmE2w+/jGWXXWCfCsTUiIlQF3Ir1hatjD466Nve8Tlym7x2
UPQ9E0ghn35SsqZmKIJ37WXb1Vw5xtWyJYq9Uobt/YfA/PcU0vu1JVgvX/rZmywv
JXZ4ewt+qngcy4u9MlP06P6j60V3EVc6i6fC44n44FXGeaXASRTPCSkakkC0MiKl
UQgWNOY34qSOHnKpQnseCldJ8rRHvvOm+3M63bWO4ki2xUA1eNFKOR01xuF4r0f7
MG811wP6vE2o1RtmaMsaqXu3IgSUd5G+OdIhEMC/c//kSaiiXER3HXFrnTJmpLae
s3HwPDRfbAqpdJF/B5oaxLBsmkkhb7Dbi3VExkDBk2WSr5B2axSZ6JmAQY1bjPll
Zf83AwrnFngzNUOWJWrTzQkGkHAfHMG7NC11ap2UxtQOrtzjZZ+hWZnYiDidFZoJ
wkb/j1R0jnQ+2XqCy8WNNzbT5R4/jqijdsWkd8hp0wohmLHtZXvyovU1W5ZmRH8v
jEGy+/F+DNHKoJlaS+GIuVfbsC6GS5ziWiYrulNm4Y/ZW3MxWLm2sDOYB6LF1JoU
ey4MLji6+GFzHqz4Dk7fkZMeHQwa8AhUtdDekIS3zhgyJ3+VfsEvDKjoC4qi6f59
eGbiPmrwDFj6EwlZlHqoNEAAtA/vcF9AObxyV6uzqIsFx4hiNJRfZEgUi0wpqWTy
7sSwRqI5mLp2TbKUkndie+uVphYPlQGWsuy4ZxiZUYzs3pLh7E2bQ44FWpbn5AS3
LepODTbtTtrNEuI6jXcRq8y+g0bG7e6la1/rPmRjjJf1O/zo3zQk8FCPfkiODV/d
a0dWeTNqFR53etb3WnXlJ5S+ujZWXbgWIBenNleIBRWNk9ggkygTQOo+uQ/56rPb
MHwpdXKNnIV1n5A5N0AAohA9oC7N/CvNIPRSJ5YUFti3pI+livpYuQ43Gv7J0Cz8
kMBmTOQfppe3IdLQX3C69n1mODR0zKxKLwmwcWm62McMtfbt1iQjQGaU9433ZLOK
8Kn+ie7Vz4w8M/hWdk3pvsdifGUjjDJNcsT+7QsuY9MHh9kg9t9qS2PYHMpZ20zY
bLzfiG9dUCbE7UAChtvQfHZ3iz0QqXXNmWgeoeWLt7nbfBg0Wa9HncOTxsBgR/P3
I93rhRFUaadmDad4KJaDel1p3nQDfOrFJizbPAhw0tWj6G2PKphjD0IZgnTXLTb4
CumHtekBV90z/PA6XZxSiOwLGmpd/mi/7C1wAblW4bqRlHbV6/2vmykVc+1EXksy
NQaBo+PycNzBigTXdi73TKOaFIMIQG1GuKYUGFRjLZpTxN3siXd/SKqrOkbIcIKp
ffZ0EqOXDUy0ajtsTRZkBQMf8KjwvCFWrpW+ePIsQbIbuJ+UEuw37eDNeC5OMbM/
ckAStwQ4pyH7LXfrqVrBk8ltz7SlqarD1ZzljTVFd4SsjZ0SlOVcnjBd5wHrq2bW
isMb5UMv6lMvxLt1PnLmpxpxhkuV6GkytqDn+uSyWBONGXCIjr3+PAnluQtZEGCj
1F+Nbd1pxVXMg4uta6EHgvrADETtA2NtSPRpwkvl05Sm5cvESWEc1Jo/LtC7ELCd
lTQCkmsUZDLVhy2/xNllbPlKUcL/C+GO2NVXxt0OeQP2RSqpc/0x0JoREHNLRKBk
Ippd1D4eIlDE4mubXP+KXWPulUXxSE25GrC41SkajSo1stYM8hLjhntz7vQ1JOLo
zeyBlMl76auZ+AXs0y252rcYS8QRDIPCBm9V4wluq2T6hAiARPdYTP2j9kKQvFZy
7XmIIrw3dL93EQ23dBINZJ3uQLtiV6N0zOZ5JIm/10I0gOQ9qqnKRkgCoBIDdwBl
Kgvh14aX31mtcdmlDE18Bgcy6JRD8yucSS4eZ8jt9UU3wuHshlV4uA5rvu2CvTs5
Ly69xfyYwEA+BvZ/7LrTwNrEyrJQLUmdzcg6OyFDkJHtvkPuNM9XHq0jNu9GCK4N
L1tXS+cCSKmkomkMlo00vTeghmp2jj6iZijS5A6LSlnXvu77zXN5gNZVlm3hvOnI
vK+H3m2qzJGU5PaAHdM8184CA8za3KwBfVbsjbtCpQMbr5rE6RL9QhwIg6elU8UP
IkQ2fiyrIW9fevgjC6QiAUJrqhS9DCucuK5hIAA8NPlUDF+PBJVClZN0nE7+GbMI
fEWe2vP/7Ck/P4v6Zh7E3MP3FGJPLvBTNoN5ZPXN7NgtUOtnwNFNt68PEOZ6M6hj
P/1T6pCgeorPSkMWatPBWvwMWvscdEYCR+N7BNKs1Nos6okzkdCyyWYWZg1scy74
4g8ktFWvqJ5pmkfAVXRY9QPUPQWhHvxcuynR8ZKYJ7hmLDVdON1NnEUp9VGFyjdz
4cBBOLX7DrmKyIYEZwPTJfsrePzQq8c9b/nL3K52RPMYAnolAlqnBqgsZYcD9hT/
LNniMdptUWQbdYnvRPpL60nJto0QSbJgrg1zX7dlcr5Cx8XKwtNC9lDVfDUJUYAj
2Qm+9queSDP25OLyHNTd6FTRYmCoTVXYz3K/UO1xUlySn5xfLgY+mh5TNELfvXRJ
h6ETlsXcOqpptm3wACMTPKthxgCYzyO/ptgLMD94lUIgOa7Gk71Bh45wIk940uGq
4ZXZRlWn9moIh4ICBhLrE8IfIgTNEIXrJKrUEbibire5KTF/+pn5xlIqfpoTrevE
7WvVVetDnLLR9KCoGd7teyFYhOM8shIAtStjPpjsT1Jd1hBA/5M4u+qzZqekX73c
8i3xZE/DL+pNSkGSU5ZfYii4Cd2ARFTsM+gL5EC1KAES8UMWCYZa3JGTSl3QWVgT
H5a95TfufU/MGudSCn5cip2Gr1AixknGdLYOGV5uqdB+MfIX5MHeS0Vx8hxb98RT
Aepq6AHfqACHBqKnoYXkNmuuMDrM5bYBz4ZQ2uOd6TjDFUfFMN0kInN8ebjy0wLn
L9deHRwVsgaOJTuPYfhqlF9DURJ1Cp7vQqI6LOXKbDAmRbgPUHCOSHMotLXF4ktW
6XoZEaM8L+JYObo0AourZn4MpzdRrO43Ed8ytB8goBlBx5ZuUWp5RXwPprc5y80v
UyXuaSHHXIMFf7N1pSLi9XdK6e/UGmuiAKAEyvKOCWN9nTwW8u9tgSqHwa9M8+rf
Gem8liIvlbKUzkJ6P4/M5EEE47UErZECr7psAm0pyUCSrxHygQA9qFkIis1ggBu3
Jp+4lTPcq/sVms8oZ6FUzYgMFlG+TCgtBFolafSnYGAfEfcJloXbbgsFY+tkDOow
TnFIADaHksqg2Un/G7D9znIuY12ywCLBr+pZ+DF4bbzjufX/xDXjT+0+djX4NQBM
F+KCTK+ETVI9+SkXWvJu5H0bZj05aj17FQtdTv6XmorA3oRh7HP+LOXIVTAKoK9O
M8AlK2tIkRsDWTcglrAvBro4JrS/fu0zfX+i2a/u5toi7yOrbn6bbzBXSOGXhEn/
2vhnaRe/boEOWGBaz9/f+QOrsG6/+CrJIc/91pjm2eNKbgNnCfrzQ1bIgWcsP5Lj
432wH0A70mSxO/ObQ9oN4tx5hcKbdkknA3JmvFanMPUXz6nHw0WvD275aDaPsnkb
CcjD3IL+fg/S7uB51gUbv7AjXNgpB0RCLTOTT25HIoFOTSaPSbGvZP+fQ2E4nFCk
qXnUae8T6OHdD8lKHev8LrrsMNbEu0fEdz0YwQIdl21orcT6af27chi4hx0Vntox
igl99AYD816iiug+K58O9E7+s/1iALS0dYCsiuLU+eYfdpvX52ocQ8AvTi6kvb4m
LcWGOaO9v6/RjzqlBCm+UUanAnAAPt6nKRvQ61uZFdV2pZosKCoVFOe395+kQGx4
KWyDUBkXKlyzVt2ThkQSqQdL7BTvQ8oO2bTmnDayek/XQYHAt33gF+uBsWSW39J2
eFCAQNmbi89rOMF9IV4OX27QBZNDQdoBZb1PgZJxsG/pubNl0p9cNJo+UhTC1kYX
EY2F5D7amYaV0ukFXHvl3pqbJ7HXFaKJdv2p07NnW4BJFENBcLmI1k/2HnzY9PSF
SSr27xRN+xrphF+SakQkc0ZTfgERuM1Xe3gwLjt3i0+0SAvmr124DZi8fLZz1Fq+
nYYTzcDGuH5rK9dmotpXt/jP5ki0ZC6gxetWhQL3dvr2lueS0FcwDfHoItBwpa9M
MhyGsyV4Gbd8cSwDo0sJ4Hr0d6VUDF3tjRTT7vecV7nfqd3e0GlTYny18ZkRESEp
T5BFbqjR5utMM4a70kNqArvyx/9tDYxXNlSOkDlhIYROHZdwkePiAf26Ua13cy89
6WWyXUAAEE2Jya97HGoK43N3k1e1/KJxMomfnFLn5P86Q+y6cUJwepUQ2W2eBBZe
qlJ0/pQUfN6p+OYpxiY8PjKtDVexvVSlZCOzJKKY3HNPvYmwxhNMuMHHHTDLFF41
CqmRseB2LQ5cBX4hli2nh0AQM+w+VigweNDj27f62zu0tvvcAW81WmchMTNt0yX5
+wFvBWESLpgP05G9yWHaFsRIV6Igd5Ch/78yoAQ+io+A7Y3nhw8dKrgIduxY/F6S
bS2NMYskMYeknQ+BlR/3aSi50rifXdTU8jW7zHIa1BsZITnbc94N3GY4k87KVUNN
ccmJDeb1IV45CDP33IwHcvHoss5zE7awsINcQQEk8OtXUqMz5krIRakN2DPslims
wHJjRxWzrXqxaelI/dOFYorQucSqk5TBBhZNSjZiWkwaxz2iC6fucsSgZr6htRMB
yOGm1uxZ4Bsler1RWWqkDBR0CCuMGyS8UQw8flOea2g6lOkzpTpZ3IY3c8mE+XIX
KDqcupNSPyjJwj2KGHrP74aZIQUpmNfQBh5YQX0M6qWTjMWGRSdtJvfSoMOBy6rk
oj4/IOS2oczTYMQy20OehXwA4xLVSUMYHZ3iolmGamoRwVpTpuSxywSVqqrOqBQD
1BxsNw+eMwR6qYfLyDKC2oxa3Hc67fqSXFbUUU4i2qj6Cl6z/6rRGXml1z2I/2fD
29OHgsTwO4NrjbMXfe3YzvyrgO/d25LvZoTqcFJD2IX2PuXtPj+IeCMJC2G4wCyJ
/aZLvYjqB2qpj82CDdQEvxHOkPwpMjPI2E6rvB/qtgb4zsEtacUpSiFDumYv7hJh
nVUMB+NbDInfXMAnlNOvlnMJuJ3pUXj6mIAUvhU9cEUP8mhoCBXP0xLnldIAmRin
kASiL6D52GJ6L3Kmybx15dVpf3hauG5GwMhgyx0N3A7F9Uy6OhC3omktf3029/fZ
opGSPfo9kWgELFDYn9TEs4mMnDyoA3yCEjx5xI17s/G5aLnJ+7evYLCmJgikxrGf
RE1mtt5tP7SI0YFfqMMloIt77DAmUNoubhkFq8QclLughsEznCQCKXn8QiCau1O7
0DW5NujlyRKeYvUxIUjMLzCzSYA3IGHvuXsrXzENlIP8mtXvINX30viMUeMf1UuV
Zl8+XweVip9r3k6JFV9grqV26UcJL6FCwTLAuBbv1VcEqvVgGxuHW9QeUxe6FN5n
jdabUCtkTfoVxGcNZy1MXqC+POhbbOf0VeGA3GxYc4hZ0uu+hbDaTMVz8dguE508
73zd7gjVErMpe2K/TCxyMgB9pDL7BbTJA5Bqzad+lhsB/jF33VZt/wxpvMXfPFph
/sSWzoF+g+W95dY7u22/Zfmx+6OUQpfVh/mxwx/2BvjsKnpI/HmNlMVUcFsDzoMm
V4z+2p+zzT7nJHmBVrAKoxqkaEayhkTL3vNZS5NT/5slqou6OjkFnZ7SEu19vsFo
/IOWcgemCKTokBJC1YXJSwqpBsNZfDW1YSrkqITNM3/Td8ttHSzhmhKRwEuSYE6s
fg32DYniXrxtd+fcJV51wUIzgUAwQdZiIVnD94BRxcpb98smPp1AeCwkaBMRzMA8
sQ2BNeP+qi5A+sXwi7GLNjV0JLPKNr/6cUGxopwCaTvpiy3zzYsWQYNLSB5rU+BO
6Ujnnp6nDMIZhA4oEp5tX9b1eLwBXI10XJK0Mpelen/eO+/q4ZsP3bYt8/f6GudI
ue1sFh6QyK5s5kF88zWn6/bVAJ/osZfrPv3tudUkKAdPX8UpL0QspJjWIg+1ryFu
IGQ8bBlmtTP3KOY7ivPTfGR5loCXj8xdle0KX6sbMjYGx0QTdNUO8d0ZmzB4E+zz
5z5aQ/Sp39FHM4S4PmxWIfuChKvoTt+kP55asa4bSdXnzHNoM/VfwLkloEMqnjG6
M5sxb0Kp4jU5FttFEvc1T7OaSvQEXwErBUIRlDfU/L1kDr48+NNv1WifyU/YLJKa
Yg6gY4eBmc0h1f0KqtBx2g0SYc3/DFRRP+o0PUAEgDZunfyRv4lSvkCcDuGhZCvC
xa3vQSmYmrh6R6mw/IDAy50LNEQSa8i7f3X1VrWelvo5rn37ZTZ4pvmcfksK9X7w
ZaRwC8ulzM5Ui9hdcdPH8IHzwrWiDZxarfuIpRCv5dKM0VPEU1emuWKyboHtc7bR
9fJvi1NfvQ+W/InnlrNdW+b1wA3/6w0otGVzh1kcbgC9MWDqu5Odg5dzyKLtIKUb
HEOrjQReJ+uA/RMpQ9bSg/rhRmjV/yX6JDzRMFgXt1Z0rs7HaYPLCOzNeLr1ttPV
WaZktr4oron109AeKD4qXcI652MCCcgODu8j28gn0igungT1bUnfuUPST7XQHDVJ
dJ7QQ9CG7um+q1DQbkZGkvEQGfvyR+NOVb4/qACvCnSjOkQpD7b5qgDDd6BZE8d3
KxxRS2dWN4XN5eeqgSH22KfGK8I7x5JM+p1gtCaKe2LqphqXysl7JitTum8fUApF
vRQ5d+0HVUiuEzDmvtZwO4/0OIk93ZOYCu0UNF+LrkrtS4+AzaOilQhxWRfd4zLn
C3W4pKXwsTpH/6Ftv+DRVmuJROH7H2LfLWWbJ+f/mO2JrVEUtxFPLOyO65xpjLiz
9vB9yb0J+uecqCDjIV1JFkvh4nVATPaPRFkUFm2kJ/YR/j09/Vwx7tw2Cr4SL4zS
AbeXv4FqygCxS9h3Z2OKAV8H5NsMvlUcCRaQIQyNx6xExhW6NfrgGM0o8sfdVz47
3uyhzu0UcEsUY5qkABXk3Bdl5a/2wxA/blyaQaOG7i1wrDmjBR5LQioEpWonaoNa
SFtOLpdT3fkAc550ET9XdYikhtJJ48To1mu8BXRB7McCzDUqtaU0PI4quh5UHlw5
sXcaggBAlNba/xQALoh4ODEIDDElq5mRkcMOmTJ+UrlLxkcx9PIkzb2d3CDiDft8
CEurUIWpkLJ8Cpiiap1Dl9jkkok/eMA0V8HCtn4EUrRDGsKNIYCoPyqgGyrJUks7
RSCF9NrJDu3jXzyTRO/SmB49K7rjs+Wr2snFyPSqfWNxSGZCjkbIVnfuqL7OrVaA
HiXp25Vdvdx7eAwmt764uIsLbP4SC4NnJAt2Yxsk1G9j+KpU86leTYImr8ylw5wW
3CTe03YQD7xRmYwP/YmEmkpT5jXBd0PV5THB7yqgWuZ1sAyD0xN7pbZ+vuzgUPbt
tMoEW1uh7dQFyrOKepXoQrzqNPkrYUiSiQIyoKBvzfG21bcVG/sMWs1cQC22DSxB
fxbEGmEn92ObV6tKy6nU2iIM4xp8ah/+X2cZornWF2um9I/F/IM6spkI2pA9WLYY
PbckKejOiUMHUq8cHLa31cIj7MW9Qa9zjcc5UdoUL8rPzU/M6pM7TJwd70n3SCNo
GbDlaSAddPAi9BicQCPr0euAxP4OvD03Jp86IhrnJObB8vUWaH0W77iOIAhKcWYW
ssnw3wWeqkb5o0EQoxJl4Q7lZIddMl9LBBEd5XFi7LxE4NJm+5eBW5ndahvBvb4+
DmixTjYmFDuuGZPkpqlDDjyRNCIDOdaTNMDOdx9eFo0Pu6bpduhcOgxuFF1r0Sg2
OaGN5ZZ6PRSv9Q8hdlzttTaLYZlQUbMf+7jJ0vdDig3fAqqbdsiBgBBuJrz8Pxkb
WOBpKJoiNJSWL7hsJ2Vue4N4a1XeOP7sNeCjlau8hs5Ena2urbHDIhcPhYDA6MVq
vghVEpX7dvIfZAMsC6mm41ayOtZ1gGKiQevf3rrIdrIBiBDkfaXn2RxOwmccsX2b
tyE4I5UwmoewAgmPliD9Re1b5/JNI80+Lh2RCY16JpvTr5EKPpkY34IGV+LeLZ3e
f4DRV+08ls68uW+7jeeBSVSfBbIVMWV2VWsVcR4L9zA3KBwJ1F4IQwjUl0rFG970
8QASdhw2JZX7rgXDHIAp4tXlJLudcqpqHQyzjjmOxU69ExIurNtOfkaF/KAwowTx
X8aScWpVoMBSQEoawu/PfHjDjJx2cxephfJyB30iSVl7Icaoj4W5AcIblJSVsgBn
KEDqXko7zNweJfn7uwrzlv8DPC9URnFhL2ya43lfy/BM+qGrccdORvMmbZiwMQc7
lO69qXhiO0iaqwO4scIcPNPUaas6sQpErZHO9B4sgrjuFDSTnS9/ldfEZhXSpD31
Xxy+Y7GoavZYoLrzUhOBPy2fD4Gsi5nW896VzKzAGBJBYkToZ2n3KOI54MUCP0ah
Faz5i+nSAJ5GTraRo9jNLwNW86sgHy1AnQON556ooH+WQNZ0H1LhKxZ5H+tWgC3P
NpzTAPsKeE58/6gGVdv2SUYk+WyK0VTfqXQrcQjnUCV8kg7jEUt4hj70yRoxpIoC
PVsSDtCvRk+kzX8qVSh/3NLlEs4oNwsKZURZn6+6XwGBdNpC5gc0WQd9/jgtak1h
Z3ufJPjKjCSQQ7izt7b/v8ZpljL1E3NJRX1SFxzzeHEW8ln1EIr0RT8uE7Ly1MSq
t27MMwRgzGi9qMXWUHNvppj8PRCTh2EdzJuhoV+Y5pvTfM+DVptrW0JMLSmVNCot
LwZg38W+H0id6PoZVnpi4hDSgmApacpLu0KdpdmSjmgyq6kGjFs9a9dLErn8mFdN
bZGUa71v50mb4imySY6y649MEZL5cb9YAhafT2vaXfu0gAh61hvuUD58kNs+M/kB
E2s3OhXZyY+kutjbWn+91A9eLdW3mXJ5GCyHyu/BfLjq/1HBpib17d3Z8Tw8ibYV
AlV2YXZj6J08UOibcuOs1BBSkT8srY8NNWn3hSxVNXHKauD7Uib5L5Z+c21nUHGB
tCPa8nu1FaoO9OzsChL8i8e8uc6pvN9N9QOOz/WHpjd7524FTihjHv6IUsuAYa5D
AV8Hze+rB4zlnnpq9P1nktrkah7x7T4/gT7/MlkLEcdtY63ysTVIWXpCuyPiXZ3r
BSUcgDnUEDzRrQTBmXDRE9nCTdYK5+OzC3NV1toUYtfg900J4IGjGJZbvKjjP/kY
S9/oqZBJP8AoG1hBYQWrOdAREK4I+olseL6ZBPyLnmP7QWpkohsS4r4Pvh7QGAwY
WtVNtaavVFgOBwy+TQfYVn4GNdSZe3OHczSRUtzEvzPPGpB9IxoSHjS9CKf72yiZ
+FhSBU+bUsW2ku8W4a/oT0Qd9t5kKFHkJv42GaRd5BSguj7KbkZyq7aght2YDZjY
mSk7JlFZmgPHhR8ttra2l7Nr9Bhl5VlVTZI4xVCTB94s7NUoTY8nszzQPXZoaIxT
9YTkMzYnH5SN10xsTLX+uxyZorfZnlrwL4EPpIQGYcC/ptDdQSFGdGuvWzTqqGWF
5zxAmfdCMydwhhL9PAYYc/dkxA9Zfncp+aM37QUIkU6+73WVws6PbBaea7x5fNhv
mB6te5Mou2pJWgGBAv+aGnYoHUPWLJ/cC7fp56FqIXRUVJEZpW8316AZ9P+OmFeT
FW2aeeD9w96/P0TdyzljaduEJClEmwdNwYV26r1G5cN1oWc+PIG9MH5I8Ct0jODv
VKkd8fqYdqlBdowINKfYupZObYo575HWSfRmsFKFx16J1oINe+jQjv1+8GYjHdZ2
dHwhWcnq9TlFt8eC7ZdTJM6AafSotEdqQBgF3qbC5xyUmThd3Qa/oe0eJAIwwi7C
HrJbUnU/hjEJ0ErSSZgapRPWsuEMYmJdMSq9VO53CXRBWWKWEmjOZpqCXM90Yxuy
TDz7I11puTvbBrR0o/76180BtlX2yXjGdriYBKG4XCIjWJC3FRz77rN+dinCJmmP
3wk2jR8q++t3wzb8lYY9nNFRyOlZR/vb++/akeo56XYV4QjWoXasgChVMuT58GiF
XbL835uj+w0PHR/RRmHpt6ggXjLk53Q2nrEEc8PA7374tU9hgrex2wuskOz1ufd5
+Qm6w8CC/vERFv0tD3VPlSgQ8ycMZMrVkIKhzC4fP8D484gBZHHBplBLpn27v43i
PvRv+NuMFtc2o+LAlKTWmT9RXiX1I4qeN5vLsapoJBQRJSaUHyZ97xJiRZNgyEnu
STIkCLHdpev1KP1tU9854Qy+V/3j80w5EedSh427aihhbpxovnGR6hROhYs9ZgMK
OZ+z79jPBpehmINkhgCSzNQuJjBVRkU7UsjIOoHGROql8YjUI8o1lGFv4pdJV4wM
loeFZ0dfbl39UjDai3ZjHuqxkLPXarV+nOIVHD39SMQuhJlXiJ29guo5oKFMEn1Q
Ua/HoXMr5Yup57ru8LzLdMOmZA6E4EJbOjtTDZjVbYRtBvN78CMrv5C8IQzyxLSZ
E4Iw5+il9NCxBP3tdYZAs42Ut9BdS9w/Imlj+wjwZP94O0q4ZvRLlSye34Ay/eax
2LctxMyazmfAZek2VeuCLS6Sey/Bhm+FVlWtM+2BXxkuc1ZplPsBD2wPrIk6oqnO
uZS5gHa0rY8ayLXdFeFbWgz59CDUKmohcpBpRa7GuUySflHYUCECUTQM1whmrU4Z
M4BhqENIhBbSV+q4gvpaoBEYlP6dFJo0+sUctZWm4JE6G5UcrOAmTik2S2dGLohE
/iSbfP0quIATMggn7Rz0dS4/K2XF87ftMU2QLawmccAK6/muLnQtRJvQF+qpKd8A
3nLAcuoNO/FRQJmOzzr4IXhAkl2ex1iAMnWD9pyAm88NnjDiIbHuYbK8pO0xpF1A
fjfsPeUMTxLRnta0cWf0W6r+uUYxsVVlYz7/lpQwnzZBAwT4qmNM/QpgMtwZRR62
UU0t3p+Sjhas4HZ5/PMPjfJ+4XHoTk14VrNlx3uktapO1ueiUdRqZskIfjS7BS0J
pXNryGKzKEhpj/73OhAG30VCSXJsDLRU2vtHfd/hdBTm78rtmxkt3vuviJCKRnwr
d9u2S7fuzwqRh27gnaobv27acZINQTdYkPpLmqR2JlqeJLEJRV95+NguJ/D24GgB
RoRDnFqWTbqXzfJzrz5BS0KtrI6idqM/XlA3m/8i4QNCUph+nmRpAvX9SfT2RpuL
YZIC5sZIkq7KzjTi/2Vk3Wd2VqmyP8+n2n+WAHxemoUYDgTchmh0ETbv7hTQVqWA
69TceeeglHbguxwA2rEB31dh+R02cLcKw3yXVGH5XoRpjfyAqS4bHLcZL2tF3j+O
eldWyU3YuBh/B7TH/cjqdd/XSel9hCQmM1h4T14r1pYUaMdExsRZnTep0Z4296dv
FP/pxTwHGI05YE+g3y0ylJGTi+06LnM3JwXRnLmRxi4/JMnL0fmiIzy8lkxC4wTH
tcvQ0fNYKaH5atVPvpJL9+CjiNuNleDe4iOAXEGHxLHn6aIycQQyNyuIYG874b0c
HlymIX1u2ZPGmn18hXNzdsLNOvym7Tq1yJPlL2ZW+F7MZ7BuUUY7Grf8Uink+0WB
Pawe/xSHfiYk7Xq2mr4oz+kHD+TOf4AqsikVLHjEz2D1/dlfLdX9LIkz6GcZS8IG
ebEU1DsKHaC90+2+d0mL9SDNgM1L+/Jb06LLO8uoBqoD4Nc7GUW47sSzwvdjvmgR
3BywKIb3WWvcSasvhO2kJiIqEdvwNSCLjjlfREdyoUMhNo4mcweH1LsLl/ifzY4J
+x6Edyx5RpoBUG7MUyQWKLnLzkVOVOjUhViag1qBxoe1Oa0+LfdpoFam8Ce/nxcE
T+Btb6+XjCgzUVehYek9JeH6/nJ+6AC66s14/1sx7BtNHx7RQtbPc255AIk9bpHL
FapggnInL9g0Mvlln1YTe3zdhm7PUyqWfpJIZo5MtHikm2XJ7NePw44pAzxGP9Qq
a3EP/QoOLU2QaLXQJFw8L9y9lQ51XrAqcL+oodOiadq4tzln6sfeykdfhRNJ5XE2
60omfe7NMTew05ETzewqhCCHFhS12ts/tgOxkibfKLTodugHq2oA7g4TOU13k0ps
YM7UWy4eg8WvGiCdLnIltWcNJMIj3cKbx4f5ztbPzF88fdj817Lnc1+s2iY7FkZZ
kgmuFzdvyCcoYLTJQqSMxdCo5nBIviq5g0mQ6L4Cge1IKxQKa7CWMBMCHK5o1Jkx
Tp4P4BQJ7iT9KFDpO0VyDSKAgo77BzpHCBTA0q2aZ0kb7tDtWOZbwORWKdA6t4qR
nHe4Y6U+Samif6X/g1mDvfL0rN2RyiTrBkKyABglOGyfwrgucLGte/+ofh/t59eP
FGY+5+X/CoAeze4urdeZBJDUhnPfOgH0/lTmEVzrL4qcFtWhMI2uUyvl1rdnReLa
TdDvomwkAL54/y4INJqh1kqh9Be9Bi6aw8AuzFRTOX+gLp7Pqk04SJI6rzcLK8oZ
e52PY+NgCmPhhWmZAH/VOfJx3rxR12d/OAmrduGQuIn2j0sp36/H0Xe4KzKZq9U0
7CKde01fji3C09YJsH00Htudc2uunKYuE+OdoObowjYNNav9oQvVQ8dkPUdu5Bxv
qm25INdBvOnPopU0ruJXhS3fE79bqmsF3jcwSM5LSWvd1+taOefgkrgzHRYu/J5m
k/T8zjOme96++XLPnS+o5PowlqDzCa6fYHuJS99qxKoUQ3+MBEyvGpy3L/pj4dp7
SC4YiahQLS2PNGJOMfGtyMQ2/myKE0M5ZrGtsj6FMJ6wgq3gPJGNa1Zi8dfjodBM
zstxKMr/2fDrpYLm7ZgpBREqjy82i9+Qknig1bKpma3WZXT1LmJ1Zx9Mz9fWCLLo
mgO1NuNOlUMdM1EvQHfaovTSM95ZNITL83zx7ibCxg/rCMxJGDN5N+ssJeivleJr
UVFE3fuwCaSbkfor4J9L/xxMQ71gwREMthHp7tDXk9+BMF/+MZS4ia9axRxBVP0x
+NdHT32Wx1q1nX+ndjP03YpU9TuZ3SXAp5iOiRiOpXJ3pomJyLQkBL9JrYiAQfwU
sl7mNPXW8DaRPoNbxgQGd5clFYkx0RveHf1B3mt7pEkBkUBXNlPr2jH8V0m7kWEc
KPrkiG0ZrrzDEVykASujmaMS/yRYQ2RiJKwqbgxY2HzBgjsH+xHQ42uX2RpmDn1X
+ypU7SeMSC+lvhOfch0okZZIQF7FZ+Ofwi5xWh/OrLcut8oE8zSmy9+hisIvcC8B
gK5A5tT0PcsABz22bZucKTGjMvtnwaLlxHbqyMQjs078C0UJWd7qjvhMN9f2dS7Y
M5E7hLRWZb24cZXgOyErJHfqIyVLQ6N52o4OQboC0RS085SJVc8R3iEpdhSIxaJj
AjvXvcPo4+URDDSW5creeeV0cyWxCNA0hVkZzQoUaKP3OSoWQtatfLg2KUwlGBJq
tayjKnrKOvJ78TAEYUsDGgDa0gYApkcejwU4CDY41EFQWCGTjo0zLO4Wilr+AP7F
JdQ6kSe/ADAoYuo+hVKUH6cRkPham6Nnt9lypkp7+Wrjd1voE1CfYlVcQlOlcfI8
dbaaGGhcGJhXEhqaTSX1N52xozySQP8tKbV58mylrfeS2nvVVBTNvM+ow/SzDz40
Fzl3O9Eq7fhzrXued8OCnnRzmrNXdBCVTgPg0nWuzJMQe05lazs12rrtYbY7R8ij
mHp4WzxahkaC6BFuMw+Ga7EF7ZNCyOp0rHX8ECqWCM/WVWobfL0wFJJxKIo8UthL
Tfu1gUhKGKKY/5D2bSFBd/HKPBzcrHYK8HLJtUKT3TmXzkB8yiH8//fcTqZXLedD
aKk6rBwb4dnrL22cKAaEWfWOvlB/eTCTwgYIvGCrzdwbhEArWqpwkda0KCYjxJw/
lDdpZ14cluzL81t2lbH/4+aBSFFIfszTiep5nrD0oTFeVDSjuCJhX8Qpr6Bsr74K
+oGmRC5rGkV3DM7pRJw1qSNvUjKgFOc/81NkA3wlzqQPsHN8eFaPn58U5Dlocuf9
h86daW5ystaxvAUl35tKAsaqyo+DJ1dEhjRCQScPhHoN6nHD2QFxaqUcT3qkB/qy
4Mvjwd1vvZ2jH71Jm4cGJy+4hDx9AjMk6egvR3R+R8Ga1LbCUQFABCssqkVgqRAd
J8iSXW2IMlLGgUnXLfOnoMq1LgpwXH4nX8nTh6USGQCBZTwSGMAmO0/VGtXIKji8
Y1qEvFmqfsL1tR7duRMGzv5N36N/dxaP2Y5luOtCCpywC5b0Rlque1H7uunUOFHf
pG4y/RxhEC1zIZ5HSTTSvwneWYaBFQAwWAvFsBhI2v11RAbw32vvENuDh9iiRV3h
YPV5SVC6kaDCBcO0eZRbiXIz88j6boVSTjS2bZi/MqQnXX2OaydYFqU6H02A1fC2
k3PS5F/eXG3DL5pbUOYyZKbD1tGXwsVo3FfFrRUWYG7xz16O+zt6aMhkddbzyrHu
eaBzRSGDT0r/GKuZyDwK4XOEZ9YUmht0SIC9Y/zMPaOW7jJLyP+F3fJWN76r5lyE
NwL8wa2ywJMN2ta8oKq9L2MVnDhvUnxyk9uFofedFHU9Dvc48b3X+td2E3HaPwB7
9xLXbxvmSNq7KIH34q5MSgJf4nzlHgvPjqco2+/OL9FGmJVgGOIRgtNGVFbV+RjM
jH22GcI9tAqP+bKYCStg6WL+pB6kANQHxtJNW3QMiDlocevaUmEIzk0ADpUnsOv4
otFirnD7Oze64AepENYStjl3g8BCPibTcmBRCe4P6otGNPD91z+c9aWT3xESSWQB
YAExsIhhkSbd3soJiY+NG5B72qvbKYnXsZGqub9ARyfbYzw9NI2jk84Vdz/qwEuj
JV3nhoGDjPtssGeF7+UJrxJLaWykNz7jZDYIZpc6FsEyp3CnEOmC1BZI+W8mH+PP
e3U75md9n/75utQzjHJWc96BkYZ2ENpKOAI8vxYZeYsjw1FHiyCzUc8GyTwSi3jR
/N8JrxxSQ3yyN8PuNfKgiokxukQeEOCO+8opV5IfUN/rAVdj6wSDMTKSst3M8pF7
HVgRY98h6WxM+9I223LBfzpi2zw4I7IA4Qc8mLiq/AWltFfxNIlrsT1D889vPFWI
W0njkA7xujk0DuSS90U3DSFefrlwh4TeD5nsHuH0deKIN4PyNkK7PXLi4Vqf8ttK
JfDYrFt5v7yB/TZdhbkTByK+jj8pf01R1GIO4qmvWOPQD6Dp7IJqkarF4fbLrY6G
lZDECYOg86r0Tc4qJpJIjlhV/Ai6JlgzXNqkQg8T9RKKVCdYYMx1ylqdVrG+Qa1m
UxaP9YWqKPKzWDInk+PWCgZzqqcBntllqtGJSVh82dbjCqB46Csmgda/rZGNofkS
LHqWXo0G8J2g//hQFMgYWOL3los5elDQqdlyAEz1Fa5ulKH+L12NLd+h7/RqQrP3
6GVnrqGOL3jbYzJTHCOPGgLHyiJ/W+1rF8fUSKnaSTlNLijxpAKq4B8eg9AtfhTN
A3mp9Yv8IZBkIcfI3A+W8J3sK5P7Ve89wVNQlw9rcenfAh3yvjYpwmGVpTNgi8Y8
biyw/cZg1V5/KEthtJ6kykD1dlHlLLvfGBECIYtsvD2CEJv1M/Ilh5wh74DSyD2K
ccvqVSEVBJFRdUdvvghASGZzmQkzYjmpEBCPOqzJF9Ht39PGdVUL5wv2KCnJJyum
zJO2uk89HnteStvA2xQWOVPV5aFA2qGD1Aij5W69SLW2aF7CeQULGM8IxemQQnHz
wNDDnFQ2Llct4rz5u7F+2CYJpYdJtI9socqK8AEEy5bSp0lPQdiElWH5R2REKKKY
DU0Rea3+03ix0INAIPEEgzXxSXM1XlIo01WT/saGpCXyYb/hjSGhE3x7xoiUQnNT
6G65DiIwKr3SpInjJdwA5OA5pP3+GP6l52pkpWwnXCjMoc4z6FLA5j7GLmh7CMwq
LzFGtM8VMmJgBp1+3w9Kd+ACTWMmCoFWbDbWQaBWE6SrQ27syRa8S6qWxx0RZSG1
JUj9mpsyRHkuoVciDaGkAP5SRRzvw/zmv6u5wnyAGD4s8ow9DqWLAWd1BvfYZ8/l
MizilOYyx2q3hI/QEkQh3VrWOWZtvt/TlXDq3mIm+VMiue8I0cnuvhz05LdfY0eK
vY/2QXvbOBpDlqyY/zkOKwEvarBMYtfJNDMzuOB24u1+8NsRNCtUgQFUMUoi+Q8p
y5ZJL1GCmvVcV+5N6bo3MjuDfvGlOWAwnr2w1n1hif+XGA9G352ESj14vVVGna7n
98G9FjUtZeiuQRvj7vy84Tj1/FjhhXcuYEejf5eyoJj2q5gdvPhlW9SPo8Tg0lOQ
X8I67X0LlXdUM+pKDQXTB5/GvHMIIuRf9IQSGM2c0UdO+3Xl7vSJnVpkfq8e6W5W
B22wj/8bT7r6bXDRiTz/xm8G5ZsDFPSj5CFyWxR3aC9sM8AHz5btt0j4GaUqzTPy
QBPYL0oFWQ5auxGsYH7OHl5vjV+/gKl6YT4GUk6Tt1/AwGOQs8OAFZSbQggU3D/x
CcycN3yMTyJhbV+/7r3eXtGI3WpsLC6xnXQZDiLfNgg5hflLUwy0VDqkgQmlKBSS
TAPJNJdT1fuodYaJ0Yp96c1VGz/Oxu7GYIFaTfuMIeYKnMHHwf/lQJX7iIb6zh6f
LBWr2hTguudC1cCWu1Sj2Mrtp1rhn21Toyx7xl5DvQwCNmW8Rak6wNada80foRHI
tp5u2KTslmdEoeviS3Oen7M40nG8N/fYDRByCSs28hQ9HEj2jSkqyvtHREFxc8Rd
lZR8a64aBAPhKQ2/d5HgRJOKnOroa+e7bZZdYOthJMjer3YFJHaqXgW7rTOdlkqs
2MOytq6IFJS8Fx0kaL1X5UHrxjWkTgvJvsR2Zdy20j5/eKbNFhJFqzm7VeyHS0Em
TSC/FpT8VyyPYjS9mS2DgB0iLbEDReqisGCHctttqIHnexuoRH8xe+EaEIvapIEv
IZ1HXm/1F0lLD/yx9vFBYAl+77qESLw4OQIzYse1uTtMpKTblfJ7ri3q+OUcTmaR
YgNNlPlFXo9n4iRuBvubLQbP5BiiEAbwN9w+eYoMaGA0Fugh4knfvk7rj2geRH0K
+BBfCDrLZGT2cQ5equasWn6tRQgTnRxEOGL8/gi/+3Jv7ua3tw0/iGNcfrEgT3kW
FMjRVOIOfq51yRa4/2ONULsCvjO5dpmefAh7VeBilG15GRjrbIFDX/ydaq1BHwZ7
SZ+pVCkrkGk/zdIfNXYNNF6KW1WM85RdQfiG+rSyj29p+lbWWnz3DjXVwY6hg+bw
Y1q1+SLytQaLKfPfAQjj75gNxX3cPgqxvqcnWzg3rnm5R5mONm8eOwYeXnFOvnUT
GQl+xKSODTl+93UubHt1FOrBkenB3wNqHUOvHc0WnGZ3L4WX1B/KG4Ku5Tf92iun
sa9yYE2XCwLPM6EKc5RqPLMkX+eFb4DjFvWPBCbP2roaf+cK2AjF9ALuuX0h3o7k
YaxLR7+9AEUYkAGGMtobfx00S+ubjXMq9/GEhtZ6VxftdBuoN1QlZcTOvfMBw6eG
WWDUwo8wLUZSxM9Mc16Cs/t/547GJouXJUPi0TYGKGzA+avNweZ2whGaLtjfO8zN
RkKTk37tXxk9ib6DPhMs4AMxKNtxqtctIMVErvtXOjhDclVCJ2BRLtN6qqu1kZjN
HgbhGdvAF/6qyjiR8/ssQUAg1yilW5yDYqqUO15GhrsCZNfd3Afs+dXhZcFsL8oY
3HzkNscsC3VSCiY9jEPAh04XLUlSeTixECefMzslB49pGX3xX+mmOd0tCKm/l6kq
x78fjgPyhy/E/DZeiVfRrEiv5tvVXTJ5a63E3Rji+4nT4E+nxpeozJpqG8kTjSjH
3YuUujrpGI32ZqbmD0AcY6BO9wnAKKFAr9qoSchmgjrNv3m+l6X82bmvPljXdnPe
NJYKRz2q7edhtl7qKbQTpjna5mOismB/dQf0duurLClmGYy72OxrspRmkCo0sf8b
rI0eSzSy9+8syJT1icslzzhooFTLB/mJjAFRNWEnw1gNZFXZ/CynoBbVz/cYC/mS
+KOVpxiMPiCx6m91cTyJT3an1OL3hbBT1f0xEKBrV4sc+9ax+Ve3ftNVUJ2b+m14
9T8xMRzmoG1bUQ9EQDvk2E1ZghH4ZdkvJvX92B4DnbOaZwIlz8sTVX8GxFytMt0X
wRhWsMBDDRKoIWqAImrqi03t9TcVUL0eavAA4USIQmDPJp70zH+E6vMXhTGltzGe
kvz9ykgDPdaQb7zkBFl+yCGyjsWCL3bUb6qF3g02LMN2t39uNrmz+TkkTwCuvT6c
6dHJx59UI7WyR8hPTtEVYaKj2nZcUpZpbF/AbFwgPkusuSUhTQojV2kynFm0Hrtc
mEaYBGmI8RuQYGfGMYcuz2N3GheMAslXSZpgd3Lj8CBR/eRd9piGdlzPKefgEq52
Vq/YGqN4BJsw7krQFNXT7ZY0KcqqstjAyzf2A5HY8pH/QjUzIPDJLsRgLmNn/ipr
wZAlRXCHLOTCnOEUJ/MHIDCkTb9qYOOpGZhckbe4I7aBE8MWvReK83/TIlfmmIwH
ZiENHQWVTaVGyFhhE4XAelxcaN5MdJgtHDYpqtDoPhtWF73nJYmGE4DwSX2nVJq8
xC0O/RChjWIT/CtZqEKqtNkAQIXjsy6T9CQ1LA2WVC4V224n/qyMrxIcbimYjPaz
trjolX0ocWEq7M4U4LYntb+U+3jKh9skdTOUXyD5ygWacccs1TD8SxfSYlnqYhf1
9eyPCdfheNl4hYua+mki6Yi6Z0QIHApsW5HmfqKIGucqgfmoxXIgQ2Mx5PUfCofW
UmBbIv5eJWcpqr8HD9q407LucMlpfaDbjANVHcglP9u6njxHB5NdXf7IyKYD0u/+
QRyPmLSUJhux8uGroKWrgQAorGlBHhmxDSGPW7DT5gEZu43w2lcJNBcvAbamec7Q
IT4VFUsEhNkUqMEPiagvY6MQ65ygn7bjknsUvLUvAuu9BMLVNn9iCtz6CxuCm+if
o25uqIOWKKvBfAVtW6Q9Cr5L5pz08DyjH4uaUZyTrEXBzIdu2u+v0BlTxI66Xfuq
INEL3tFKGhjj71obNYos3DDDnHubyfC8nkgKFG/zvHM5Mp6Z2S8mXUfItwlBl5Rl
lSfyNO4dmb0obBiItiMKSvs5W9QoBuHoKLulCK90z9N6ZnMKl5y3d33OhHdawNOM
fzEKfHNggAqyAo+OfBIawGMkhzfZAxxYvfaVfF0kz7m4iDk5x/C120Uoh84o+mLF
mb8lK3YqJI5PGFo9I1YBZ7ZZgXGxWSUHInAYv1Tps0S9OPrG5HcdzeO24TDPvAsL
Ukle82kDGpNkWghzM7sjVXjj4012EG7UQ0IYviGE8ISDs5au4jcCfZe7TdEBtLSb
TGNMwqVlPLZgQqTlAakoUcrAegbM5XxmmiasS43qVQgRsEqYvzG41MsHLrgP79DG
SOEBSdeyQGIK+F6RULFNDL0CthiA6H0pfjgvDSrAE/VxPYA2T8JgteNaKKBgENAe
IMyX/atRo880QGaNgaXFwi8CKjVoKhngqLflB/FF7m/om13rTLK48iG2LaArG7Go
2fTzGkX6EoIMYEl0WB+Y5fTt3+ep1lObYAk2ezoMQ6h6gcklgpM46gYLK9kTyehf
j6YQBlvqJBH6qTx3hZhQ6cevktCBZ2Dxyyx04Tdi/raoCE9IO8YrUE6Ky51lCfar
poLmKF7/H7Vgvm+nDFDqFmfyq2I9e0cQWEO5E75Sf5xtPB+4qkBwcB1ttkyMJym8
TomvlSZlmKKup7X9CY5X7bv/LYEGG7x02jDxWXLkLBiGevsdoeP8xJ0k3X7szXLL
hbD2Sy7QJuEAqfz8BBPd4FxAZI6MQkwb3Z0rEl4p4MM7rbMAEqSN+rhdXXJA8WH0
UeUR5gxQdoWf1qS18HAqjBU2Wo73VHKPP+/7sQpy5U3J5LsnSlJpje25nBL+w0mJ
BR8lVS85VS6eX0sNEDrxaTcNCpfG6OX0bMcvFkE3MQGUdy3/FFkEOx1FXhyTj6u4
v0UMFkYl8YSoUSDa1ceWxw6uBnYQj8um2dY1UwGSM9SWJGLUAKA0rGJVTFXwHYy+
is4vrfPFjCR4kH3DutUHSUyo/14EYST+KuQQQf1J/wMeuNUuhlYxpd1L4f8jrQEz
tfjr362/rKqe2uJYoOaN1hS0aaLwJ+g76wBvvY82tOAhb0JAqv9yQmNbqIpXTZTw
VZgo3g4oiwPDmBBLNMznjc/ESB0LY2PYDouiRDL17UodMsnPW3sqigKxodtbvgEI
3pf6AE8A+BeE0esja10S2uLVJSUEbvwMzMnw8iNWyywFBS8lu68g46V6v5huC6Yw
RTokiYNCwl3OOriqttBHmbl5AkK5LxQ4bLBCPy7O4k72QYjKLk6Nb0y6YpTtq6Pn
XsUIYUuU983khns8No5ro3n08vjmlINov6PA6Zl3B0j4dwE+uI02AUwLr96a+IqE
oDO/vr+hXMEfNFgGZxqFwvG5PlqWYWRbzYoGZK1SMm8dUqZwnTHcAbKiaf3pYc9d
4PQIhui56mNHDfb2oV8e99e84f9C/5O2zOgTXju5ZBkH0pDXtTJ3/J8b+G86IWS/
J20zfCg4W6id9DDkJtuvsoBiCd0EvvzfDgFGyrGxHCj/UnqP0P2HhY4DCNSDItC5
edj3qhyqOktdyb28+oxpr9L1UESn1bYY98u+uFFnrXHa04ARgiw48Z3Ckx+0D6yk
LTPtpEZHxhyOKN29gJh5U2H1XILxdOcjpO8dKj/+WCJQSjx2I98wIEQsD/fIOqLS
FlS6OXyKDEtEShdFlFefsfQZtvUBBfJzyprf9B9K1ELc5dd9usPUcByDhdIN05nS
TfDgbwq/jpnEQFgHmHPh5RsKPr3KwnleHDwsYkl8I1uEEV3AmhHu04NkKqC3uXeU
qVQN29kL/a25y8fNET+vaZneUJYd/o5J2Yd+S4F5EBu7PUtcOw8GiyYssdK2Oc4P
aIwmRb/6fkMtKcB9yBqkIPiVqbey51bUBU48XouwR4/TY2eJW3DV/v/wysa9Kvam
2yZ0RysK9w0f3eSmOrbrLe7nAr047cr2X7yXqSE7mEj9ZQ8EyK0W+R5Vcdg2Fa66
2Q4do3WGbWyiJL6wXRfKU6HG8x+O4wpOAeP2Z8StFzNc5GGYBmJfi0IUsYEAsMfB
VZze5o7sBsVRElU+3sJF3DLIHESpSQbF3vmuShaOAx6LxUyF1Rvh1hPpZD2phHsK
sckA6HgwZEfUd2SUSRVJVC6bKK3b/unjyEKU7hslD4D+bpKdV+87SrGtkU7Hw4Pp
0mvq9uOeY6bxV5PUq3npxzYJfYsiP0QrgMHkGzXzTlG0J1DabnAIBn0b4uLiIGJA
fDthIAMHMUyFrWmvgQBuHJyzrWzCx/1VZaZvk+VAE5iBDHngzxB43z6oq/lhR5q8
vT9K0y9y0gyWyFPOH+m79BP4NHx+QJXvWpOobD7BL0bIZoBOuHydPEPV2G8yJ9Y9
vEZiyxXJRZtR6lSaoJNvMelBz6VBPXAsHkgPKPng47DmoehOfzpuT+Bud5qjjInp
WPSUjpsIFpYbVkY7WjTWN2EFduiRSejnmcHzjUZTAqVNaEAouU7hsNCqGuIg4aD9
t43B79+e3KBmX2DNNv2WEiitZOx6dvtJJNW6tPsUnE3c/vVtji4SUGrdsJQLPsT1
GaYhv2+jfNZ5EYSH0uURtJBllRURl3/MEo4swlK6pvksXvWym+X08zpw/hNf8lmW
xPKY9kgXEhZPC+Opm92ZTOcA36Qp1ehiCpUAvvCmDw6kKQ6if5Tby+HKqE5Y4SHW
YK1q9lPuCEASWNeMecVINXzmTM7IQJDHaPu0JemaX2ji+8R8bVMcyUX8qkW+ABMv
Dm8nqlxKTu9YzLOkfAA3lVtW1YETTeMEUWqm1BO2bFvK6legk88Q1AnuH08q3lNk
Gwm8nFw0fMpwkpdaMXsfJyzeXOHs5hqI8A3qcNi1ts/KsMWFOYKhDgGkPq5Cft4a
dM0/lvTBNfRLtDTRFaztge5uaHyvYoG6VMmxk/ep0DYz+07Y3tyICmP0tk7OsEhs
vkNIiYoaEl4fWEWhAMcP/oOuwTxZqoZIogHPQuNrDIdkx/G7h+D8GG14VXF6NeHA
Yxkpd323L+EjjfiGjtXQmpxFMYVLGAamTxCLTsKpkkQ2x7LcZCcrZOd6mzNb8uxX
y6T4XA90Gu1BFWCdDmYf1xrArSivv3quKbpLZSHwTHpuHlAblFfsrAJ4Bvfhrou4
JE+hOmaXvcIfX3taTgZnZH7xSp1Cw5CVcV9AKTkYqGR8EWj1gTRCqOFagrPMQf8c
YqLesWeHFe/HC4M3TGAIbkR1Xu4SU2l9wHNX4urgv6VPCzBFSanYdm896+eNGKnF
iwfnYH46uaHjDgiWLRZrAga1i8MppJaifUQBTv9dgmBjNVzY5vzKR17m10aMZKI9
sTW/Y52O6vjM+C59Q8FXe4IGnjEMTND5PeTmNz7ywKSTf6UGfHoq+R4r1KY8GUHJ
zxR/NNScydn41hLUz4UfyXC+0vdaRrf7a7Qj0xmZpL56CtFZf5CNFHHDlDd50tMq
SVK6c6zFE4qduh4UkS6DkcmlNSnH6NB07tjmtTfeEDJgaTQWY7XRKOgvnso0j1cn
NrrabhBmC4x3b6MOHwAa9sxuHkykZN0n8Lv7Se1DQv1wS0/XtAR0D5kl9HNjVEJg
txwn42T+OcbweekEn89iLTYdzZ69oOAgHr2n0k3HSoAvWGweK9QtvaE0d5fYyblx
6oE+0dGHt9mi8QgCill+egOogWPecTy8GDRiTOyuIcW5G7B18Y8TQ66QDXNAmBTF
595hRA6lj7DC/DO39cGJXiIb6/6DnhEa0pwTt6PZIacnmBm9fWhOflZOz4U9X9nF
EzjK7/zG5V/tHDR/Dr2SHxInZfrFeezL1YQnaiHhk5bGZFYsMhP4FIG+Nj9eADEc
zhaq6kcAKcq8zXcL2Gf7P0f9oIKgqvWbhOvQlNqZ7mWu6CYG2qnc+XRlpz/tmKxO
tMSvqYzaWQyCxlau8X3zqFWs8imCkAz5KqUGdatEvI07esVxoNYFwqX48Tx2A5dV
RAhJsiUnLAQzmpvDoLluZdnvHh1cZXw4ienNe9sUs5Gjnmo+N527Fg+kudLDnWig
0VB7dEw5s6pKf2sZjmistE2W/+jWUAq/6EEGnBeFjL4+xT68sDxT74INsQqXvTu8
GbV92Tczu7veNwqcO9GhvMNsLhIg5fLFF2JpOboF/hKuXvIY5kzswh/rK8/RSif+
pQn8/5dqjPk01G6vxSuH4hSXspBsRmeG6FD8bBQCLd2KkQORjws+l7NmDWu0H1d1
IOcTotoi7ZyRQr9GJN27T+8m3yn7IcALbAwS1hccMPlU6WWFkOKq9DbZIM5LfO71
DSJHo/hEfgnYiUnfdCCwnqK9dd4itV9SPiMcLFG6PTCYXuZPIa5ZG40xFChpQ5j5
1FVJEJeBvBl2vonPfOfeBBM6RdZpHJch2SmRki06klI3b5tcMJVJbw+eCRTWbVtB
mko/CKr8PkFm0m1q4pP3tg/wYrQRY1zdNpItisu0R7cFcWGn48iJgc/a2/g0Rux0
r1R0eBBXPrS9G+FVQA/ehDBEq1690oK8kEVvdqg27ZKyAOwXo6X4UmzEPWcTClvM
lDptfuf0F2JqruJrgoTLi5q6YTwQ+KU/6CdpE1UWRE6PMX+CMx+VoNDZ9YtKREeC
V4dZ1gW4ayRLowU63xfoG5tM153fPMvsf7uHydfEi9bu8476aIyFLupDd7dSVG8n
UaZ6mfzqreeV6Ye4XcDrrj1nd7P5I+uNJciEc9ovcCfv9atsOtjmIeDIYM2CCPt9
o18tLNW3ZA9G3UgomRIKeJ8WnpC/pwdUT1RZrsAK1RuvnBcU/nPX9EvRrSA+T2iD
Xm4S4NP5RWidv/Hgrm3zZ7Os4Uh1L6hPPTyqJDLO4OXospit0Kvghc7mgEN4tJxT
lqKMblPk1kfleIGgsBcHaxBZMHbKRWyYoYhnNGF/AZjlcR99oHzKDKbKTPzRmCsW
6Fj6iuSgKiX9ea1MfMMQ4ebLWBj/0Blgy8Avdw5T+wgqQmu4dhMqEPCA9vgBamjd
Ocw0eHwqB70xEPWYKFDmb+tI7p+PdVvCQ/6kvUQ9SQS6S+59muwAC+wWDCHqhSt6
NN/qzkDGo+/D4eEclemJjk1B3lPFR2E/lfgfTx4a5Lu8bqcbkoSZHnOt64cOMxrw
pW+bJAmy2pi01hjT92VerHj24eu+l8aB3lSSGuzCNrrlPTzhL8IRe0bcrEFHyJM6
v4llcTkplXnivi4lRMQ+H3M8G2udP7NM5MRN2IYGSQ/KjXk8fXtMrcEK3fdMvvwr
GMGbDBw4BeUjHSH50Qc2RczFwz/7lEX51z7g+K02w+VqHHsFaNcAZsWcoWc2/TL/
bmwwuut0DiVgrRWoK3nMpzLPfu6+qPBArSw9PTTzBr01K9oGoLEYfyCzAIE0vrsa
us2FH62BMn3B8TOmITwglSayc0BNrLSl3KzGbSJZN2oNQNlt9R4fcMffKwyaB7ZH
QIqp9kyj5zO6DsIHse/a7DhfoJoUqa8ZuvN+HTFoxrhxiRP8esM5LKwD5tkOsUyZ
bOr+mjLD/lHmHO7h2Ykjq7FrYc6O+rpX8ExEG/9L+/T8zhU8cOGj25jSPc8NYBBs
Ti9E0PgyoajNQcpOHF7cJNEVRNuaRArcxn9L+jZHZ3UU/ZBA9EY2fRnDinskwg6d
Sdj+aGe0CRDp/MstPEIFx01wK/U+Mgo9EzxwZWPxLEOoNk/PABd4Uys91ILyt5Xf
EE4XFyn8F8kkKFcHybQJOvwdAnqFwCa2KKsICosd3KgQONsBUuoWdnIOfXDFImpu
hZgFD/Jt9830Ae9oDbzB28JNF5qt2l3JooAEZdkfCs8NXx+Zmf2YXGCrvWQFOVDz
0bPp4rfuyyPwEiKiqXPyI62WUYLaoodYKV8m+mZmI6YfBwLdov5dhKR/JB+BDQI1
YkUdcGje5doq+nTj2z5Ire0r6ggoRhjt2LM2qVTn9ltFSs0Gjx0iKF3mJAphqDvA
NFD/altcEfIuOeFPxqoiTNgP6Bj/uGCRzG+/2x2b3/Nl8PwlQp35/g8JXSr+QqPG
K8oLCIqP8LITyjMaDI/eghe0jWDGEErUfhsO6IXVsLepC6sNYw63/lA5OQ64o0mh
q0SR+mBx7AbkSgzAzViDJtIyJ8A59QUE6/iMXHI9RwwbJHHWzZhlkzWCB2wbCaS9
v37KB5Ax6+usHo4Y0b6wfvIke76UhWHO4nZ1nG+883IWOE9/tHKZ9xcD+YeTjAwp
6IgzpSZhYOapEjkHxKOD6/o/i4McdwsUkHCMCnnZJS6yF7gEioRUe7CmO/P1xSyx
qdKfwUc9Zg3O3wOGJi3BbFgZ3cxQCQi2TMXB6YK6XC/jLWCeviBAMlC6PUtD/Hfp
is//Ldh5PwB2Z4NglhUQLmgw5O2wEeeWGfpU+eMQ4sBViIY/aRdJNv7aWHlk0Nn6
tLupcFbphFbYYDnjGGA+PkFN9NCawWwjrIfSq8NKxnZ2eubo0s2N4w38BZgcVaCa
SSbLF7wpOpjPIQN96gVPZABlZI+BCh3PVIOB08Gm/eM6a3iTUy2Uh+wFL8JoVjqg
L3k3Qt+iUahHK07dr1feJ6+xUxG4holaW2+i0wqXQUfdIYWExvqAPauB9L4CP6v+
3Oh8RWgyk5izQ3ZjOJwuZeNC5zJmZEWS8hpbfulh29Hk2OGg8jMXy2zupE92WI/D
lXYY6cCmKcJknM2ftmvSP4cy1IxBOvmhYX+e/+stA5wzCb9mILmU9Bojlqo6tNhk
b1qYai/zp2iFooElDDFWLe+xDPelD45+NqPDCZ2XpyuQkB8Vg9K/Ngy6qMi4p/oK
JPqfTCkd0KAkTCLnKd7R7utt+zrwpviutexKQhyXwrpX3XVC+aGRMsB6baeQzuj2
ABd6kf8L2Tnfa0g7x6Aq8vXKP7LNgNlkAULLiK6pmYCxj4kkf9apLIi7LVz+hpnl
oQJBMkh4T2GIAzfyuL9JXTBZsOmLTYq64DBY9rLPlqwATENw8RyV8ZB3ZjiMrVFf
1Z1zwLdLnl3t1K/FP6KpPPckuvIFN1r9hcJrNIChOoeztjkzg2ztTscU05L0e6r/
Wwj7KmmFVO3BbDKhQbJo+M1puJxw7VcuOdMN9lPVVjpuraalbQyCPPy+nmJvlVbg
sNPnlKGMZBC7O3ys2nD7R8fI45eRcNHjaeFRD7oiWX/fLnvt/rny2qmqiHTf/uoQ
VppdsDGX7PQyH4JSXIdu2Rg1lq5hjy3mxw23nQK1SEUvD3+/BxDN+25Jt+wQGDRj
AunYqn03a4s5q+pjQliIvHshCCUfD5G2Lp/4YBIPJmJEl8Jma8Hfup24TmY93KJZ
ELnP70ZqfxSPId/S9SRrWd09RbkfSO6EGP4B+MKcLcSlwpkygNVyiwxNn4nTS5B/
Sh5v/QCdVeyXlVuI72jYZMU2eoqa4U/5N+m/DVq8Mp/IXhqyWCwQHh6Lcgl8id2l
zf+Sbn/nrNyuu9FNw1IfHknEVufukSManwql0DMpBEnC0BWfkGLkWjtSfjYNKFFM
MvNFggjIzP25P9jAEcZRuHQMndoUS5sCbwOMPhzfCbe2NDscQ+eFWh41aUEaqBEf
cSKAOYhbaKnRsDERLrk31efmJnxv8fgNKRmD8EkhX3MR9BcvJ6Q4DFAKnbuRtHNk
DEo5dElPCW3DW4RIqRJZddtJ04J/pSludS3mWdwmN/C0hKmF4ekFhL1heNjBWfKJ
USLfEw1BbBmB+vj9GEg615RA/Z/dWCxVPIQ32F6jtytYFr31bOsqZ3scdaVMFlLM
HXGeem2I92cNqVYyyftsMjTSDM9aImT0LWFn1PsFIuBpGTJCH/V0D1mc/VRLPOmY
w8073lmYz2mnj5A6rUfRAbmeR+HyQhNzmOf12kkyrcIMHR/GRaDr/i+Bs/9fhxtr
wzVAC7r6kktJ6/917nMvvcUG1ScMIiwpb1LG974qNQZtttntTFuV7MfuRksRyB6L
/WjN94D2p0Kqjz7tdQJZw9pGwjMURobEvEqlqiGeb3/Lx7nSYJjLFmh/G+OlXUkT
jOj9Qttid9KB3SPDJJYW2LItlyPFbuXpL0OeKasYHMYPLgzrYV5qB3W/QgRRSA4m
jE6OYodNFE7Z/q0ZHh3GnhH1uEy7Yav2S08pQciwgXTnQ8fjyKtdPeNWB8MvZAl1
7QZEZKymZUDr4k0Ct0RYA01tuh5XfALZWuqBBj/zKLaqnt56jvO9ZeHlBSSLBOfd
RPJF2iAVBe6uC7yQszHUtf4Rd9ZqYppiZOSJZvX2W/2VkGOLuLvKNIhmmCVMxF54
Y8vd7SVeDlcU7pRYiOwAdQALHX8otfiMoY9YMCVJFvc98S5TV34wWQwTG/RLKg9E
c6MZRhVOyJsfd/tLAa6KDjDZZ4pRhIY4kDPGxNygprPJFxG2NRIGYC4Z1TzY84bU
FCxCyN60aa8jo2UaAA8ZDP72K2tKzjQtyGoE+6w3XlcIXDubMLp1fuvUHCBbk3QF
6uADktqzxT9W2+dy8aAZY1F5i9UGeBy50MdwZ8qj543c1D6so1Wq2BATyfPhe9m3
PXIhG8wO6h9TpIvSujMpp/Kw7Sl+ButfrsAuU7b8r5ByHp/71rgkuhyU0JBi/HHu
xiUy7fi8GvhCF5v8fo6035MI4G4u469KC5L6swKlAEHuNvz3qAMUhAnAaFYYC1Iz
7ke0TCc1BuvDxkJ1fbcdRLTxGI14PAywyFLbz8Wh4Qt1Ox16NxfGD+315OBb1q+s
gXy/EU18DpVJ0QE7avVhPQgFqlsV8R7NH5AEasgiHLOMvFtwcli4W8GH5AQE8eLT
O1HZ/3Cm7rYtpaDg3pn0jwmjquk2CKyuke7chOO2phIFbPrLDDezCBk++cApNBJh
ZXEpDOk2NVBsidoBXkAI+tQWSdjgSed57U8u8/EPsiRJZxJimlf4m/Vve/SqeGzI
2BkUrbjh4dg/iuYvO0BSRGjgBfNDCazTM/KF2qHBJ0V6Jthln0V+5qOi4J0hf08N
MRTGmgPKNTpbLCD4Dim6SQw2yac8brpZXfsAG2pvFdlnqoKNjs21nrCtDTbVbBzs
wuH0Py1T4LmvfV8r84PW2pdCZJaTPeTP/LF5288uLhJrKk9MVFEwgjr7yF5FUrFe
6xhacTWEIGTPbuUcifQ/GPVqu3Xy1SdTA3OkBrlMfHr/Ss9OH6m52zmkOTking2Z
lRwOlfdNhCWsBtnnyyGvXhleKpIOPhbmAy3RhhGEtT04KQnMIru3klY/f/y7mhO2
+CwoxWAxX1e6L2WGKt5VR8LC3h5wA+uFUQDfqpW2lLa7RFEAlg2pLdjvROVWnGDr
snhmtGs87O1t6ty7RqG7NrVMn6qm7vWf5zZjoCHwSFA6qzz3MmegVuRZbL2XVKi0
C5ZJsL6D6DvsT5HmCb5bcEGm1457kvUuPM/E4QxOseWLHh3wDY2/3YxLXf3tP0Ky
ipk5RELu+H3RecNu53urVetWH7FGLrz4iIJ1cHuuNtXXEaZM+E2d7deaVeKQu00g
YV48nwR2OCcNV458tdLyTxU7MPFWv5SOLu0RHGWJNufScE7WgYZGOQR8psZKf4Vp
+OjdkHod9cGuhUX8vAyNZB1WzZ+HkwofgVOwu/PP9VaFk/p1T8GWlWlt2QuyyTx3
2K06QfCEglWZVPgJIYKL0jcN0pAS/sFR9DToI/3Bz2jfSMtlgTgISGj1+pCGFUhJ
5FT2nfmWlNKzXWE1qvGART/Az/Hb/Hsbr6SIwV9LTyPJaLcCXfYXOwb+h0aJcmk9
kb2xIr6mKjo4IU8mWw1wZlooaTRfJMTtydebXjg7nxWRaepnt4yAWm0O8cE6SN9k
20lxmt5SNsEyRTaUjSROxjErIYv8ySwH0AVBohkOu3Q9X9pe5Mm0BbZSDA61XT0r
4cLLRoCCrSBpNZzmsxsCJGKeRA+x8JgMx59ngt+Z9b8K+u8XK9mVeEpxrymAd+RT
1uiVcf6hc8e+dGxxHM+Rn9FffmRavUpY/NXMxrDV8+ulxXFHt9FKBeukECLqt1Py
FxZnMoSK/GZO6bgCcCSOtaOxjLjWjHy6yvuuxysQw+RQiVucvMQyE0c0tmJboUK7
HErDwnRJeknt4/n7QelIOMZDhYSgN4A1zvSP83jLfaycdw6vQJnwKjdD3ERZSOmS
wL83r2GO9GaYjeiCiozi5v2+4hcheMXCYfs21yZyXPZa8/Bb66RyHk2r1NZEwdwl
AgMOGVJaCn+uvTwup3lMMhxT6PNgFLstsq50/BsEWDZaLkDFqEx8FjQgb5fmJ/Lb
J2VwzeJnbCU76hDMFEY+QqkzZswRJgl2kWD1CpHpbuzzOaePJdK9CIAT1rWPL/52
1DdKStNhj6DZCiLduQ0QbrdfJDdJb7KX12ZD4zd4EEt+1zEvAYxM4TlKtDM/MBkT
P/mqOSgFWIH3O3kvTLhOvYVsoS73Ve3cSQIg2QuQELFXiqnQT6IRxuweqTOYOK67
Fsb9MzL6jxQs0Izel5YY1bKGBKZJG7Y+pShLRLJb7w2wxmUth83X5B/ZdOG7kQja
orcHEHGj87whkKc6pvMhNJkv4lruvVT2CgN5FeTvAMk8MKZme+9V59qTmoE93LES
klhqf90fuRmV2ceUYk2wpkWw6hB8P7M1ApeRljGVJtRv8G2CJyLlB0MzUa31SqP4
4SaJm4zg1QrGH7ZPu5Bww8NLV0qV19tSpjgHgB5L6f05q9Zxdz0RpxuTkGqOsf1H
8sGIrMudQpDNsvqlCkStnwhoeMVfhaZZu2tn01XNExlDByuOQzUuEXL+B0jSissh
iFTQQMHZnBwdarBNjWDFqKLnKFTcrZ1kncWdKWSkKKTbrv1UPjbLtIjMwfcDEBXK
KpOW77X0eFYkrcThabqspnnrByw7oyqu21oYuBV0/UIVryIWXVQoICMQjhsgdKVa
zP3N9k8xQHlSo/2wU+j5O7+SBkmAsbkprldfXrEJLOO0vku7/VD/hs1NG8CAENjV
pk8BeC7/MwlLDRwC8LB1+PZCWqCnWKZa5w/V7HslI10DZBlOsYhfULHlWUcCrI6g
HIVS3Dx5LfHwcy+GjfkGjDGa6LoOp5u6zA1+olFad5eM9C1TD7ISeLB5M9UvMMz5
AL6BYO2CbEAL3n5mN8cuahtSrVTFrqcL5sIyB1gh0yseYX+4B5QXf8Wdupt5iT51
cxcs6oLqvpl4dathAvZWKnDcxAjR7HwdK9BGRn2f+YvWmdroHN2z2Wfy5kXxXeEO
C7bMGDsUBo8664UM/pphqh05WXDBF1WQdzqKWkXIBKQuG1FGl2BEPqh47ov90PPd
mIY2HGHARz9cQZbRypXU4qHG1wSQN2P0/l24pMlfT5tZI6D9WKQQ0A8dbPwK/BdB
4GOk7o33B+ZCbCfz/uPbs1vDuelQXkvK5TnOlTrJ29RkT/8zN+JiveSMhcjWpK9e
LE1/RpE6Fa3xylRMHwVdEaem9w+sl5HcWaqXd1634z3TxENJtIAruLTFXL3nR/yC
3IprhXNG2VPdHsDJjJnHYB9ahmDCG3PxEq7KbZ//vj1wgkCx1Ed8+KXG6DOtZf1p
JfmfpNIblOhOMme0Wge5NB65kj350yNk6bnkfyJ5zhg6GyoAxTq7EdFhcTebvTf5
mABzPI8gS8D9SG/yZd4Pryggnm8dQi62ufpWI+ByAB20OnIPOfNkeWJhDBqGw9Jn
+KZm3yHnU36mfMmG2dF96FcG3X1hNDy/zxcVHWowvTVolqTnafLk+YgoJrqpFwK5
TjvjZAFDY2Viv+qfdUG9O19p4OP85gyU03bW5rKsqZ9u+mY86/kVIBQDKUNmTz7q
sjPTRWUUPY92gxEqdG8A2Ci1oWR9fTUGUVpvaxT5IFJhhaKY4nSrp93Mqvn8rtDH
HwdDX+OcBJ5DXRlWP6HEeWoGQUD28pW/VBaEbYaFxkF2V3rFNwEIWApT0rbzcSyj
Ly5ESEMIlaquDOXCVjgfpa+4cK7S4fj1VL3gNgNhppQtpNWtUfDi/gftCmbSLWTX
4OxC5pyv4ErhOIZMLdm2GzXYuEqi6AUG0SGbw+BYGcx6e8see1taTj3p8NIbnRUc
ckw1Kq1J1QAVch8oIyBvXcCgaoKbrbU5SaehE1jqBIV9fOa6CXMNG8ToV3ha1UeN
C3kEm7peh30D1/0wM2hav0Vxr77vs5sZmoWpucc36t8DNtPxXFa4pxVnDH3AaYOA
cR2mhdNqhu5cprVV0gMR/f0LURaBmA2edRCx0+wd/Sczj/LJrIhKsOdDC2BlQrtX
HtMcW6Mt9i4IkZduulAMWHbMN8Vb0tD/N/xgow8fLDrTf+tP9GDCxdH8GjoMPE/z
ftIvp/UZhl76cXRKEiMwCL4s7RJPFwTbkbYUDxXKvdTi8/v06es0KqWajsqe5o6x
63vn+9iZAf563Z+YQ7qKpCrrCBVy/u+ydnVU61M3kEC/sxgchBIOcJ7wk1NWphpw
tmhWXaMYhy9e2+Y8u2Q47b7eZH1bwkMQztw48kV+Q2vJuXW1EooOG8lkOos8GkyT
AYaUGCjbDw/19kgoszh2poa4gpOCBywjZ1BL627K191ETt1lPcHRLFRbuJ0KQUOi
3Gv4yDbAib3pq1/R+o5tOSzx8apRRl76lPC0jwxdg+Hp4XAktdnwe4+yXNmlQ2K+
DIRxmJrUSNaKJ1HcBBfWxuRMhRt3tX36gTCucvsMWRgBuXPHNjNuPZejAHk4lQhR
RstNIs/ydB0gXlSj1+tq7g3igw6IGtjK7NFWEXLQAyW42Uq2LJPdvcMtvgk6XTiF
lmoScDgp5e46f2cE4vH26ATTLuJJgf3BMieJ0w4As6Rdi/0ydJFjWxurZuQrDB4G
xD7JyKNuWjJ1mGLKqA0ts0aLXVBBKdb0VcjvrGfKhkTn7WrjxGTy6EnJbe3C12Vq
KrW9ehMsS3SYllI6DfLu6IbJHXpMdbtHWOl3QAunNfZsw8ZDsrYH7qrOifktHllF
20zQq9x9g9Q8cNkfQC8zzAQFCtj/BUti96fWpH+XZRAYqhIT2XXQNNe95R2VITvE
IT37Z1VfWG17Z6dUsYpzZaxV8G4KiKx9xMwQ9n6e7KxtD9L0RhsLsf3RIe0qNCO4
9PshlG7Qs8DgDYpkj/DtxCNcfrDVW49f1Ohns402oj7YZji9wYiSoGDOtNzBx03O
ueISq+eMuqXE1KBShKfiI7mxWPyesYXcRYqBHwWugoBEw0cKYwncOom/Wm7PZ39b
O3FYbRIOGFmgHpIyGDdRfS1Wlo7UHceVMh7e3Zuwzens6K1hOUt4RRVBUVSHiaNK
5objTCWZ4olUiAgWPHzwS8fiU3XLX5uJesPQbkAqVt3mXWvJOVnJIRU6yFlbGf5f
XES7zsbtKTlSk10FKq0uiIHCvc6z0u30REOKt44ykR8VkXUj2JCDVQDSBpikjqct
DvKAYDn8n4N5b0pJ77elluP14JMDoz/W7rds5MpHWeERVbSy1g7VagXB6x6qXKZk
uPOOdLwRDeq3RCxQAN2PROHFRXL+O7znLDnEdmAWaGBwFZ8aJwqmehlCoiQK+8ul
JO277u7l6lSvMa7Woyw5+qlS5ElR4LQLGPt/TKxqjoGwdHojuRVfJr/qgi2E6TrZ
ADhg8Je2xFafS95BrLFNnGhB8kjw0masBdYHU3m7sw1mfznTDt6/4HNCmtdysgLb
FdSq4350uejc/ZCURDZWaS9q0UV4gWM6ktLpJ0sdgCTPZ+lxraSIL4+LCL6EoMWw
uK/HtspnrBLy/I/9CPYyxyynBRbOd0v/ZbTgFPdj7wTnW17a400TQzutA5mFbdCi
c6RgSKZklM+oMJSJrlMaZQsurUJ+nM+cQDk1AupEX3CcQcM1J8tIGmieqtJRhsx/
UO5a3pglaYooeVAplNrf3F2ELs4qRNfKugY1j6PD9YwiFXSOCpjDECrUeMXSowL4
cGwsy1uDuOBr5AZ6D7r6/8uFwlSNp+kQi1Z9/3S4dpiy/w8YwroNsAuTfd1c7N4M
a4kd2LfgW9/aY2QJYPHtAjVJXWoWF+LrLpfD2azgJfvhsO7F9qUy8J0HwLLmcGjV
xKg/TD/A/SRpN93VjA06bas+gA6FWRy1/DptMAy5MRBQu29umR9C00Ylg+F/xrrC
xt1dLflDJqFNEfKdPslclvflg8V2LT7Q92bTcDJwNlWlfuCA/Xq0g2HZlDdV6TKG
JjVBu83Kj+qXXvvpd4cDKZUafKjVZ74f70Bv5MgLNOgg2r542+DAEVzP9dPuPa7q
2Gu21o+AX1pjRSPtx6hhrmYokuXUy7A98iO/CI8fVjxYmNZ2KWYE4a3zNFUd5lvs
qgX0uvXNIhcGvloZhPbSHsd6pbUbuwJwKM4nt3Jn/ZMkAM7SMD2VYjo2mLBB9yWh
YZXXG1aCH1vEQCX1QQr3XeLIBM89rQmOnGlHtHYYEJavfEfAIi5bV1m0A3JbV+Pw
E9sqwce7GOBhfzB6b+9UQibIe4I22VmuijGUW1L8eS0b2rqqoAUJ58I5j1T2RJKG
Oiq1c1Zbkchx8zVet4URnoKN6+EaJZ2OgDdfzrugLvULLQzR0VyUch4ooU5BXpH6
WilZVdxxSj+NS8MT69YczE193ijR2j62v1jvxz6nPX7rTEtv0n2C4IiK46q5SAiM
HitbpILNAOaJ6kbwnoBfMTaFHgfMSK1Y2r6usV71U8FC8K5xWiV1raNJZwYsRHgI
pqPQHAq4GF9ikEzas9FvGg7yWIiFi4aG1QLDjF3Rqmwes1f8KIwLt5rJsGy+k6BU
A0lcYu2ZYd/sI5AwBzquKpMcadgQ5UO51AI90IxYQIvsjGRc4GAzDSLRRP8DbuRJ
bOk0iV6nliIE14r/pfF2FQgfC+loY79DMvvSJ3ioa1uM1KtcV293i9WKzY0mUZii
ncMOhS5gjdJy+k+JMP4y+wAzeqnKgr/I2kY+aMAPqSrsHO79qEFIElE8lOJiZCUR
Cce/W/iI+adCxhKH+flwMtkdCad8MgmDNcxeqEquVwWwnKGXfajmuwblKHG0BEvc
cV+q8nH3BIEMT80sSctUzTTFOW7HdD4QKL9Z7Pq2NVbWhQAghRf4PJcmynb2t2yd
zdWQFMJYe94O+ARHW7LZAwNUbRM+RzuT9IBJtuc00Sf8ybXmfgQof7u/WgDVfz7r
YzZ6eYf6L/ftfoRGpBiJHMOKGY+IIrgnZcBzubTDs/0JGTFLezpy19yTp3Tjq484
QQNwiA+8ZPd1bP+LPfrEgt0Nn63drE/FdmlN/c0xoMpgp20582zItX4ckixxj9sW
2s9L6bxhj4C/EkQrYpxS+GCuZ+WNu5y6LwlRFy5i2k9OSRl8P4Lue/3YFZi2K8VM
hhoCOLbStvyI1qR5jbsjqwD5ULxdK35aX2OIyj/HxQhsYLhVr90+a2sCZtLuk32q
jb5Glt09hcny4wnsdXJ8Dd4YOP1caNRg7wqZl86wKnlPimGZMePdibI5EY6KW1Y8
QFJ/IpSr3hp18SBzr+4IuWFVxKi1QfgdHgjuGwsmLCOBUV7IloY/boj54aZgI8TS
+wOzbHHzXaHl6QcrmNxkrwuB2jCYF93IFXm7jxagFOPMJq2ntLdZu0kjeaYjVLHf
SwEqE3R16sksSUQBXd512wIf/aeWlyBc3ErHo1loNQW6RaUsTrVKepWq/u2rAtwY
VZIBLl4j5gNaQJy0hmzzk4dc/1YZ3NgTt3OOXfMkKPr6DwwktoOkz327frm858KE
6pvGbnHRlXGkcX85AJXh9cGgEcu8bZgrBbNwA/kwGaUmtahDV6XFE1SAfi6mqW3y
SUFm5e03pvH9IDDZsZKNO0t+tVsEOJgXdvHN0HWXOnO0OoacWWQv/w6n1QTO+11U
aiZZ/VNKCPlcftVCrU3M3eaeO/75CYfBJZvPQ40NNHLKV1mR+JeJ+WR2csbnwWoQ
hcTnFl4Y5whY+GM0uyyicdBDf9ariJZkM1aoG3b1/GsNoPc6oB61/K0CLlkw5gzW
+t93ZyCFsRAlVs2cIDVzWgfC164u9Q2uV15PqNzM5Nv+VT1jxgKaBLJSC58GiuDr
wQmWlxAB+Tbx07c7PMWpBxtXBfFnJJeaKS/7adI3/vYdBNRiUSDXKoR9MXM10VW5
RDAlwc2zQr8r0tj0Pqh0DizjO+Q+q4ioOUpzOWZmpVK19F9qrVnb/Ay4iEOLF14t
kXD2gJ/hgUNUVpSEOECeat/ZAqMAa80EixmUKWBeA1EQNKeriI2hfK5SWDH7xaAs
h6+sNCdHZLIw4ZjHh90wMYoccAx/x0InX7TZ4/fD4iTu1HJuNE59hZhUx5GyaGCC
6KoPsIc3zr1Hp/NT9XdcDG9MisHCXs1O5o1H1Jm55dOPy4jg7JeDErPSiFMkIxd/
FHJ5ykrANoUXvsJJI3HRQWOBQOJo8osx6GTXZynKp3Zhdcu8rb4sVT7fhEoMh6jf
RSIPKks0EcR04KlKP3ptV4eRBCLIY1hKLyhjBfaKANot3t6Gf94+GdIfc7Dflq7M
+WsOOcpV28fYsQyO0zsG2IrmXo1RFWLvZXif/CXdB+N1d5UVJ2A+2r/2KWLnnRi/
ZT7bpELVdK5s5zK6vN7VpGVqRQK+ID+3V5MmpT8wVcirDxawW45kk+QEs4WNt+co
HRgZgoYu29lOQmYlKXkTbaX52IruUfugAVqYxU3lLkCv01NH39Mqf9KI5fEMRGGy
WsWpc+GGfuQG9IMvWnnQtm7H/kDgI3rrl7A8y4I/2JQ52uPcY1t0h2tckqaHMimw
7EwRt8sYEnnf8jvIobGFz8435ED1oILc6nP0wnxL6zs3SkdzfJXNBW2cIqPdg2pU
WrfUXoMM2we3A5xaNAdzCN5jCuE8irv9c+D3T8zACexvtdoA/j4BnShVxlMbqATQ
1SaYDokgjuj9dxo5TqK4QrXzEGDal+IIRLT2sLBVfAJIJm1S9Ll6cZTPOtHFR06b
F49p4adUZg+0QPke1viSsfgvZyI/6wjH2yL8cLdR5kVaXFw7GeiAKA3PKm2BTGwO
dIGNawCDcQHu9oV9EBsxsbgNs+boXoUO1YCVZONLyqiXrII2n91yr960zl4F9CG8
T2tRWR9FU8AK4AOeGIroje/QYnRsL0hbc3AZ0QfSyhIOKp+tGqXupDzNh/XOG2+w
yAk6qX+g+MkCCV45/+Y/8ul9XmlMR6QjfYkdrce5SAhFPcLnNxN2x8p0RQWcurHh
ruX6+eJOmAkJEl6gyrmPpivKsM0q0Cjo9XXa+WWrgjuVIFkiu4hZEjlj+RrWEzPd
A6T1Ttr1dKu89jyHotSoqZtbtJPwFsPKYxv+WqLwcj/pRDy3U2oncLFoBRVhu+Iy
Y5CSV5w/4ExYEWFKvPwuyWExX/zvpEW92F9lSC7aZ7/vcf0SlTs2g5FDz8q0nys/
P38a0fyFYUAs9jMbWiPbOrLG5km17kxy+/ZrsNeiCPqhUYSnsdJoSrr36pw5E7nP
jpHfkrXsvkBVv/AekJQjEif/0QH4L/kxucjHQvrHayUS/W1UyAhXb3UqgJ1YarBy
JEBrgLOYTIy1VLVLilyZ0q8K1ExxD1LwsAAqS/KwlOj8iqhnh2emg5iDdni0RjRH
YgCn1n4uU2PJunn2vwVJfIDawx2RxVjk7Z4Lf9KXEza5qeV2i07DcjeLub3yFBgE
s73aBEAfrclWDzNLj1ObwKY7HkPGbPgtW0eNyNiapjhXmcxDjHzUJKqETbggvO4a
ZvzeV496BwZj9vM678wBUAZT5mam+TI3vtveJ67WSExf7y0rkI+5s4j7gHJgP/th
C52wqzXj6o1mkVkyRrUWK4/wPbhTFcb9sEQpAYpsP+8x56ibj68bXhhh7n49xax0
WjJR5/UWQUEqjoUkGzHEmoooI+EafikLX9VvJsd0azJEYumwmMiNFnNaadHw1W2i
FvfcLBSm81c7V53kDQ4XSupjLVIJbGucHHWAO0RUbCJC2yZ9ebxILHUDhb8i+nDf
pQrV/8P3NEgV1uf5HiibnGIxfQxldvVb/Gb91GwPf16SSarRt9yFUhYxZ/UP7qa4
OmY6fEkZguSoyhveDic6AxEGUvpIrk5WMttNIx2JYFYMVsayj/MkUniT3EVDC4En
OPoF3Pa0Asob4oNddVD6I6iGD6e/CcVVPhlgrQUGnkwZTjbWTSucUEt5l/uALrMk
tVtx+rwGjBRHZ6UZHZaczCkQSYFOlZvUtKxU2yHgcJqzmyJ6vY/9H3SldXvh7DU2
0plI6TY1lcOeceRRNtjcFVinuSSjI9luRUzgnXe3FLAqqFWmJf6pCV9kzAy+4eTL
S3LD7sPiKs7kx5PiN6vp8sLMPEF8tjJ88Fu4lBLVY+60Jf6HalIVBdk+DR5rMWfG
M1ZqEMriFu2EuDVhOhhajxdgs+GkCb/RIroYaW8Yw85qDbmy2/MvOM699RJgHqP0
v9YspS94Hlyad//sfOhrBEe7S1sKJJZmPXqj2VQgW7gd9urC6hVyzP7HV2a45dS2
MNusWYacXhwhw4eWV49N1lLzdRz63KXAl2c71syvD5RU+TpCFmENtJ61gGorfVDV
Ude/80AM7pCf/UNeR35I5kVi1NVKItX4FngRu3rRNo2NBA7q+HPNuLY4Pi/X4fg2
ko1ZZ6gE8OV28OKF2lxKR1vcyw+UBBfEdWSb6CAjqGty01xjhmozhtNWdFBcPbbn
aKjt6wM3YVsfEfc3U+n0ye0bwSRkl31yNP4NfNVcKMrDhSSN6sRrnhlYL1dhih56
bvbS+I2QXtRy8KtTfaai7/17rrXuHVA9oKw2kkSwlEBFfHDUMc360BRydt4xlSfG
j9lS7wsHeWpxNdSjVt/cPbdiz+02vGI1IpRAo5Yko+0Ati5FoZxhYIQpE8YCq0KA
66j/fOemxRDcWhJ8KVTtscpi9RpT/zF8W1QLMFkfT+oNj816HHMhdBZNp6VWvyDh
McdWJRj486SfF3OK+mB+eWAJUwlnv6+rNa1vkBz1SLDt4dQ2hhj2gGo9P9DyK4jg
fsdGEPjZ2I3YNvR2/KYd7pJvUlKJNx3TA9YxZLda3kHhTGvUqIsat/zTH7VpJi2n
r9dk/pd8pZlwC206hmtB983zio2UgFeXE3ATgDVCVyIEgq68xnM2tuFW5bTbWHx9
1motv1AHuTpuFipsHcrLvA2f8Mq2AYUqLQvwwB2fe0b9Q4GC619yksywzVvSvjeY
eKb8DL75QjRRTwHXT+9lgXE/K4XsiHVA1w0Lyys7PNlKhf+7gMZB9YEFvw9BwKvh
WryInbURdJa94nlxLJoYvM8Lhq/Rjis30i/3TQZ8Z0O8avTGTSmiA3K7kkxbMWcc
zqcC3zYI29WtpzZIvOj270E3SxNNmiV8uZhqTnW/skem9IXlfGwyDrgH9HfwrrqY
wl1oGUqNLbrlVHbijS+k/WLx6DdRg9nkC79IPITYBKHLwuNluGMUfUIB9yS4s7js
yNr+U+SFfNGi/07C9IYUpa6AJT3eVuAiuHZvKulfZCauZvLUwNVymNRC3eFLeqmb
zCiEip9d6Hg+hCOL/eYPvachGyKKo9WK5UD4+SDSxzvmiL9cWQ3YhOK2DagwL5MM
N6+wU/nhE/rZVyt5pTMoUfLp0W2a21T4ieZk2F7SxGYuS0uEtBMU77a9aOFyKRx0
5s8lO0PxInrxcSQmgINzf+Tn8VElJH6qrp9zmQzF7O/Vkcw77ZfltPNgkKij4SdF
4T2O2kwQrX209cB3R2wUo23ts0saF0gunsk/k60Nlzgr/PkbJF+UyeQF+kIXsWpW
1HnEvfBRg5wZK6MJRGbMHEO903oEtz6maOrRFM9czoVhhX/gA8GPLms9dOXdWnns
jpdcwYrtqBt2OLsI5c+K/qag0OcR51NeYoZ4XveMRW0JA20c0/WRfiMg02LarGyh
0bE0uYyVIWm67ReuXrabQbp6gqlv8296TH2QSipS79jVkbD4hgr0DEDknbLAY8XF
mLoR2FgW2a3Lst4x3cbcPTAA1NGWNk9WxwqOSNr0Qndi+wm4t+8bul+J+MsEecvb
c3So+ftwnq8Cx6e7mq/WA67MWZDOo/xGCF+7YttqYnhc67UWXWW4vT47yTcVf12C
w9pSNGvc6rRrtwZZEuBHELVS8az1umIsa7VqpnT2HI6laEXLZMgJRASj2wekGgDP
wSIqnoxhhZZqb/cJNcMRzzgIVXJVOchMWi3LKI74X5uDCNnTxgsFCJab1i6G03bQ
KWdu+bMcSL8ZHV7H7wySDpvTJ6hMQREd1mhwjKF6sscaVRZK53DQ2aIXGXazAAgD
Zdw+iavKlIc8H6g4vjlst2aTDgELkTp780uglftPXMgIHQOp3VYV1GpKUzEFiz+x
TXojdsE4iScJUZ7mwjJhsXpnVbiSC6Lh8f+ggXWlydiS1maKCg/T0Bq6mHSgw9d8
BuMx1vlkRxqGc4P1inJcOabdd3VW0GVBh+5nd8DrIKgTLoWuIEs8HwQv5YJkpVuJ
CvSF4AZT3SofpTt6uv1EFvQ9I5eRKz5d5E9qNoy8svqG+Np5gDEy6GHTTuqAwu7s
2vIUm5JQr3Eukfwzsmm6gIEKk63966lGyTqsf2ujFkl8ABEume7BTWBxAaIpmCSC
UWDM2DyPrznX4xheYkfMxkEVYzvAHkbp+PNycC0SxZSYcG3zwgS33XYdhzrgikPU
EiRnGji5ReEDeRobzhwqeQiYq7GU7cq3gM9CnSb++4dS2/MP4BxueFr9Io9fsXV4
GAuh5aeSaETDgYgFRZbl/Qj4F0zrGwpc8hXXfVO/gsI1d2vKhzWUxTRXI5W1tLnp
wz/oQKwHZT/0yiOrWeR19RpLvj/F6/dKd896EkLD3kRwdsnNywp0eZwxCuD1Rxrh
d6hM7V4WlgijIjWueSKLPq1YVsglvlKYHxs8r4XLempWW6r8J63uJJmvGi/SBQdm
QIUvyaDKIaObQs1oQPNH57CNduVAs3WAtcCb8TpmAuosMJR14WVlGTDkOtWgB/wk
BOXY/G8k0UIUPgft+kAr7hPdokniuTJ8FyndF0zOReRP+kIVAlVI4IXLE30AyFw6
aE1y+8qkF54FlFAiYGtoz7smQlaKFlDU6QfphCs69KiG5CrL/v3p1qzYL6540fdi
4NpHC2ltG98aFUk97xaAZd4jrY/xMfdxtFKZMq84oRUqq0CuQsaP1yTy6wDb5ZKi
9yfdWlsSHkw9Az5YaszySPjlpEX4iNSOKQolDg0j+CP0aN/425P5VgunM1INPJ+w
palzt4NcBE9Dln7jA0A8VRntAoS4yK9+zA4tV3mKCKBdKwhVyenIp9AKXTz26vhJ
S1RRvYHNBit+TgZzT06ahRhh8lVCAF1ZswjfSSiwlNQQV3lunRgR/O4wvomiQWMP
mDOfS51aGBDyeYMWHZSHuBEhHBWool/2L/sgPpyVEBlEIJXdVsgcXCWE7ZD3anGk
iQy9gxnvktx3GSQ1EBcEhg+isPL8F1j+N5WBsIRpCdbM0ULtAkqHQ4KaL/yDy2nw
HYdqXmNHJd9IqClMeXGI1vVShvSH9vXeFE/tnUAYk3oZyqNSe9TBIPhD5Pn778Ti
lJZ1DPWwEWy34+R5HXlrRlkdpuWJQpkC+CAZKn7W3RFkeeMPwIvpPNOQKO12x9R+
yeC6d8/aqnVBi6MoJXHIO1SSpmo5DIAUtFRJSUdlvgURL6VWx6qGzLk5VFjLDt1e
WZmdTI+gFRYTLzOZ1TqCZvWBFFM2v+/vHKTntLnYTZxXR92WW4NzAkOvYsbuhj6x
yj1VmIVRCHqOQL6i4nSov8jquHxJRzqVDBZ4fYi0Iu+VYyIFaWZtcrMppEWOLEbS
JASdh6A3lIetwSDs4B1fwZRe1crcesBpp81laMs4dIP0Srf3w/OML2l46rF2B8p9
6oNQTYM9JL9VHosiYQ2SF/FXiz3MeyB6og+2hZdcSe6nGbFjXpr+6cquxFhOOiNt
ZzWzbk6LoY6GuIRi9N+8lb9930eKQdm9IRQ56Bt41NJ3G6rLJcJynM8Y33Fq2lWE
m71P+CFiYm3TztOSr/TwpSCph6jWsgNKvocZLVDY7celtYOTJ+fwlDwosWMkkkSW
qqmE1Wur9ndPG9t11KXE6wU7i2yK6sx7cUsZ7sFO+zoo/kTW68fo5LRVb1HiMYAc
d9tgx7Em20/GGZrB2S1GulHAUeqrd3bMWRQBgjCUVLccJUSam8eOFKTqh/Q0dWML
8SKE6C6qk1tEAYUNSp789NN9vzVNpjr6w+eJcy23uphewh7i0aaSmUimdegRojl/
t4EZSmN+GlwEyWZ/4Y7fmlOR2D+kODVK3bp0w2w4WGebJQi+XpVW1IVW82NkkNz8
M+oxXjdEtbcK7H14bsLYKaNkK6bgSMRohFCf24C7m/8ycRJiBd2jGhokyUTI50C0
CrTcGh0gViFXIIlqdO2EOilaqF9X9RIllz8MqyT8NnGZKuQ+tQRdsrG+POFWLZfi
/e/SQ4T0rZvW4Pcnczr4Drq2Uxn83IH0b7ddrFsC+Yphqs7izU+inoWhyDPbnHPg
uG/2QZ+p5v6ZdU8Y4m0ie2OVcqVx56YquZXRmxsDEojYIUuOqilFM5vVfqyxvcko
0NF6jzgRUGleQbgzA6VU4WaIqe+/I2ItQknRW+u0VeEzKaUEBbHpKKxB7r1AVMfw
J1fDxYL8+5lrZ4g96HhMlIZU/fz4m413peWG85GAdhoV8ZX78WUX0Rh3gaY2Ro3z
fps6QkTKGHQ4ERIjTOPEaNN8DHs0eVwcvtRmBLj7VjBaYcQX5H7XOmzNVrTd2gcC
UOS0aqosvSK4IusCkhK5z5Ly2+xQ8rSbA52T68U/bAJBebw/47fSORbdWL1C+8Db
y4vUcmrhKie7jQpFL/1J5g2FZeEynhFs97LEwgeYe3orjd0Ego5vcs/nbYiRcOrq
fHNp/TOkaebNnJXeZhGTR64VvrsS8zSPyVn6aWvtSxln6wibYifZEYXl83G0nqhp
EdFz5A9itNSDZT4FI+bS3xSOMGJH7t3kHtrTt1fEy8/Gi6S6V4vmC/TubLGeYEFI
xvlH93lLuggNPBycqiPf4Fa+YOQ8Vds9Z5rB2z/dpjNJZ0uUSjL8peiCGkLE8Z1B
AAdc+TPxPc6QUah2uc6GgFH/IY66iZs/nCftG8ZEwRCn212nPyCeWe3ItJ5h2+9r
+j9ijO0mUl3nZRHpGESX/IVWXJVV23MFm1JBcs0+/GpWj1yIb6TtdyxUvjmSnwpd
C/YgCybPFiOZB/T6oPEk16gbJgo3C0T7502LJqOjoNpT8CAdZtEwtl9anm5u79mp
TWUd8k1VzuJfPaWmpp+/cWHweB8Sg25oYQArShxbtJntsnwuZ4I2v03QRdIWzZq7
QoW+cH+NwxTCjQXyJJJ8D358s0bWfCYfP041zaEIMCZ9aEpOYkaiOrouEqmJlP8T
T7uDx8QRAIax7qEHzRog/wgkoETCDO063v6bV98Pe9WaUw+AIr19agSZdljviIfi
CiwXVS6tDIL7drJe9i2VY410P6xazPzQFWEhOoqFGE3t0hi8I8MD5IzsPxflcQEV
Z1IQJNT4KU56CcRLXfMbSyxNccZxsU9Nu1MoVcmNvuhn2mPaGgHTxPRDbX+5HVDr
l9HMKR40rv/E01u0W/mndUCsVD9DE+68yVEow9ZVGJQCEBMCj8Ga3EV6ikBPAuEW
Rvi4D8r4j5B8UNUBk9f2zWs0PVC/Lt7JFIhbgNMVrOi4v0aiLOErWhDPIQdYQxgA
Riz7+XlBrVl175M/CPQMbv/lf7/4IVUJRb2Va2vw3yI5CFuQ7LLVz0OyN+CfRVDh
tza2BIV4CfUKA/7B1m8wkNDrdzZauVWCxbQ6yhkHJLUWKdx1gOwKktOXx46/Vk1w
XcsYyg18dwH6nS29OySkZbeXl6KTrJVfLUvJrfTEeKH2gvS8WwAGnbGh6dpPbSon
ie38zA6rwuFqsnGmcBswUIW/KFrUAVp3RbNRQeHUDeEenDutvI1ms5iliJdH4xxj
7GbQoB0mYQz4/0UQZYeCkhUcSOBeT3dt3rPNzBb9NnrncLxQ/125+SL7REHIUlO3
TURVxntLI3jQIw58AKkgAga/LduKXh4od7c+5UjyhQWUQ9wEKVj06gSnfWXH3ywI
dOcbyObCQZpQ+4dnd4td9ri6V+gbdgv8Q0TpL8PC9ETsSpMmUPwPnUJqWeG92fAp
HySIPpXTjBN5VeC0Pa2tHVwtbbX5jqi1CdYKjnRxBrkzux9SIphzyCtY2h2AsqEz
59mqCJi+yu1F3deMfroq6O/7+Jj+ZtpmbrQarLuHBzAAU/OOK32CEFpRqxOKlJks
i29jwYNy20RS84xdHKN/F+VoG8mC7xsjSW49HPguHjRlw8mu8jechX+K45nRgPKy
MEBb9MeU0M4ujWv4mWtkBDRX4tUkffFkr6m6+ceP0gW860jdXnSlLbGmZu4bDTj9
phHXw2UJDQ95hiHI50tpYWV/f+NfNxACozS2FS8VNwYhcPKVaXV++FlcLPdcAFlT
myOICkuY6+TCUHRYG5jmdJ8qvMMhzHENyitUJDY+NkWS/DmOrYFWChmNuGG8YYKO
nU2uUBmCqP1/OH+CsQNgJiy10oJ/HKmmpDD+DR03F6yWDqjqmelLfwlLrIRX+yJ3
T7SRbOGZV5CuEyySl6QCDxF/6VZ1TsxMqOqgzGMgojMhKST1lGkVwW835bd52huS
ObE/PSc58v1NwIH9sQkaxveWXrPPWdVppUJlILoaOl4YQQ20g8jnb1VRBr1oqhaX
OdePPI8szlI/r5Jciv2MwEtzhw6plKMrU+JfQa1dHiKGASuXg9W3ZX9pKCo4YtbP
43t2ZWIh7vz+AWqRO9JlMh1EWKIR52rVJsr9hmhhFTo6kWUkYkil1TRnoUjrLNgm
l3zyd4dgmVQgyARf8KCWih/2bhEeLuVaf6vcnkiR91MmN+UDtWvbwwUFt+LEqceW
HTSztapJJYk6vlQizzEIe7rQWse4YyGSaGozeKbRInwe0VtuKXaIep1OP7aFxW9D
xP/LY3+MUHIXvd6XSqTYPE3OSdYmZ4TZeJCy92XXdnnolCK+0HhD+oLT7h06B1sP
v880Kag9zCxydmET4EsfOUHmSFZAmMg5Is65a0NT+UYWo3Ls51zkPWWPvg4xCWfJ
fULN5zZQAXt4M/ssOkkMsKdnaFE+IpcYQQuyh+wqcWh4SbnoRzqLqY92RPdllQez
xQfO1fCCldiM97GsAUGYL1jrIO83wX/SwYAUtmR1dqTtOanoH+75JAmjCZvg6REt
w3VVIgDvgDf3YuDfKx/aksAP4JlokqJ1PfqjJVZjrtLeB5vs8WkCvLbq6+5s07kP
IxcEK0Kmzxt0u86tQtnFAs0qe5l3RINiYHyiOmD8/NE3pAoJu8nArNOnouXNwRyl
y+HjwAIntgp8yrLrS+ymZTKBXYFcaLuxAYobl2ILxUDy+WWEtFrx1Jqp9+noi3Wh
OZE61lHr7iOpJWNSX5uMch8dR0iDiWff65Nuq7F68SkccJIwM6ro8e2H2D+7baNy
MeA0iECCZa+KxzmYOGMqYX7v6Na2aIHViN5FyCeeRZ3BMH/I2vk+VYqRr9hdaCmy
LWJB3XrQu/vuM/yIZFZRXUtuqOUyiH9adEoG9enYx8LOi89YLMwjp8TYbQk5AYGP
U+yDigKwS3hZ8YpEIArenNsFzecwLJO6pZHgmZzYdaKDCLUrsWar05XFA6a5vX81
ND2bXMQcGQCn9Yhj0Ug+uixA/DCprfN/PmLypUXUfJHPpqwqruQhtQvpT3klQ1Vn
/NfUKgD93fsiWsJEo5TEY4rvnBOTDRVLNPtfm/jNK44B7kjGrlhi/9/uLxyEGlbF
5W2AQb8g9Ls8dsNKz2kmtN8LAUSkA9Tg5/2lXxx3sJsg18dbDFriSanMgYlkhOHx
d+xvteaOLN9nIQZ1SrOdeKQA/ZcB78WocKiTEmnnnA8wg30ReX1o6Yq8m3fQtMfK
Pv+o/+aUK9/O1qWsucdHT3WNrfvwzQIV51zp8YCDAd+b/cI6ezfURILW4tLI1zcn
q4wj7f7O21kqDTX//4p3r5OyiHK+xpand6E3fzTtU9lvtiGo6zvf94lBUpd5Z3lt
Lxb1N0yMfNVBPX7AlIg1diVrvBVyT4teTLHEibU3C/gEgIjtP67pQTPS964MMclM
h2wX7tb5dFdkL+4w5KBkt9hv/fFubOEx2vnbAnFtu7RkvNr+TQxo4vofxq1KGxuo
DcMoDM5z5Jt9z5+HUqNKPc0sAunuv6Q45D5xtsNlDtWiIYhv/3bvH6aE1u6clrS+
4GlnV57IUloLfCvaXr0xU4vVzm/eoaLe4O/RDDxgJaiBtoDM+6Bd6M20Ocn/z02i
los1BkNO00nOmWViRnt39zXVeeHrRshsRUsL/OVJqIwAwCbS5EaDsYdYYFxfSekU
oBhdSu1oSQ3sXkVuoDawQ4XINIFyjFtHddWAH77+jq6giivOyHtwM+Chu/6e10gf
5ChUetcZlKbdKmDlBFILJVhiNPk1O41YfUTQEU4bc414kUTM899kE9PxZBLS0tqy
QUr0Japq60yiWhe42xsrg+aFNOxKhMsDXnTdFPpGKw1JngNcLB9Hnbq1yLWEe9co
H0PzQv288nySNZQ8L0h87QegAAJqpcOR5sS98O/3Zvh97YOXabA8YDTlf4RKTwwI
ouJ5L+oaiGLBDPbH60yRy3E6xuj2H9lUzcJz2m6f7F5+DByT936XJVf09QHkysKF
kL+r+qFChefBGlnHo2+Cg1se/bNhRJB1uTNN23RSru2pF5ATmWJn7P8k+kjuZ1jE
OIeU8p/amd6vYosge3CcG2JYGYJImtZAZibTDnXRCZQmRRIGj6Df8R9ZEXaGRU75
A6VUjHFwcXR7L9rKbPmRRAs42psfbOkGt0iYA/IHdC8545qwsP3bXwB0lEzxGo87
HrROrG/ls1azVuJxUAtw0HKa3ZWOBNom3NGCGBr9S2VWl7fl4hs8I1bq5o16ovf+
imeuau3mMa9T3vdE2Qj8M5owyUCvObqyGXOWZ0TNv0Xn703Pwcr0/WbSBm13UYk6
+oggprlNjtIiPi6dDXOT+EjdndIXBA0D6gyOK7QFeaP9mOD4VOxcNDXT/ToPJQ74
uolvNiam1/bTVZuVx0utL0a0rCg1CKM6oOslnyANiZCmtaTXMA0UcwbhWZSG7iHr
/L7dgXjz0eQPy0yrNSJnam9lU7IGa7pdOKUnDHi5RzPXPcCvPBmuN0dEWIDCpYtp
QuyBQZkn17RdeKWjJoLep3QxP+0he02owZw8I9sFR1PHLzZTAw5B2dGVKpQeq2Nl
eONrDIht2cbcAcW0QmXIVcEoP5aXLCXfmmVJ0PzRWMlnKiUHwuXPxOXFPZzFK0Fe
7Uy4tsbGWUZ3LQKxdfqaLkOvDehuXDO3E9qZG5VICyu5VCsQ+vWpAIn/WZUoCOb+
hLitcmBhHiQqvFeLr8D/Eo7ouuwb+EqJ7Y7NK+/PxUG3reG0zY+7GoxTcHtmTm8d
WX+ZAebIF+mXyo82IifeIjD3y0z4lRRHoWdgQi917p0+zATgbzSI/uj5+Bmy2HHR
r4UiYRloNg4WhrIJ8QrCQLcpFQuNwevCZSZi/9NnxQYVBYSeo/BJioYXdqRqL5An
YpX/bj0bAzgKprqIIyb5WATYMvAKiPfD5gRyuP/LyqYHi1ACy+6q3BYohxZG5Xl/
25IASgB3klF3KAJSNCKnkYsLF0tMKxsYp/V8VQDKRw59PMz83HdS6xx9NP4QFUxz
1QxtNo2WgYezJvY0Hnk5uR+VTSUZXQIXv0aa6DNWmD/wRTEp8ffTSBDc+NtDzm19
e8M2G2f+RWiwPHtYwbICxmZQY9VzzbCnEtGXhMEr8Jx9P6blXbEAkQpv7uos8zE1
1WwzDVT5xtsV/WlMOP5bsYfc5TgwNyfGcG406gDJPjeUqI0PA0HECAE1tuAPEaNN
4PP3r+x0RRCIO697LEeacftr6wkJRdHODrhIpVvSEMaFu02++Jf+CGTFNuvJc2Pd
cPO86uL9ltDPmJHDZBTjOIDZrhFYSuINRszvbhC5PT/MZKzj8IE2vJSTBEJvKjLk
A0pITOft7VLE3P+gJwCxXBOynbxFYAbmGuDBEItMDNyoju094ylVEh/xKOyGX2Uc
6+zUq0346STf6py+nivd9RHT7LqDo/i/H9nst2Dq31t/f2MWpiRz1oghf7Ygedg+
At15HNADOzee3O6U0N5IAMqubJ8ku68Rwbr8fIhlmWhL0xOKzicL1L2gP5UCElfj
Z2xcM4f3UcEtpfVXQXx9zvJmK4rUuGx56WrZTFN+6L7uts6EwpmAlggxRbb9SV8v
kCh6J/OInCQr2Zgl3bOdk3pyb06o7YMHcTGSd/JPNgx05pF6gwtJ918WnbHC/jo9
FREdhux1Xifsd2FDBq0XqKUJ/3p2yJ6ZeVDQQiFIeF4wDEtYAYHZODbzCXmjvJcU
7Z4t3DiM4+jWfXG/y4FZXIG5xKjlmDB0XY17eaOi82vKhcOmq9airwyt3lOSPmKD
AYzZxgHjK2x4iCkPCWd0BCp+e3SYdHE/XkSnzedxRz3U//OSsAwvth2JELmNWRQH
8Jz8sSDqTlp/GtqpBcIkKD3XJbyeNl3UpHsdNPTIHKFK1SHg5SOSPcqDrov9B+0j
pI/Gp57Noc3oWkd4k00jp+PfEOJbndwO2vQ+xiUs5oWHfcNLKmwStQ4UxSKB8IJj
QQttfJOst5F7720xnYE681YLiuRqoqxtTYos5lxsKwmLvgulEFDZxw54b8kGpSLy
NpJEESGqn2BfwyWEqG6ceGN/SGBe1NjHWV/rATAHwqXj9MFitlpX+e2AUfuhl3bN
fAxzs4ujEEaMCUWYX6dCNwZAFcTAbfGA3XEWEtGGTUNkoYpWCYe/o+18H1lKE5yS
7njlryv8YGtJVpmcRUPevTMS5SRAhpsL0i8c3jMy6jNV9yxvfeq+AlLdeKC/ufUf
ZulNY8957JBZugqRjPd71wKqcBlAl0WGJOauLgQLyqiLuD5SoOOWeW/5Fd95w0MY
HqP5Y3lNu9eMQaMUo5mrsS1aEAI/WQb6p5gsiASYuIVymXTlhgn2dX7FGZ7woP68
8zVzr5uV89Rj07poKAHSRFUJX+oY27ZIlH8xM6RNW0ssoahp75BeHpKwu2lmHKB5
jDqRBe1IqJQFrxpAPvHQu3+QRoJJwEn1jQBNEcqZonUL00lEno/FornggpBKZX9k
Nk2j03fiLB4NwJVNZTzV3YzEe/FXDAjasigQZRACr0lLNOnDyeLaYodsDyVY+2IX
26opSePBqIkp62hN0Ym5qepaGsWFVokPCEzeDu3LJDfiBXryt6+RqnK0wsQ3Qmsf
g7Qu/o/B6TEtOOYI1eRGDT3QateRcgmsCKgHt0djKADjG1BrowWjocPFcAdCiir+
FgsoJiS+sqgMffpzy2sgS8f3KKEoYYiXjmYs4Hj5BOPQd2vYqd0DLmI0afp8AXI7
FfjQ01gIvn9nA/IXcbInLVZt/1w7X3Sre6wYkadCvFCvTJNdL7jLZ0c0A7tLD/zI
BHefnaUpDhE+zpXvBm63QpgUDlZhbUP1m2aku1GAis64gsogTYTUdF2VJz3rTAL5
NDe0Gatw/qSX7WyPz6/GLcoEtVkTtnGV4+BMxQnR5ej0aG7CWtCGkA1lvtGrcUQY
+YQU9ZIJZQawP+G6USvSUveWP3eJXf9xJ7RQYdAyuR9yQNyK/+SE0PKoGbrJtU1Y
7MVsXMQNNRpKanBRR4Tfh+JqMPr/abLyuGqFoBZZKk5IQeo1eiEpG8EeXwUHI5i6
lq9aSmx4RN70tus2naiVTz8G866C3fj/Qst4ToVXSBIRhsXdiMaViw8/cbdtNVMt
CdYxrPClpaHt6OYS/2byap9DI4ur84GT1FMv0dCvC0CzagcrimRtlbp8pwybR/OC
eqK7dTkEogjlWm+ZteJORwu/0AWTzMdb/+2da743JpZK8qlfl8/5g4vQMuGJUM3H
J8Eq0fPEMT5oCuG5TBZz+j/cldG4kNXJ5XlPesIKvcjpfral0AM3CH/QL0UPHvro
k2Squa635UdwTtlOI0n05PL4NET7i3hCCEq033RrSpLdSd1M5M5rKhNgZS1rK3Td
v9N1245hwQe9DOO8FzoHV2hqngGb4CUZ0B9j1Y2UWo+BxqsUMdqNVjMcLkuoiXM9
asjmiD/ZsjWtAHTlU7O/7Ik4ANkqLoOXUCKMpwub3AXPiDn4YAsqHCM+PDk9ThxC
LroiINaPskMg/NGdSNCmO+Cb2YEpFCtc51REq6cKu6kW64LXPO8gyzuOILXHumbk
SOUYC/mkEc6f4o/yRu9p+O+aD7ouLBPWi1F/I3HlM1rjInWg4Z3+WQlAlh1fJ8SY
9Tk6I1YG3wMrZp0VG/5vPg493bAmksNF9QB9EaSsgN6XbkeNgucsDyGsD1wvKTrK
q89tsfv1igYzLcJuAnVd7/mWnmE1RpChoiqI3q20N/O8Isb8+oH3cwgQJPvIbldp
EVnnWnr7r7Ci9aAKbFgBU5p86cMM1Htn3nqzpMIgq7otjQFjncq+RggaNCdmHpOx
8sHK3ZY588qNZykA6x9pP7dbeHzkAr8kWE/cIMhpRdXHWVuqjwF+1R7x17boNghp
ln9J07SrnTxdnHIbKLULbLEczhlmyiETvOFVvi9pSGW90Xiug6b9QKwc3+JZr00y
uYnmg0w7Q0/I6ljuHLxO7g7hM278e4Sbnd8IRKcNvdCBx5Fv+0lJ8S40L1sIz0CH
FzDCZb8Ph94rA/7NdSJxDdD4jZfldDJ4Pf6OewywELxCfqO602zR9jbwUpfO9qde
r6NUndDk6d3J1wPKEhaRuX+7DgtsvLiOgnxP62M8cWZNieWmpL36JzWKgcrVu26s
F60LFlaVYSYi3uzNoNbO8t7GoJwj5TbDOagEA8/VSzMCSfGZfPzjofXuJ67Vt1D5
OUFAtUzWLd3yBLNVrXuvOGaqwQRwF82ZFbfG8ItB2fWQGO/7IVWIJMHuvBK/iyOn
6zqRukfggQMfg9m2PQZjuZE2ifNdE7r7pixVf2Sv8y+g7S/foyHqaRgt+H4W4x9F
RrdnAEc/POvEoN4hKl64x4F0DPub6jYg+Ru9VIBDNQigpQ7JCR5UkFo3vfddaK6N
9/AU2aTuXr2jeaRRd0u8y2tuBD44VDZVaPFAY2val6wiz+fl6qe6ik2fIwhYjca3
JtFr6N0xchAcYBGRAag30rNJchFZ1HvX5W/tq7w8Il01iIhtSQuWP01CutgSnr94
tqGwv22iltHq6FnXAB56R+H9HDNFSiYoWNgfjECPFbxC+1v5IfOsZPXKEhDwGELw
A+XICAcn8y8HOnyKgDD+MUOaCSFxD51wCBTaN41BFxg19hVDYkq5NorbDvO/4xBi
rukQD6m1ulMRG7C2VYkL0O++vS5RHUmcQlB+W0i2JDOqV1EXuw7K7wMXBEM58c73
zh5SKB9xj03kgSdPu0cxwb1nJNRC4I7w9t7V13hqEOrI9vIKnGEfdnT4EshINdIo
+XvPe+BejF5YSwSQtA0vk0o+EB7qbmkPRfJidsRlZbvEawQcATw/N4k0yuP9B/n2
zpYfDfGWslSyTDTXcBrd3bkUfU3Xs5PuC3fjQm/3/YQPc9N7x5dBt334p9FgVNZw
Ah2D2fZ5lc4YJ8irVM5DJp5/M5mmvQf83aMdIgKnQ/9Dv0ZmLVpOppIj7iEQGV/7
Cq310XjuaIxkUCC+FeX9ZT4v+QJG0kUIYuuezKEW4tVkX1Wn00NjqdadhbkwFD65
0An/HP/SA1o0TikYdRNfbPfChdznDf4QrKycItAG1vhjRDGiQiBSf1JxgsMfSeFf
PXvQF7GP9BWnBk8pvYn+sRblWvHHqDonSg0/RfukDhtxO//Z04S3Ds7bdJwi1Kqe
2bCm5QSQFrGK8lc/W3XI42Nl5MZ5Yhw03I3/VbsBwZ40DDJPtAIaaoA+inPeWj2H
vc5+6bCYgZjFEmUTqUIIvfy+t+GDRDEzBl6V90+Eg8C91lW5LM5YKDlbR6qt+dRo
UzY6bszGgT4xju3H0vTFlB5iobOZjh0HeesADSkLpb1cz17Pa0Wh90LWpGRy1dQH
qw+0xjhN7HwTWBR2njUVMmFYccPHmqifGnh4dwXk5YbogV3UCk8NjC0zIqJVVgpF
MgCM60Q/uR+Df5ugJ66wMtgWLW/BuLN66ijy6cDWmY7bGnTjOdkuUVvis3UmP76H
Bsyqg33Vlt2loojgceWOxPPb+UQ3H/uzRfCNgCSDSx/wewDDJICRIbXIFEz//TXA
hqTQEii3RGpd2tCFMt7F2NLYM3dKuezoQfGQVNlLlLZ6DaxchCoTboZWRooSUYR/
IiSzDfiOuBX/xb6bYhLIvZrwNkpdrUgSW0ZKQ0eVFVgdh0QkvHEEoAh0ylDuqQ+5
kcM6x4yhZmR+HPdiuvmbnEnhyKnBf6Ogt8tOty74jYigsET7dSrW7zp2DeWVeNP4
lwx+btRMj8tThqXtNFSOWGkjVm0c2W3uJDTA3o5JmTZRKNEJdSogwdeT1oyJsLcc
/1OWd92oy0eSyaAbL4EjAesik0z2RXfjdsKEcSdyWYR9YnIqAG3Q5FDJ4Qr1yfiJ
GTWelTlG4UCTmoUsFwZdZm49uDBn4XE7E1LhQzHW+AiZakrzoFC+krRugzTi/6vt
y/rV8IyDM0vYB/jIfpAM+YFyeSse7I/27rIFmOFE2WtC86Hb52GfUTvTFLmwUg0J
DyUbSI4SAEXfX/O33ZGsFCP/Y0Iv5X2Q3UyJexHcHuGq3VSY75nN5QAW3xjblD0d
VzoYKyw5O02HQ08LLScQS/zT4RzwfigPDWhcSTlEjfHBJPLFE/9rCyEdD7wehbNY
6WC8x1i2ekQ62iGV9ZBruXJnGztBHVDqpdNXjdb0leozfkfbjJ1rhPAearN0WgsA
HxOCiv4I8/xGYPyzFE577mbgE1e7CWDPmdcPWMG6HAXr52aPGn3CmJAlpbsn9IOu
fO3r/DY71T3mldHQXwXSIv3fnaGWSlYuxMwVppcgO/xyhE13qfyOoCUcrrF1pfPX
PA2USCop2gTjDlooVyRIKLJXx1sLK9QW65hersTNvzofcU7ZDd8XbrjMN98FcHbs
l0MN1JQKtDdhcC1s36jC8dVxNJx+KutRmmbVSPdd8vyfZKA5keVm+Thp1KP0oPIn
ll5ewLh6zm5pr08sQ1c3MR1YGu02c402pq4ynyz5g1zAVCt1GoD6ijMCUXZLLmyg
gTCNkJ6JmCfSBYzCtasKvUGKV5lxw7BTYP7oMLD9uOFH8vFQDgQkZVpF8O3+c56A
FCCnMMmrse6vc7zyUcrzRfZT59bNM4UONb/ajxiTbVaYV3WM2J2a32f3x33WnPr9
F9abr4ClFMe8al3pEhdP8QLaLEPG1wgm1uLeFZXLGVnqr3xN0kQQDN+SIiKvlC9R
coszoKLFjEkwE5HYeJq0bQ5JHJ8/6lnujiO3ucquj2y2w+j9aG0JoNqrI1TBhGF/
yIWaHl9x4OsCIFN/vTngxUBHV4/upbGUjadshEffgioBe96mrj+ClmRoKliDKQop
g2hJ1YpaIKmyCKhSGB6BP6ONwIXw5aAubYxMGN9I4IIWNL5ToAA4kbtHjSgKP4C/
8a9BQnmlVrcCB7oV2/3koJ4kKGvtAIzDZuk5o8XseO8mL2iGUJSdoRLEvyGBqv1U
/OOYN/yd90xLGvUoTvO/1hbMROJORHHLJ1UjjbMRdBXYennuXYsis8HxNSZXrsGM
OlYw9L8Dzvbs71Mom2maa/CSMOtk+K3bfCm6CnJlhSRi5OD2KvbuhV1iT6zb4x1I
5vVOMhqxR6rBziOzsInSR9N06IO73H6X5aFIJe3XrkUJ9Goob7amCM3mUFEQepXN
iIjwk4tPI1rJ3VrAWX/7MhroUX79REFigF0gOxYeGJ23b5D/FlxCDUFY+7uf+M15
BtxWuOm1nSuvZHbE2lgPFGNdHpNuPgeiScx6jpHla9La52HxEc8GbYJpgClCm6C3
t9a6JnXIsFKUOzfQIz1fdShpBMRuUFiiFZNIwhb28IjnapP7BIP2c6NHrIw75tbL
vlTU4A0hdbakGntcKIXZrp/+ji8D6BMcpDRlLFByXwybgbWOTs96S4IcVifkdaMA
zznJ0VUvTcOyiu9aoajsvq1PNoP1bNC5YSTcoXaz/5SAi6f2uH031NKC50r/fLHZ
9NMAJ06/ptDQTzGEfRbr1GtuP/jkoiRZM/77L5zfhM2ov4Efp/ZzshxMcspzXTXa
eYEsNOfDlLUPP5nUUg4+fwgxw3IrA5f1oZmzBsDziaLCzbK9o+YGAwnkCCqUMxnp
oNv8QUlHP9DhgIGOxWnmH3E4tZBaKGmLKWZdE1shwGIP3RlACA8pFmXNKSSaqmns
En/6LIlIT7FXF9QayAI7VG3WAmSDJjIMNYAuOZDffcNqQpXfKZao0JP3KsXwTO0W
DDGSDd/6uZi5+wzHXrxU/9Yt/f9tnkqsgZpoIOzX2eqKEf/xGMtUMUkUH97U7Ma5
VzPq7IwsLwZ5l13E0Fnw4bksmlwOvC4+3N6qvNAaKaeSPeGhRNi0++SY1nT3li8q
FpLEYtiiYz1/39xYUgL3OPNuMKM9D3MVL04zfzmVqccLuD9lLyk1acEDJTCTZ99y
mHZBvSxmVhFaCw1zaGTdQYp88k9Xzjb9kWb2bkGjFwqVFdSgJr7s9JyxHCTmSKm4
NoSJeaWE63+SA2u10nwFkS+se2PTiUI7367/rKSKtIJ8qpsp5UaHHWHeKP4leiMY
3DAbECSOOxNVNdh/6NldZHiKHGSlGa+mn7ulAp/pf7m1ysPTctDoDCLKt/Qmh36C
DJMRA65ACOrDNJsSMlzkdI973g29/Z5ohODSE1muSklIOlq+hLGHtOjTDx8PhqXw
u7SVYmyZMF9FxCHLfJo9sa7J5z6iuHZNPDD1612poC7lj0rv28aihJEKKs33OLIG
9o7R+r8ET43pbzBCfELldR8RvjyAEmsK3JDlkvjvFEOlMFJ8B5CJXtAFNskTdAe0
5pldzw3ECqQFT8mRf5vdnKi96lSHJhqpha+NIsdZjCjp0dO4mCANwuBWVOJtJqqK
YmcTkjgo2z3kB4eZdJ4ZAxW1NtnfVcQnt6HNxmtXtocI+X20rRTp6uOCNI0I2dZ5
T/IunSw910h2QgLUrf1DIF//KD7Zh5TeO4zw0KpAb+ufC5jG7rcQBqZLUVjRCQMD
hTMsLQzwFQHA9DS7CxhOfC4RQseHlbNPRPmEJjZo95Enmdc6Zhfk5v9icJwU9mrQ
552P3EcgQOuh0PnkZsptklhVXTzKzeHppOaneazK/H6HQa+qZpgPdRAXR8LtrbJn
VbnjYJzo1qc9lwJSgMlXE0vzHwvrJ30h96YB4DvL0+nV0SQCbryHca4MvlkIU/6X
OkWVXYOAf7jKTbjXtG/vcggaK7TfAFQ7Bmp2LpwZ/4xLro+iXLX+oXWZNoBqdWcz
DL57TdY0qWy7alumvjajicqmeEw0DhBq1tMKlkKBD9gyt9vuRVXHlMpVq6PPopPK
q+Vb5wB1jlLuvVF2qP7Yt4MIwp/4gz6pu2aHzsm/QwE2ht2PwyFexK61FpD76ATo
SOf++Vtv6rvemTjLoFiJKbU6MiBz5JSl3W/s4UaxJpIWIEX0BpMDUd0MoZSQ13go
V1+cE6KwjobdITaRHhxEFD5kEL39gXP1HBG4afIZo2IipNw9NgBlZ9cg2c2y5j3T
QhJOCYdCpEL+pSHXRfznn2dqt4kLm3eqiQHcFVi2cRn1wV0KI0S7c00pSYYzGe2U
IiqizbG1r+DcmB+ZPZauamF5c4EDRWOiJFOetNU+jYXs+uXsmwmjZiGQYGIM+ubD
QF6zDduQccuTLppuX6dDWJjf7rXGF4VYqqP20bMwuwbazRiUGKqSu3J9hvgqtYB/
3Hn5i/1O1rywFUJ7dG5gSIz/HErKInGTgf5yWlEWvSAhOBCDnHfdDtPFC+VwTulr
NPCwRUlfDp+7bLVENsnkNIFC6i26bSOFTZbrKfb2MxDygJipM694UPlIBrrsad6z
EU20zgJoYX4rqsMTWKCcnm5HgmCrM5EEWtOHC3ZCZpUcWayl1I278Rc7beyvl7/k
bhdokBP4B1GJaJgkQXMEQ8rJTpRBCU6kZzJ9NWdv+7GHDCrQ9g/EGoIZp17dGWRK
oyIYZpOTcx6Q2UamLL7/PJn67uMPkqLNbQuDz+zvTVfx5XwVguj3b0x7/teWiRGq
xXnFGDWGnTzUbhTj37GXNB1IVqse7Ca+6RM/3PNho+hdyRzlpsnOnxm7ZR9i6NXV
IhvAuO8Gae/BK1VNmHC3hHoYdgK5WpSVsYoHxeqCNjrOaWtH4sWL0k8CljeA49VM
kbtrKWVLiBhMByMSUrOiYK3IkHOiu4+AwDG2weH0bdN7VYxC+aCKNpzDyLvLqPuO
RBeVFVKiPZZX3+nUhkqBWEbhCVE1lJvkd/sWj+FFc+1l1YVzQsOTU8LE5ywITRoc
YUzWebMuU+jawsA9UfAvMkfjGHGDkHZYv26kmw6n5vC9YJYIQiQAPajeT4Az7apy
G7YZXr0AphoXRyBPvsVjpmatTOFngGvI9QiKx265cncIGT+udrDPIv01bET5UBXI
lw3hjRVuX/h8f3wST1bdrnn8HZStL3DRVQbSGbdRAJwIn/wLmc6qNGuLZGbJ9imq
big6/gD406C5KepZpVDfiu18iBbixwsFvNXlUjsRbJa+cd56kTjEyX3izk0yarJt
L6kHXRyZSPt4TUIw0AtLbuL6prwlByfgtILJMNm0YrZ77cZGAmBYcsazfeIj345S
PUej8hE3QnEAP8KI9U9FolxZi6Rgdm3521nW05CKHcZFQMpvW6ppRIB8jT9ligsr
EJGAxjWKkYqimhIQoIz75su+/ffMkxYETVHgdnE7p7n6BAqrYOVl+EvxHIXhwThL
GNtIrYG0gUhIKvayHTm6a4FTv87o0P29Y27P4NkhUa2KAI84fRdGYWOhaxd6gXP9
W5XYXF+rxFu+CUpVjDesPfHVlLo0G53lsO7HHhxz6z2ozmJTsqeRNW2aW7CUEBLP
DelbsElP5thfI2pYsavjVZM9sjPe/sXY8Z0PRJIq14cDzbG3I4w27cBfYV3QigEQ
XwCr0TPOEXbw3uCg0Yl44A8PtziaDzJzhQTF+13uS8AuRm2eWmfGKiQaLlxQcfl8
Ire4TUOagoLoA5ubKo158GCYBCxrsRRCPrhO6B8Hc4FEpe9gmcvahXJbcxG07Wwm
RbyCHpzvP/wtxmSm9QGLsFVWZMo93dtnAOs44nDGzUWzsjOnXLTxLDO7ZjL5yhsC
C6H3RgTeV3JeqB9eVKrKCeGPmDrZR7/Lt/ClJiwsVvL+GYIJ7eiF3/+dHmP/nXxS
piFlbnyPQswOjTlkLKC4e8m5xxiUjcH1djmXKvKutscXFMYi1t6UwuTKttQ5p3iA
Q3jwI0wQTG7+kxfRIVA1NJAMPXAVnLEQ6bCa87Dq7wom0be60BWDBOs+hNYWWsUF
U5u3SYw0jLdigc5wplx4USPCKzoeznqTKeBbkv8HmGnfrHFHMm5zAaDJa1WKlGom
SWb4GX/O3PXmApigXkBFyqetYo58GHhNQPyclDaw+uP4z+T2LHg40taaLJCTMTTJ
+iWtcXAfhXuXTfo1eXdX6AwEDAVWmPYp7svLEtsnZHdTiPaA8DZVrjcfWke8uuI5
7ldPaLmm+qpysC3N+I6AQddgcSJDq4NlkTYPaU/DB2qmnUmpkRmFbcrHAZl7KAvR
GhMkR+F33keUUR9OIttvGqOTpTiz0Enbs+fLWZQ6h3ckxo41hXpf3yvXANR32ou7
EUPvHHlbofzfHg3loUrJpChOeHnP0B7cVfBVs61CHbHQsGQ/JtIl9hTxRCLcltmK
WEhNNrqGlZ53KmezS9FnEEICWl06NTFpiBzBlC7UNS7psWAaACznjDpC+Ay05uxk
SpSQk7wxAXy7t80vQkuS1X02/opAo1GxL8lYXz0Klh3nvEJfquRNg/yvnwNRSn0V
3ZAHKoanpWZTo0ZBvdz/KKn0cn58OguJVNtX0GX+8CgJjb3nYSOOOGSn4zJO5R2b
JnKB+1R6/UZ3nSCqfbT0can90ggsLbCl2G8a4nLywxMRFKAcxGDOp0hhVMbCIrum
3VygKxt+XIdWLf5W9IYSKYw4nfXtIT33oQGS55cdfL/MhZjyOZGb9MEmEMyqj8PR
bQTtrQseGWQqihiSAudno99bbChdbgSToCmq2zpKiyZom7UntfH7HWVlH0Q1R7da
8iNa/3PyzhB68YVdPgoBH6E2L7d8RkfPPOq48gphfsxSNUwTj0H6aahiIQW6wfxV
B/CHlbczAbfqJNAAy8zjmfC5awP8/ViKKNkcO+lOHJtPJUFakXkS/zgBE8Q1lhQX
UG23azidrRh9k2JaINKRDcmdNS/EvrZqRargoXiXciv07kn8HPFsebQeIHbSvaAT
0T4Tw5f4bB4NOlGhESkTHEvPXJoBoYT4L1qyBAMjKzVPMnusBrQttDklTQFHm9Il
SPY6IvmOH26KdBzfxbTVjffac633n+U11L0vnZvjop9IUW/HUA2IU16Iy/ynkx6I
19KcRepWq0P8fmllZxf70mejP3yeH9D+kKNdgJLylrTyyX3dL2gT6L6FD9nBhEs3
CKkoNxxafcDswwdzwkW+gvBwhL+qQVcLM3kyvI7HsvPjSWaWcVSXG62KSq4Cfapz
SaHa0P391PV52qiWZd5eMqXJkPE2sAfNOQYyxzY94wYulq9PKDLXF7oCLcTFwEhH
w1INjn9KP7FRFe5HeHMRFL5B41e4w/fMsAcDv0yle1qLpHEbVLQbpf5ES5to/TmX
N5rIVqyNWHF1u5/CQAogr6HWVrhcMPWJJfSkqqp53XD5g6Ck6jfPe5Wi6lZC1YxI
sfX5uaPGOo5ph30Tjc6LTOLTYn25P7IJyGLP3qpijzJ4ihqAeGDc7X0pzg8C/cxN
6obW+QpdwC1ufBzdK4/u95vMHvg9QUfG/DZhkDw8MAceJ7hs5WXUd7ycemj4WoAP
w8cwoSzVWjcYca/ky+M7omYOWh1Avw0CSVDnRo6SzXc4DwfA6miH/EGe22JhiMHN
Yu1uMgFMEiinXU35bolwEy89myDNyao4p6bXCPF+5xHqR3KdN3G3ssd9BiqWtiV6
Pk8YwCPXCymf7Tklb5tAW1D8HjkHy7koFjv3dh3MZWefP10P/eb2c2p9sdrsN738
Xok+t5Lkt6J2s1txLtWkFPuCFBAolDGI884h6lHtHBAAN9WJuj7xQCW9LrBfl0Sq
3FEawdHV700AVfphnwoHT8tS4tJgq930D0pHaTFZ5FfUeAI6iBausK767DGnb1A0
3eiRtxZaQ9uo5aGNLyLlnk20il++gR0HpDnxO9bpMy5YBQIYNqik5J1R4z1v5h8O
+4sJh6DEq5WHMpx2eNljYcyb9ENfzaEcLOv+a/rma0dEDOf7/pEkILTB6OSG2mbV
NL3D+bYoFBqpvEfdq4Gz/sF+HgN9OemvmFjMjxNHiQ+Mhky45yieJXYYTO72SxtI
Ghn0hUObH7aKYyr8zC5LjKElHbH0VhcwKR8BvnksKdHVGtZWCkUdFBwvsOJYReio
AKsPZXIgyibVbL9Md02r/QGjMXkfdvv1KT1u3E39ESazYRxibMENHgs/eXaybqbU
weKVk8Lsc3LrdVvFYtVeURZxvoFA8mIp9CSWuQjFTv3HyW+LcmLaKbcUWCN9BLKS
x04lOGYBF67oS5WQ6ftbhsRy/zkvercE6d51O5moPjcnUKHNHl/FC4V1SMRWJq5h
o98+d4/CmPOb8Sy4s3qoFJUp9v3m0y80/RX+aoGSCRWV67Sh9P66Ui0h7ZyK16Ec
cjMHBzNHe7wMd4ugmsmDoB00eMzkufn08tNqxKjwchAaX8UoLC6iY3So+aUIQApQ
r+6eT0emFC08CC/mTlhpsUD+/hLw7P7bniv2H63iBfK7xAXnkliq8BOmEGLxH1pq
ZYsDJugLnibAru858J0U1fHodxsBhDPjMeeOESF0KAtf5tgV8TOd0p8atyr0gTYz
6aidehU/EtZPekXXHJy/O7iI9uDD6/WHU6DC4GKO1XrWr/FjG/f2gPNvMeRLUjE/
BOpERyAco0jTvZnIAPhWLT+B8efiZzKQwMpM7PfBE9Vnpwj5RumAQT4Eri1Pece+
N5qtyZk+HZQm5lMqMN0jqwNVmqCkMeRnOWamy7a71JtryD9iSjiqaVbQsU/r8sxf
mkxqtwGMkTcyalvs+JlNeaHS41KXsbokYOjGeXL7PfFYWuvH8c3tnfcW7R+CTCRf
c2H7k3jFFJvfO05NGaf4TkiZRrs2M8inicg3JD3FZgVQMZV703Xm4R0xgtszzV02
dmhF9Sa9Mgt0E+mjP+N8bPBilXs85z5IItqI+wprqiSlpBZv1NiDZg+tAR1TQfWk
BFznc8fLAXspFjXUwUtmTrCeQXLKcBfxlCF149TPcK//fK6wWY5QXA2azxFi5hw1
MZfKUlZkXyOSozS54wQ6KiQDj31WjvrZyUuSei/4DZeMrRQDEum81OstgUHc/kG/
/aw1ot/9bRvUIDHmro8N3qDDthm9O8XeLS5UsPK1vepmSjSZwGoBFn+aidOg5sNO
PO8+j1wvLK2RaavJOCu/M/1qHs/5W3mpOfgNVQ+Y2p1g1Q9j0I1JZ9VcCbZcZtzc
NJwZ98waxUffLPu9KvuKcgZclOcantjXHhE27uEKCOC9OiDJQNowVUPdCyku1TWU
mhkFEZyZSQUaZM/45rEnfuQXo+IyAI61hWpuysbHemFL0QPvyO5P/sO44G+MSDLU
siMjqvWzwU9mv5A5VKuNv2zDo4AvAfK2N0Z+f/NZPZwe4BJveavYRsaW2BvqCNht
jeaZgMv+wN9VH05ULoUz0xm7vz38lX9ZYTkp0i51FYqLYco2NaFNkEqRsWoYUJy6
WppKbTgj8isxwAWUYTwSIlnfRVhR6uEtJOjQTd6zKBGELuGdxRGJ9B4BlgMwED0m
d5WG1yvfRoWXAmGUw107IJtWiROmrYT7DzD91eQGy//ci9apzeNv57nvRilDjUmC
E0QHWQnrGg65aHSsxawk6S80JSQlxiptHsmNIFUZ16MnHudAiaVuywB4nXRK/7kY
YoABj2EHgI5z7xPVO4LH3UrXeyl4vmTx1mFWxEaTK0/PaZfZVApxh1o55V/gujs6
neipPyvkjw8QsdTHfBbzy6fEgKfHO1NOkoKIcHf3vvwjM5ilh95VaLJU+aekukgN
BJlVJLEEvX+ZXuddYys15SCN/lBSGCk0P3jrk60fmxVzcCAgxmBa50BrykY1MQtN
IYi90imYdAhXcZ1zmY7nKsRwNdj57GzHqX8RV/2AKVBSSvd1gsXKxh2J3dLNrGr+
cGYZzEkm3HMcBokfVbC9Ih+ve+xomFiMI+dg93c7mYZ6HKGy+iwmE+tcKc4tFq4w
+wvEUmMZwrc2xqWkwQmGjH/ExGNuncjrBROcoydh4lftt4B7YkPS4tGCll8VPw1L
1JvrBcjWgpvc/ftayW6M68157h2Fh5qnKSKsNma/rebYVxDMFx0hbbK+Dk0DFrFY
TtbGHB1BD2jRQF+9FGQe66MLPc/r6ESC2lAOx0bIZMy3tWWj5tFWu+heXcg0mn5h
jtWjMsDpEbwcFro3TYqmLlDgf1/IphEZZKgYnuDFRszGGUEI2ZdT28BJCKuaxjy2
XR73fxAVAqAYxM8q1NsFlyCWYCUVOJrMXpr353+ZDDRzPbecTkivBAJT4sq5WlRf
VI9oV9td9C/MuMDc9JXy+A3knacahtOS8RjNle8jibz1FfCJVmOHH6DdlQKdeB1F
P9e5EVcJEx5YECLKy2XrXQNPntlQEtBqEk1hcQ65yWJ+FVpaaeaal0dkcVnBysM3
/OtNe+sWmSK2Sxj435w2F2yhHwnr3QiJgKelpiw20PZOrMl7/qcBHApRPL3L0aVO
zbNU0DNsrPvgHSqhubdp97S8mxBRtBY9fmzMVT6ZfaTskBtAEdlJro1JdKycJiFy
olp5U6f2LoDb16Oa4gjdXYhT4L3zG2xoi/85ui4KdaAUzd5/A3k6XAHcxKMQpkGT
jLaFd9/4b0rkNoGR7/V6PfME5gZJ8megI3V7v9kVQsvDAvOWCIngYb0V4lWj7ppq
XSc+BXqhgQuheZjMCDsUWRVDvM2pstOLyh4CmZnB9E642QFC0Yh4mCs3dncQHNgm
cCcXwTNyZ6loNotLXNh931FjsgNi/YBcE7bWgjfwYhV25xzQgD4OM1r2QBos+KD+
3y+nHWnTj97/x3zI8lHPuexdLZ4Xc6uePc9BZElZUaTsBVFSGeADPajCI1ntPqNH
vDZvWRVTspz0iAKK8FucqkBExgAls41wyHzhtXymPl7r/ue7hzLXtkIGKoCrNzNZ
XetXtXglwNCA2/X5m6fnwhRrWANYadTfz03OBENOWaJCtB5ZwFoQyxzawafz2Pmm
UUDZIvHlRKpGo3wMu3AB7h2p8FOOwPZSKzWKECdnv/2aHRcxGri//49cRg4zEURT
9k3lGC3d+CqB7O7rf08q7Nwd9jVXMXnjcMyUbPWOrO8Sg2VuGiN4w16R7pT/oNHT
1ETWRKuersJMiLaCRbbPUHAe48M5gD3UtgL1NNChbrnxJu7/OKmY3nMDBQyBnt9p
56f4fcYpIly/ybft9LLpEKxqvtIw3oG4mjBjaKuZOU5w2d5tg5F14pHdit73E4Gd
K7kLxU9gxxQerocgYBZISPEAHl+rjf7Ms4U5Qr34efjjXfx/wzfALhr1PiJMZYoj
QxDRn7ZyBM1gAkh01ybr1SOaI7upn4ATZfkIO50hpp9ccU4+Nk7PI7cD+3dpukku
nVtHew1cnyAU4thfwfU+ova8KXlwXZF1/rCTt9DhaRmmHgwgVSz9SyLcrGbWSQse
8IJvh8aZiNoTkk1zHYt0rypOcw9tUavZyleHq9Np8WMyyMdcdDBx/LDd3ZIlw8ze
yEJKeCWrr6dKkehKjwmqNLeG/XMLj1xDoIv/KiSYthguK1gmq+8slqazFvN3jHkV
E1OGu3drGCB5Mrihe4HpAlgUtn4qxJilvj0WPuYn1yik9/nEphqCBVNz7iZbFgBz
iWGZa2QmTpElintNwi1hEVyPZJmHIRCaFmWYEdfP1XL1yBax94NTMaNnAqzDUwAS
hjtTcrB4CQE6dGP9eCFsoi5JkvZr9qbmA/Q51ljcBudKQ7Ca+8UuOEUVzWCNzVTj
sn6uu1ZlSoQqF0ifmkeEsA/NQiL+1lCU9y1E6ldyBcigdiQ0v9+O7VEjNlfb1lmN
RxHe8IA09NjcIBKiZVaBDYbusyD6F/olWqDcE1EEnAWC5fnjk3w/z+EvvOTXcC67
rFpNbzfe59dDJGGeuST8OgtiMOAaoORxcpCmB4N4XnHvWodgBDOkpIweADC0tcbl
iiQHNoahuEZQ3S/YBpWSznrt+AZRlxjzatHsZsto5VaFbiGHKdmEIS+37/gWVc+g
pqqB+BZ2eJY+xDKiRdXIA2224LthkLrigmLlqgcywCKkCfsMPtgZNMdXOCcs/aSW
72irpZwJYYgbdTqbRK+8y/AdQurdzIcBWdr6bZkv34QfIB24+bYT4qo3D9KP1wCC
PbsZYAqvIGbvbXtJtuAPDh8X/VPnbVcPTr0I+cSn1LETYtpcZOPps/TXc0K9wIrm
DPFWQf2/45t1PuuwqblId3WJULnlAaJ1hltvntTMzyDHUbbS8jAED1F4No9t3dc6
40VoBpiiHVBk3XJtLQ4WCJUMJo9n8+RDiN8VLJC8lYtvxqfsKH+iAKX6zuzAP85X
bTH9eNgZgcVY2P/HdIdn5yK00NfzRbx/gDcdzxOt3SneHo5qDiAsbWSWjcOK06yu
oZtQvWlYYR6ZPC4Ky/+W7gWXQ9hGscwVuGIIKbbOUev7iGlS5sqjWDKekMomhpoe
2TqS2sqEE5aMD5Zz7sOJ7h1PScmLs4RBECG9psmjpT8TPb4Ze/h4gUol/UA6Lhqr
yW0fAq5LyXP7oKkrqzTnOW06u+KVMVz9g4f/xWRIpQUsgm/+Z5clzug5v4TUzMMs
2x/uiHCAHA9JPpBwffIMf2ci32CJ9sNyKDITUkxpCZwl9RYiSxr1hx7Xq1ib4FHx
oAgE2+SmuPb+5zCJwybSJBuB01aMxtWBVHn9VJJFWUWrsOQDNGwUJYhYAG9ALYD1
PB5xhy/QBQr3pB2jUjo0PuDbkDhKHuyswUJ5yRpksDnlRlbouxQp3Tz4ip3cBT24
NwPSJ5yz0QOJNETr2wacjhycy3zKSlYxNtbkNiwXcC63zqV0cFNhSDZWpnkE6eJr
Dd7s4t6fWObzKLIsRwRvwxgUUbxf2XwxTdnXxbtndy5BEs5YnTrEEDW2W4z/bc7e
HZJrhoD4T0AwfZYuCAEcxmL4gzBcjauYoMaZ4eendkdpTdi4enqPmKziWTbvlvsJ
mOUpYTbUG/pKASPB3vMjBejWG7wZHyn/D7GiNYCaGu0ie7UEb7TD2reMZ/eQQ5o5
8DYQbi+/FdaZpNVzLccV7G921Ydxilt4hqI8cASKq6+cMx6t8j92GO9l+2uiSAD1
yccnzpNS1zNRzbqgFuvNV6zGrJMxsRa/tuX4XPTKCrP3Q5s+AsJaYbfkSQjnHtVl
7yBIXvlpUivQ4BOrUzo2bRzq7Gt+cPEZ5/MZDV8C0NsdAUqWGBmOFAW/uZ5/2BUM
3Jet/GKGaonAQAdprAXwDwDr+eFuIaiJ9uzN8U6G9eJgG2kPc/ShNNJMvTb/CPNS
3PkEjT8oYlHG5ymf3M9W5FMEUf2l7owTbAKzrZNw1Wm94sXUVupB8pIYMsILjV6j
TyngqpFNyh8k5e245wSxZRzHS2upAjeEIVu+dLkyBiSD3RkpWqkdLQjHt6cz+QVB
CjCBakF77aio2mMdNG3k+KpiVVHLG8nzALBnh2SnKgTpV5k2Ol7r3Dt7IavBB5ga
sLDb8+AKoyeuT1x4bHqCQol4Udmfn3hrgbGjmlNQLs6eW2dkasWMHhQ4qWItwgnq
sfMuR4aBhE0SSjpiUAk4xSzpTWd8EqZea+MSnuCGNZVPBPLbszUWICwG/3JMtqYz
qGSydv1goYQ5PJlnsc1MYxGFoq0t1LwViwieydAUTemWmMQuAytJoLpcEjHS00G4
2unT/lspOCFpSqZepewaB3bQF7aBifxNfV16/MNAibUmUshbrzwpb/3o3W6+d8NY
leQii6k0dLiSgY3I/0RHyuRTckG3ESoZkilLDE1J5/CfXq5j0uMxVwutwi68dN4p
O4KEqwhajIv6TGVmdSAsvtScRznm06tliYHFFGAhAyHghTZikUpL+8P+ycK4IKCv
L5GxiVOzH6OG59J7FEqkV/qLz2XvDTSRVtQs6VlwrwG6+itsEXXTY6buRWUuNAZL
7FUOGJr+OPt5FThQqVOeHWXqYYGc23YzjiQXqr/78sJuZKSrEM3D2vJi28IKH/t+
3MR5c+072BAda7hpetEqDOtj+pvdYJxt6fIZwg5nyKbQGmg9dyZblza8cMa6K/tN
oG/aMBwW0N8+qB/VJBZoaMiIe29rYp4V6gGP9W7iqI3dpdoOagyHUtwOMoBZpLLe
y1AYDDESAooY52c/jLTKZt0T7wzvQepNquhkJqN8RBiKr8qQrHS1hx1buNmdxVoG
M3P6kVebskS/xXbjdK8vbDpg5XvfhT6IZUBDVdByHfFVlLvmBt2SUETpIi8mn+mB
7tmxoO/kPTbKgkEgmxR0hJLBsOOJ1fjWtLH8Zymz9Kk+R/NlRJzTC1MQZz4w0mw6
Xzo2GP6DYes7q3A4jA9w3d+ymb1sLHkN/UPu9A0PXkeicPQ7FJ96Bm2GqoxiRsp+
flG9m/4wYZz7kROypxkqW6JV6goAyOp9d72FsvQV6n8xuTQLmUzoUnhDYHNKMAgQ
uqw3R1DvX/eMVEf64wJyz8UfmPTA2Naus3lgtbd42dJtzdv/ZkOpU2BWyCrIzdN3
Jf5WBQsSB1y4TC5ezixGX7Dm3B1NWZNBxBW5V3PkWmBkl9EmKRDl/ie8rYJ5PwFf
6splUOna7hgOXrqzKosx24mBO442iQZxqC2+M5X1lIN6P6Ud5ISG5E5bbF2qM5uE
9dl0auHOmTS41amvH86jWESCUyHL4V1Wi1TMhYCUdeY7lnTKlbXm7Sl35NAeTJxD
dFAGnFTjkxwFL5uEL34iunsJypVs6ADACPJDu/UTLSubWXUeZZgjsMgmyywYgVhl
1P90fspxn97RE++/f1uxKbEHRFX3ejaxrKtotArk3b+eCNC51cQokPM04ek1uMq7
EHEslQYtZYRD8WUW8UCZ3QhzDhgGAJw1C2SqzFzKkBpCCPbHD4c1xk7DfDuHQ4ix
juk6enANEh8aYFWKF5NsdNmIFXOCOO+Rq5StygBYpWhpADjWHGiG7enARm1bhPyx
WS7fBBUFH+JEoabHaeCfcCHC5JQbY5UYxzD+IRHI9daCrcamZ9jWyVso7tbsbZ+p
gTUM2kg3VXOIdRjEB4CYbffhVz+iEO6ioqQzHMOyUWPSGLMLa4k66MAZz9RNrBhk
KV8WpboNNZhflPbcaYD8Wg9hGRYBZ/dz6FEBCsbvXMAxcy7XPuL6AiFQOqQaaZk/
c35zwcAgFOTnPLNWbdaLpUbyDGSj5IlUl9cgYeszRHjAITaZnS35U/EzTCQ8MVHm
QC5Mo5r3Y4tH30JVQ9nCD3rOFuRrtOoMtcdZg7KCVQs4XqutPhux/rG7Hax92CYh
GC8JufUDWrJSJPmvrAnQBP6jNeWbBQQJBywyqZuvzLN9f+AoKtXXGHeZZHoh5dM4
LwP0911j5D/t6nF2qEpX6x+nOzmjEXWdAPazfQPrOirjYUrkuH4dh7klpL9VTpDJ
2hchEFl4dTJWvfBXLvdbCmwFc93+SRrp3n4m0eavIkh1kHsrA2hti6/zSmrmHxHf
lBtnB+iEs+dbZo3NRkXRizWsb9tNPNvNmytW1UFL7K/EXFbDdXVJeENd6EuM3fgo
cHdCS1NyvtGC5v7qxH9cPS/+gpVzPOaSMhpd6PQ4Z3v0jzdB9CotlZzIsSNVloQV
WQ2ZPKSC13HmINkHVW06aJXCCbM0rnVRjgqPdQgr298T3kSoS6w/qImLjG+jxvOD
FOuM/rge2eybtF5varMD+4hmdtl2sIeGYJ/y8mHzaXC6ydYyqjs+fRr8s2aETaCB
Yf/MVs0LMPJZdTUNBItDfy1zxcNsYfk/cbDaw+ef5lXBFRPeX/2+ifKigNR7IuCk
eAiA58o3x95fRzEmqseGKLROqUnTQ3xW9+mpLmHjJqHIoZ/W+xHIFQ8RbKsW9HJ9
MzKbM++CqdDvUIVjr3+8teHTVVEUj964BCAsXuRNCsp+L/HOHYG//DsBmuZoeAI8
NspgH2u/5GgwxIMcn7E1qkxWeKf7twVa3nHQkQYh1d+8vYvKh935rdpAzkh8eJiv
icfpfWhXdaK5xBGj2hLGY/wRpnh726aHlW9tDcJNpaHsEeqJzFM1WXpykAZf7Bfu
iGTcE/tDAhiRE6tvwlK/8fSCRFS8mDWcy4c3SlxktsZz1xt1QCmUG2LXql2tiyse
g9GHS3XoIvBgvI/Kv7p60BHkbCRPCPYAjz4SPfUTeXCtKMJXTsssptqaF7x5uV9I
vez3MirAJeB1hs4L9ldl+QWSMII7P66jQ4lQVi5tWgjBjKzKyl5ypshJazzFkY2F
Y1NEH3u6TDuxOsJAwSnncD1MJ2plUTcH5QJQbposrMV07mIAZSy4dd0veuK+Vb9V
AF89F66YFuRArMWfqLj58NUkE+0y8k43SHxYRq5Zt7hl8jJanf97v+XdjlSz24DF
SqDCR3IK2IAu8IpyW+Vxz48ZltR3N8Ozp9Yneqk+mfuSnBxpiokE2rWdgLh4nOMr
dJUfaFEVjimxLbRJyrxeylsCuYYdQfopr0KrL/zgSOuO/b+VUViZb0R1TmI8X7Ar
2lszMZMw8QRW+E7k80jCkpalVS/jVwsAxj4zGj53W03d1TqIE6Doc/CCYY7KsW5b
nFrZmaQPmN1UkErgBj01zz0cYbMTgQCPeKUtTuQmzcUMslGUD1VvoKDSq01Aejbw
tCga1XQsA7HJZKIGaa5dKO5owBaP/HBrwRJcJXocQ2MtQ/GI9KvCvlW7dgAo41si
ITXFwMlicZwftt0qccvs3+QiTQoWI1vcwZjsZ75UwMqH5Rii9g31eY0glnOzr44k
lhwiKZHGWci3xaIujooqmjl5BBeyYJo7Le5T0vd7BDh298XJvNRcaK0qUJpjjVNi
sMAaLAD512e7McVqT5FPJQwmTB8XzMfp98M4Cu15dtifXcRNcPY5Lbn7JbghCPwm
HG9Z8b+NrpiVZiVXfDLMepDmhFWq/q8WKo0abaTcyBu3fpRgEW6u3xiubPhM99j2
9EoyAPhfru/aopV6Qk7gCtwWZ2Z21z/Sz5vLHzZm95lzAquMjecpYiLIfYQIL5hk
UBkOVQOZX+kLnGSc8kqllyjPezhwFtFq5ptpA6H7uUTyfBYozigt5X0DtzhpQOee
zpi1rekHT50U/Tgvk0+9UV87yHnYt6w/GeBrHh5X/ZGwYHQYg2gJUs4c4IL45RWu
YElVELDUz01E0v9fF2kH6T6dNuWSYGPTpGvODyS2nztDgPzH5VwfTMzy+Ct806vd
RYiN3kksFftmMDt6K/ZwOvgd/VXl8jK1G6QJwqUd7TZd6M1GtnS4McpHSPj6H4Wn
2+mayC49VSFqbTXmm+uqyE/jucZIIz+Bgasx3rOfY1fFGoZi+2DBUOKi7ikJBkQf
vtPFfg0OqXduHGTRNHB1/2Y2SEgSd2zGJ2VEh4ZRRkP8qlIL4780JoEvdxeChV9z
AdlR2pORUhiTp+eEz+nB0fR3JQy5e6t9FYY4yvyuuHBKsKT+1YmVHPAugVfmZb6y
etKMH3bLI463b69tc6mlEwxzs2x3GC6RBwSMF07OZu55O5jhgYy3FPNG9h7YLj8k
4raf7hNXcLCrGxwXoJBScNKGo80ElGbOVjjaBG7eUdYXHLjds88ORwKP9gE+oj32
DlJuLrwJVbPQItYnTch6F4UK0g4S2HGqDIuH5NO33AlN6AJKIf0s6XdQWp/jNKe2
fn9q53ZpTTifP4O0bJMPYjGBhgtOAVOMsIg6mMXMAwhFx1XrKkEMtt68FdAZkiqt
xyCKcyEW3qR2FsJb7NJ/oBD3K9+8rXnsE+jpQL9ZrcC5cWX2J4iWAmqsBz6BS5pg
syns1PesAO0ZORcGFXW+uo19gXrwbLOXBpLd5XqGgzjxFRO+tRBzyFyKxeMUMwgO
lvm87Vrnc7cqOCn2IHxMD55NRVvoVy0I62F3Ubm16gDtLJvXlH+mEWFJXk81c/3L
L/p15TbpftuMxL2P8OvgT3/qyzDHHsISy1lvsstwyAuCIsonTtavWVW0K7TxY/Io
k2g2RKxm6S3HAzM6LDEMoU/CMJvfqIGYY4vjM7IC/zzWpDjVEqXb1/488oodQ6iq
FzRQ0k10jo8aDWfTIHsOOG+85rmLXtuxbLwLAFjySDk55RdWyu49iB0RW3GExZ+4
Y6nZZYcTPwGsBBDhHTATQIfrnpHMQm2bZpLBtNejcCJ+n6aInFpRl8V4ADGdaP/b
ePNlunPe6nasE/90oaSvYcdyPh9XsV8A178Z2XLTDJ/86G8h9yT6Qdf7oPfuQeFD
+KBXCq/Wb4ZAv+27soxBaHMk68oe1+7JAQ2R89GIKemplBTKRwkFAX9D4n+0EKBt
W+g81DM8tzwux1EphyX80/B8wZxQ9CRgiBk6nuVKhqKoAOxPAhlYTdIr16+wSiio
yPXH3OBY9+XGMYPZ+uHIH48QRNKcVmaF7imEzE2YoXSWIYmMOKIMpQSlpgLpHfNi
z/BIls9c5NE+85vAk6utFShc8KeMCN2/wQEEj4qm+SsDWv3h9O4KafsMPK47pl7w
NJQaZXSp3BRXzHrsQa02ZrTHT20DyWFO1Zu6P4PhjqowUTWZHpSLGKOFJHQDEtIR
1wVRUxGI2b09vr6KgC6O7xMD8A9KlhNoZVxHgdxs5fblQIu9KB6r/sYd4M91G5D5
wZvGQYqV0zCeLN9xr9A9IzSenrNrs6jaevftPa9lA6WDMnGT7THIpQSpMc+FoSFH
bjrGPpWJwdqGaPq2I85IgrW1+sUswsp5aqYkU9Mi/G77O9KAvtqNnPr0dJS8msJi
rt3b6eCFpVdtoNSkwhaqjWne80fgXVbvvI4AOGZUm9sVqW5cbsYPL6WDEiImP4xz
ugu8FYwfKsLtRkuot/dw5QwIBpWy5+cTwYrqThbLKvNvEc62kU+/p2VjDt9h+NZC
ITAzoGQhvGmSSFfHNWHjbRXr80ouqQtL4A6kLjPASmIAxqv+muRxzy2WJiGwkENf
qYSpv6H1MWV0YL/RxrLsgVi9usqtEiGZco9+KAeQlzycLOIp5jwAhyPQafiuLCXG
cwYn/X3d0b4MNI+KcfdDy2Ftvj9VYO9HZ1NcInRhPp2W5H7DDEFvUsulk4yMD8ny
zxL6l9+DGDe0wB/CpdFJa7OBtGcJ7tuGAi0pGN1objlZ53udT/dAcOzobnVyBsKa
wojKJFlCqQDMOcetUU57RY7zUctIsd+5+St3iOZn4UEIPwU10NSKGYc2jMTWJPfS
eYFtH5c/O+u0zNGVeBEYUAg7feI8t28c9kbNDUHrr+gJkawPC6GvAKOQR9ddc1qw
099R6/4uFpNvLuQ3X10QwHYJ+rRu9g6ORNjVM01Mr9ZlVLZP29v92f72t2Wv1UdQ
u5Z6ZjfNfrRtKdNkSAcKbVuxDAbEbrxzCtnMBIY90AK7NZPPMcKeAjoDRv23NdCc
XKRBTsYXogVtDV4yH8WFFemNu/pInfApMrBN3OKKHiJJobspGIY/+y0kufLJsDvt
LuWCaQmicGri6ovQUdn03jAR5dnIIxuEHO39Tx4WxYdgSuQyFRvnmeLO6bZdULjB
8nARBJur1cpJlRar8nIqwv9T8tGt1CNa/EHgslxvzG7a9qSp26A7O+28jLOtzGn4
rDGeWvsEnt6/VRa+MeDNu+DYUCttAJ4QagTGLI9StOgbMYXk087pz9Z+6h4xXtSG
xfgIpou5SqbCQmh2Orsy6F535us+gxD9Pypl79Tp4kouINDhBMhzNHc1DgEb97DF
YDj2kcAezvhkISp/9SlTX4g7louv/AoBL5aotO1Q5sNsCR15tsvnY+gwHlukNS07
25qbx1/IqAKpyDWu7VyVBRVjpvcFSA7V5tqSfUOGfN7WpM4/G7QjAIEZLfg5LB/K
5XiHY2aivkJGncPUEOLLy8o5XMUAde5Bqa6DdVu4NsEY1XM7ZTPq2U/cWT3NjkdN
xLAo73jKybekJ/J5vEvNXxaY1X6P7LvD924HNSjjkJVfgZff2hOk+RUN9oWlInaj
JexmSASY2uADwPdLNgUcroUYi9oBAeHbxcGd4QX63i3ScSs+31HUYLZ0Q4KKCgye
AwPT6w5izneVL6nM1PyHxaYviJIcv+zIDOCO3Pflxh85hwdvZTM3JmCLCZW+6uFY
H3lkuzS/7gx/NTreNARvDFjlI3yzf++4IdnwcVdSxLWfAj7x8dEqEXlOfbIbSOIy
2e4+22ye62s9eAQ5CtpTbRare9/A4hnaUvnADINWM+3vTRPPFTtf9XQ/Pq2SjVle
n4exVmoi7RsoMAnh9+479yAamXnYfMBoLOdZZxed7Yded7p/Mb1/2uz8WnxkFnCJ
9TtvHyy++uJ6XWREzBNqrrEG6ETzDg07wO5lpzD+kRQvKYi4DeH7sz2Od42xXB7z
vIgwzCNzqMkfpM1GeSTLFRiYGTb754iWiUSVYvtrudloqGzeiktGF0ji42MT7Ad9
ouh6AFBkiIjQugHMbja9FJPzEU4NXPAmSKNHN34NqfmcQTEXkUYwPx/ou8xC5cHI
oxGBp6JYH2ysx2EP0WNTHktruyCzPEk+2nDSoBrmtUck2Hy2IO6RTRjsAeRu1vAT
qXEO6jgci0cPhs96WsgLdxkcP+C1UKb9gNZ4Oi1KgOjRKQQ2AzlHuqkAfHWs3w/N
4jjnG23QAOWMfytmXQP0B7ZoHIPlcr489/6Z39saxX7ztcMyEBuTF332FgKYzen7
mA/9iqQAeCUVZWc1wytylIzNv4jbGWxEJhpj/9EdNWo9uBF1dj6TgCbuGusIMenM
XsVhE6NfddmmokyBuyWRHBjS5LLaJug3VPTKesSDpDY7OLWFcjWBEP8duGRY6oIq
VTp+U82KqQiuoOva5Qv40B2Oi+mGpZ7KROdeeyFeqY7r6+ZUIUq2s3ly7TX9oRQk
WGPby48cPw1mwtjyHOEUE66aF/96+jYJ6QgtNd3s5O7BcjyiFJ/ClXK14P+E3WWF
zW+Wur9X0jVjL+1CT/Vo8VJE6MD6OZw7ezTyqth06gXOn0tJjVZjjq3roxGBDfGp
fNbJnNW16W8AE1TAnG/Vq3mCGWcBtovZt/O1oZPMXv1gfQ8+z1QYWBUbPOjtl6Mq
OXf6/f0HzeROnfRtEbB/pTJbbBf/ol5K9bKfNzd01s8iJd8XGFoCrXZ1MiHGHv5T
Bj+XBaQULDxYu1DIC7HjmH5/K0IH/W8piPMrwgQbEiheTxCONG/4RKrJffqBPrr8
qhAlaNXhoruDkG+uMvtk8QAHdH1aIlYNoQAWDgGnuLiL+I/SUaHGU6HCmfNbkmnc
wLFB50IUVqZRL6BUwy1EJo15sWFlX9mU015vcXcr3LFVPyzJYa0ziqKL3mSrN2CZ
YyVJLQE8qB1igWi8995eUQSMm/wT4WPc7LPPEVeg6So37w8yh+PTs53f5DPx0Go9
IKcZ/F3DKjXb54QXoe8LEbIQSi+4aOn4GWJ4CinlkE00zOmkgcIFmAk8nc/AJOTs
og3XvwOC6v20Gq60xzBt7V7RmhmgIQPL/0h0nxE5/8IDPs3AKT1S2rg/NZnjkhY/
yh3BgiVWL3laemvPSy9qhCXy2qvxsm3EyF+4czRZU6oOdwVfUHqeeJl0wkXIIcos
qAAwNVFCuLGPbqVr/LWryrerlr+jWEUoXYCXSyUXLMn7n2kWBsrxp686RlXXoDLO
42LZy0MOGIFfV3croQHkL8lfg/I0baWo64bvP95V5UrPh38VOxL5/LY8ib0U8ZKF
sTmm4kwc26qly44KoZHGeI5RxR55n9elA6YRuQjsZGGRUyzcwT+QDqPSXLO6lFhb
A7doBmNY1KWrmEAcnPnVrBI9BfCVOFt3GgRTpsFIqaTfh6/1aAli5LMQxtUDGcXd
w1JcR6JqOemX2vKHeuWhLCiL/aSIIK/mjoUw2SxzE0kq+H0HgGtfvlBDFXSj7DHz
KfY62Rgq106zw7ahT7d2hvaEBLWmnjrc8xlp+0hbv8pARkN3Whqj30fGDE4Xay8L
T/jlZmHOKLfj+DZHjMsrjDZoGerF3fE7r+MKpKWYfz5f//GkFBA1VqgG7cpMRNb0
VpRl4vdeBysW3XoX8BXuE37ykL8mBAlw6rZMTOWIJWGZvPMsiJTnesZpPIDt67CS
BZFrxEd2VvsDk9icbuM1nV5jdDhTf76QDpb8sgeq3h7wNIxVLyNGK51A/Zylhjj+
qhIz0+TYWhK/vJDmnKEq2ugJgoU0kpTqugKsPNR7vADNCPuCnLyAI2/iAwUF0j/k
oY2NNXNte9qvm0TTkinQDcLN42vsxYS9/CjsGqs2DEoFCELBX/otTANGqUeDyjFK
sO0UWoVAYSsoVllGbjzBhINU653Qn4n8U/6b4IimJN413o6oFpMM98xX7Z+HDZc9
+llBtF9ezGRVGoUZo60noP4bdVYkkn8rpzvwxvxD0XflD/5zVCoSlLsUDLejg424
w+j2u+EepNODrX3AU+ziBVKPtYwDhM5eXVGxVYzpCKz01kWjX3j4QwRSioPN/3jQ
0Si7zo3ZPx68ycWzs4uihPBeUKECCefsw8HCjVdkDQG85o9rBgacE+GmUs9OBiQk
wSDk5QI/9Wph4xJyLmbfZJ/YmYqXuN9U6yMWLeiEm6IUexUOQ0PHJe3FjEE7qNUt
j37kNRvexq9VXWZ3P99GhF4udSaARZLAzK4gZYLqcWtgsBkWuhD4LQfHoXUltWbQ
CXxNlHa+GwXV89HrJX9s+ooeZmrc7z6L7QjWuWlX2tJVM/mqdLnXFq6mfbXGrhxv
fU6Vv58fw40v2q0UIv0jS+jfZ79Z2ZCNzYJqLEdg96nhZJE4MfmQZZ4M6ru7ldHb
4wiIynNJ0DSZbTuN66jydwQrvI7BrRFdtN9Vv95BA61WwImXFW+jqbQrjxphR3mM
ifKuRhD/NCWwcgdHVzxL6VejCcI0Kzvp472lEShF6qXwZLMWC1eG8jhkiHJleQqK
/jha1INSBJf0oIfpsQTohNuGQmlnRSQecvhRYxigAjzTyW++DvOe3lQ1Zfzb07/1
Sn2RiURNUa2GgmdV51HU3fZtqGJLHgLyoKC04thwPhjeMLgfFCI59sP8z24rkU7v
4CW04zK3GDe9pgzFcZxry72/ChYaTihOIocbbihQVApEYabqMWRvOoVh/k9sTizd
eoVHamSJu9QmQHrSSH+iApcOMg7d1X7497m5v0MSfmXdCdG287xkOmnbGpnCfpyv
YdnqgjSPXT1pu6U4s5vDOwNB4HC1eyi7+QVjOngaPKeiQ7pBuyv2TbI5dEU7LxXw
1gJiEKmyWawlAjAk+wQr9s7F7EeU4ZAA0u9M1jaXEZDGsDaTlZYTi7z1cMAjWeyU
aH5G845FsjICzFgXdsQoei7MKmAcVzQVKeprWOk9+OVqUBARhMjkwB7rRP/5CXZg
Ui7Dso+ifJVRWa7tyLxlfov01Kp6QKpvdGq2UW+/JqzpRmRMDZn7vIoEA4tlf9ny
k1LlaU1uJsN816Tn+zh6boK8ljJPXy5xPI7pb5KZhNgMjUTIGUc4w5iFa4NelG8z
33LrfEQ9N0FbjVG2uPLW4QtM7KCv+2yt6/BwKtcDFTlWuTB8t4Vp29OtVSQAt6Er
hhHMa0bkUkjgp8rGAqEKbdXK3SypJkPEYAKmFchWb5svKCfSzKgBSSQmzgN0cZ0+
N/HTgnTA5ztJGRxxUPs/TLZCVWT1nUM9cAZltA5Zow5ZFlMN1UnfHifc5EKuZ/mN
nDQGeUs+vheoBcLaDxIVIxKFgwgZT6BqosP/NyHjbH8rD/4650AcqDlBWsWG9xA2
6afROiC0fN0hhGMHMEM7KnPEbogUwcU0bUqWJ8JNkWGJmWH6xtC8Agr38iJkQhVL
a7EuP9NGM8jsdu3+t+PJTYsmHGIeS2KCHOrKkCIy3rrFRtpWtf1ltBsLbINDxYvx
0KtJjgrtLTouWzmTjpo8ttQA2pwaaBgzc/htO/pTuDEYe44zfO1yjk53a2TlxdAL
7e54VJW4n69YM4uQ4fkK95vtLx6XFhINqppA87mOmKN6mikSQejkpRC+2KKJTD9s
+jCwMGVqPYzwfRbQR7XQgbrYOZzaauRcl4R55JQeg8yUQpkIiDzE9pPuHhC3CabC
Cu4sEFoRarVF1wIrjzi8YhXdx1E7IBiFXELrVrZ78jrYpPWPnhn7j9nAmWsK2wIE
HiRAuPNivryUORMBjA5WDyvOb8NNEiQlHs5XR0PYfWbt2Yfu/9ZFbSqqTJw4ERRp
RmGh/i/2i9iMBDxnfT3hfqqG4fewgYikEaD3f+LGa3bC6gBNAZMrdLVlKehQcofm
T+GPNVr6Q9vOlaBA/SA4Xn5zDgBUFPTPfMLuBoFTcCRqDfcJRTLUo3dWFSLbc0GH
XtMfccg3tm81QjArWyaDHqK7SrTLctKbr0nIwoVMNc9C2+7EakIq7Tlw31p65S3/
OVT9iYbl4f6nLKTl8X862CTCUccId54GCiXUBPDdTonSiuZtt4RfuIXLWEuNHeZ3
D92wr0LcN+ZTcyNOppO4dO4j73ZUnzhnhh+yfcIUX1F8z81SvNK9WkkpOuGb2cQe
pwPoXI4k6YLDtMMSjZD5rsfkgbYpDk2c/tTU2BZzmJJOE5YHBfxa+rrxMqMSIZC2
uMYPEuISs+d4JaLrGy1Da6sT1iT6DOmfJmMAJDjGg/awI6fEKJEUL5ooe7V/KLDX
F3i93DM0epbGqD2Gz7U+qTDqqU2gofRPt5v/GG8lrUBj1CMU1xXAMUVB5onRruE7
8ywxBO1VGbBmIdee/kqYyi/wgvz5pCNkEaT+N+Sz7q/8LFiSfNcsxW7F3Iw84D4l
nn/CIlm+P9+nI88SpRXPrfIYp4r7YriJVJ3VbAbg7OHkyC846b1kjjoXt4DMN2nN
Th826f7FzbtiqXg/SlnqE+HzODQTqnnBs3LVqQIx0pIoVrzbsKttqlGIIfCO2CNe
uXlndG980rS7R2YyChGgSaNLIclzo8jKfzlCMTGPOm450X22Vc7z2NSqSEpJ3M5Y
+UJRwVEg3RgytVfgliBo3m2SkuM84llFU9sGKr+KGUUBCLAXhX5VOZ2bsZUAuSwR
AtpUas/kwmjVD6ksJuOZuxUcel2T1EnILeCnlhzbwJ4NjNqlK8ZxCOUMZq7l+OIz
RZdNdU2tpLhGfFptgDVE0nnCLQcNQ9xmy9yxV/NhpOEcGyXD8DdkVTF4C70Iruia
kQApo9JbgTOOwXMi4gb2MD+vmzjCLe2DINyIEDaHLgwC1i/f8dnGWG/6n9MTYS9i
QXB2XK5b/c4SXyqz+KuZkY7f2GH6UiLIrv/SlxE0MdF7+hDOcTmtJ4C3DUuSzPIB
P7O4nPM+uyFRvZAdiVTlgBjPTjf1Oedp4lonb4XwPeQgQbMEi1j6Z2qnB8yJ9hmp
5qMtDEdaClUx/7UpJyYvu+2N79jRt60sTIsZbNwLmXOBEG1a/qtCYaETrtgjmfm1
a+GdUyB8NaZfPK7n2FcoqT8TjnOteaYrbGBoAhdR+334Ca0HzMKQZsnmRaakSgJJ
gtx69sYQJLJZDlrrjyMZBp4hnHBuJaXcMnQuvd2cyYVMklDkYFgidZAt+Ocu3kk2
siuer9xEvzWzLE/jLSUQu+gTCzSjkyQKI+GcVN1PgidJBIyyiOTIzeR89cvqxJma
cm9f/iy5KOnjiAC01R9y61eQtcZ4rTDBPD9Hi4BJfwwuoB4eH0GCdfJgBVL9LKI+
2y3oxHY/b1+D/89FswPHo02FOGh91CEaCdfk4yig2F1mfGITRXyuTmnKeOcW6RRl
0BvtCvaPAKDuSWWFXgxH1VEm41UMT71In44Taa5ciwL3NBxxFVhKJgxG32RjCHV8
CtR+IDHOwNSBYuYUg6YUYEMfLtivdyOtvNarycT2HNM/mO4qbWVIL+39Q9DJ8DB7
B9WeU3OtQ4vebPVY35hBuXQD2vveM1yp4cdoyn5QVXNItpuePbZBRUoStF7vQMZI
ZIoHAanfw9vBxYHAMy2EMbrtMBErJz5KHENeSp2qD+giStti23qnXpxE5QhGOFie
lGg4WLUw/cB5H1jOtKDxtvrXHAVJe70/OAO3K1ylXoi4XtDAy6UaNNNyizXVAAmN
h2XnM01n5yLqtpf1Thp3EFFdRt6bEi2nedF+qyR2COaGrrg0FSFbk0HeHJIy2Et2
1UjZ6g58I01AQm6W2lehUiNhX/7uRqLFw3Zq8BEv1lVYfrg/q46LfJl+3zlfJ8BI
rMwB8JMRqB9vsBWsT4wSQS3LNAyLmAkwascdX+6ZwIIYoRM5c/pyL2l0fFvG3Inz
HoKbhHlF59e27N683B9WdX9yGIa4XeEEgn0f486NQjhw9W+4rNFuU0EwvUwxwehY
eo3MINvmhHaKSSZmzIJLr0yb4LDgddGI2f8DX9jlSWVZlU3Dg3qB07xV+Bnc8g6Z
DQaLoMuoMakxJzj2vjlkGgSDitmbSZwYpW2+6iKr/Vev7c/kZvjJGLE+DrKZ1ZcY
pD6jscQxlRPycTcoCAYxlIcDvPG3KTAe/qawTB5q7jPqIQwVxEcegHXyTLHCVRmx
u63S0nd0e4NBTTVmDL9hztj3/pTapd25Y5rk7y3X9mATugV+vfgin6zrf7jNYQm3
7KboauoL2HeG6lLsyqLD+dU04vALblcUOSDoaBWpLzuw8Rsp5AmXuV4MhwAEqXcn
xonWSzMr1ZPm30dJjjxPytwi+vPjf01tcXaZEXx7LHQi0/LdnWggiV6omspb6K/d
n+v3v4jOT32pvweM7llDyVgsLmGpkiMg6lcjuAR/HAQTaZ9LS8Xe18uCeBgWJ41z
14FLGdrYR/eX61jiTRfxkbpovZmZvSxYWv0Rz3PLkLsxkSbfDTtcnzsJFefg3MGF
DBU6Dwomno17doZn4slWa1LeulR4oz/JdA19qECQ1z4kDQv/lCdjfGJLbKMaFswp
wow2DYolgg87wJMjeMaDOuXXESTl/xO+Qj0ksLFi2Ql8Z3r+jjzfK5e+I27agddL
9RLj/tyLw7GyYLgkRXoRY5geYoUbhDgy+2SHUYYGPKs4P7bllVrFMpamsYGZzv1K
dPPkkDhSNlpVl0SHUAQNoM7j+teOXt/oZhwDIBZ2LP/ksRjVGcl22/cEvXRPR866
Qk2/BaZFC2weUzhBOU6to6WS9588v8qrEob70YYQzNuIuZPf7C6eVlivsSiIQmK1
Jz4tsfhIAOBxHwXtldSi0qXrPRw9QoHY1UMqj+rubWFdc7XcoP2/N0KcyWpQCXE2
H2gDglnk0uW/82bX7XkU6OBMm9JqanfbtbRDQadVBz8f9+Aczqv5ivZPX34lNEdd
kB3tdp/qbeJBPmsFb/etWNgjdB+Kx/WK/wgJsRBhORWzYufowRj9lNovjHm3fc1E
EYGLD9HKjecY1KrVKYUc+Isg/IY/viFM6MZ1Lmj6XqGUP2wh/l1U8HbaNU4ogGdH
GUD1349OnlKHPmLE1/zs7cqfqLcC1W2v2ZVmZaramsPETpD9Lujg+PfP//yhhnSf
hgTsKuvNyERnPMtMzY9qlTOVYAMbRavmj2PKZsBOCx2nW3/oHHCBjJeKLtwDYF26
eF1lnIFnVlEBu9M2VVXO8jLU9NjvFS0mo9iaFU3Off6ngFCSbvQp6ME/qn/W5wtE
SqGSYtJ6OIfTK/Rvy8vvwOm6080uUyIOY/+IWoEiGx3HcDSGnYqBqpjx2P4/rwKJ
lONFBNjBsRlfmiHwzUp7sJK0RzswCWXwgeZOQRt4ocm3iCiBs/+2blfULtBxSm89
76htzP4hktSGtAlGhT8Dm4GkDf9Kv6cvIVUui8CufpXpQCjAUcJnp/pIAc23xdWj
B9aQ9y0BCrm0CQTupXpwBH0E9h9bwMO5ESPz/SRSn2qvRA1VoRROzoCfOrNIZ0O2
/I6lfhmYCURqqWfHV/hFB0AokMW+6ECHtCWcxsUxO6s+99/Lm01sdXlCkkKHU1Ca
bE9KPOdex7KjAlX6hI44nqtI4sQ5NywMUsQLD3bl8ga+MDUyGHgLRQInrDnCjtf4
6GqIzeZlYb/eyCgLjr7S9MOg0hxAHeXNubDrjPescjkzwCA+P239R2b/EvrdZBRr
DiSZFHxoxZQTh8NocsWnjCZ9wHkFvg+uM8CTjDsZOJ9qupMKVB8yLaYleDtD/GKR
uWEQ8vERn7Lmh5DrpsKWuyZqwaa0GLjg53A/P0Z5SUbQQ6QgGHpsQvOh9za6aQ3k
Wu8wWKts1HkjAauMWsA8LnacbX6mcAhsoLUdXEoB7mBn97H31uij1D9mHtBOQgGF
yM5WDsv+4g/Bc+zu1hGwbPqfeVOO9npUfYi+enXCA6/tWXUoj3irTPq3BsjrGstr
iRplyfZGtnGiOel5mNju9ENnLvTW99LqaWo2H11X53Z1s+WGm/McpVKi/bR78Rp+
KBCvWfl1B2H2LmNOHVl+v9DmA2C8Ps8Hsu0SEp00bA+1NDL947s7OgkK3OwB3PL9
YbhxDkAKMbi1CooxvO/pNW43vtAOc+nV5SXEgTgaLEGFV1ovMaIHFNqoMHYpSSus
dQ7FUmfrY5ILJirN09aDnbi8b9CsOq7vZ+t5CI06YNLYewhRbAtquIbdWduBOqWE
q4tbuPDSkEog4AU8ScP4kke+Dk/sK/L88Opauozj48d/sxif58WwcxlNk/15c1J6
jybE/hmHASgbzLJPcYXYi9HcG/ZHjNqT7Vcij0tRfC39SSUiIqVzJqg9OG7Bwi4Y
qNN7lDZlnoaAo7uHjY0+D/hgEnYIXHDVzVHqj3gKg6H7uRl5J8azbh1p0ds+QwOv
Qgg0l8IKaTNnvTnMe0McQRpmT+nWgylOdxbOTqQHVvGxEmdsiHvZ6KNlVTLwFlFN
22hHMY6m3eOQP41+TfKGAtpOpGUjW9xSsp6oPsHFBBwodR0wtq5PSQi14sOO6bNr
nIGOutV4XH2p0bZdO3JA6kD4RpkbR+SHty4C8tvosbjM1FCZXFeSqO4gX3dZLnWi
MgAsM6cVr2OJbFvmRujk2900iTi0YeIUcrbBg82/UOWlC/YRuF66pyVvzVvLnrWC
ox35V0BFeySTw43M8A5oZae+gbUFCSdXc0Tse6DwbwdNUDoe8loLPB874GApZvYr
ftMXXPCO6gAqbhNz2uydaedauCQusdeMnkXO1lhNHQfm2BpVaxnMBN+zk5Xz4odT
2l0rSBwFl08qGdMfQ1T2ESm+DN3LMMhrpICY9jriSLp9S9YWoEAsea+J6PP5GBrN
Iszbzkt0ncH2klYx8UnjwWPK07FYPqu8nciHDctoOEsROGx/Gzz5ju1iRrJqh6vz
prNTebFBJEntAe33sWFJ7tpZBVsoDmlXCLgMGjsfzzP3N0EVg0cppj+/CIXlRESf
I0L+q5izcmkTzkS2yzStFlpJvVCUBezSz+w0mheBwqUb+B/yNhGSfzizJpsOjxlJ
96oteg+Js5UccgV8JX9deVO1ZKpcqp2JlgdKVUPfqJnpNgRc71QfuGBke6lORcoj
AGRsiWTYp0NVVwtsW+CrSlq1rMIZUoTBoJWRGqhxOH3eJtcMQsOpiKo15Yjoa2Cs
JeWBjqHFd6eaDwQKznP6R/MA00pyydZftN6+CSiGim7CXNZfma59W5sSyf1JmaaN
pMS5cbqLWJ3CPTDeaDOUr8UxfGrW7y60xwo3oyabrimQrNMq6Z0Dx61Y04TaSIBw
zBNlbMtDUeKbt4u0K5S33dPaJMmfY/UYF3yQNBhIHoU1u/1jxcbkfAon+cDVCGxX
/clfaHUcYgb6LDzTqrNm3uEL08nMASriwptA+E8RnSON1L7sEim1aEjrq3oS8ux9
5S0Vxg4Vp0UEYAPCvDDlZAS49ai9QmwIymSS696Uz0OWQ0A6vgKsuw7/mBryWUQp
eyUiDEYe8h705qIjHSj9AteN3wKmlnu00GGT8JB/Pn823qsWXyDzNwn2bT5gb9j5
PDcz3by/UAeV+fWeZB1z6KwLfRgECCNZZA9hFc9cX6awT1gTd2eMjQzYH2J0gJXJ
nCJwGYR+I5BlJpFVgDtdtX/yp/TNUktx6744fiXXhJGZ2gwx0lhjQBnxWh/43cqf
E4gmE79Ms5UmW8UlRxVM53s9nqBorCplOn6LQ2xqXkcbpT3NbEHtCvieRZkncDSJ
jrZn3bK4fBTbK1hmyGyuW9JXBDK/EG53zN7xwiG+gvh9d2LfYRA7c48jpR/Mkv7V
zELvbvw4NqrINB3hQnDw7dX/I93D6ZczcxdGJPPs7ICPFILu/NJh+k+j86KPobuy
mOARI7D5tr2LbrfymY+CbmFuKC+CK6valMQhTSnM2raeZQp2JnWRey/DsHlvkPkk
yxey64vnpt9Aet/q9JI5Ay2m9k26ZppDMEyQWnDUUHgMqSWa0+xOJCQgleVlW73k
jHzp3L8vwT/RJvs8D2Rqa8U7zBXY8v9kj4q0hhAcWKOvn5hdSWTq4R6xpibG734E
N2FVqKWiXuq2T2OmCYY3QTZeW1padtYd7dAOLH+OJIqrwts2bkdacO8qdnOrRtuQ
4U05WZfE8hVW/w27ZiedCn5OKcxAOpU2jOB7qPRHT8+h8uijn8XEoMb2GwYcYQAF
Z7lv+ONpSObGus/XlCcCnrRFoaYzLc9HaeSJf7SrgX5ZID4f2Om78AFal5GVjM4B
aUOjaIzxfMZoTynA1dAcjCk/UA1d3A+M7VXPsI4wB+cTV2SEZMblyCmFXLh9zzoS
4quE7Gtf5INgwciULZwJeAiyv1ftyJKpGbSPIo/kZIFnpPxwYfkeGtwua25v2Azq
fnoYvxo7lWbPrWqj3HsMkXNpyjZL/9XrK5APClh6YiZXXmMyb0jnXBZ2F2MUdr9x
Yf2+ptXRYo1Fi7QXbbo3tl0nfBw/EklFbJm0CbKwnrHEqy73syx940L1DWRLcinA
/mLaQNh3HcKSuIbruB58yALwQSrIJQhTUGZWBVWinab/30xLWnLy2SMd5514UUYg
H9s2WPIYx6mvpFxa6GcAf0Cx7HTtwnbNHSKXDanTNLkFV5HsBvg6W4axO5sdPW0W
QzL0dwBE8sP4l+QGtMCAA/I+SLTm3vE3fyzP8Z0BFV8FpIypmTJEFKM8PJRdBQ2w
Tz1t+ch+6OJwYwsa+a/jL9KxJgUXKiSmOc92j4bww/Rax4RMdHYX6CmR757SqVqu
C6pgAE0DaB+8qdih6EIYChGqU4VMM7a0tuyv44Ex7MdoQs1rKU6sXqdXEupz458G
rxhItgAEnINuG9zKXt3PrQ0cIOzz69yWJ1E6uU0LM2e3mbW3f1KEywWbLEDMz1s3
0ehPPXFzuLen6aPKbWEeiTk2u+GuDzWOHj/zCZyuprUn73EOFazXzBRjlpevOZRy
mhgnOyUuISZ6kqMSTlO8REnrJFLLXcmPbfEmNZbZbKbDl9ZPYsx5IQYYsTvArqxl
xMwTRqyz+lWOIzy/udheWbHFtVLVS32D6wFmRON9tSnG/INPgU+9OjvRpfL8MiQD
PurNRZ9hO4CQtSG4hlj4meFMGtYa3/ptOyLFARpsZvjDdiwcegfKZ8/xFD4OIzS7
+uX1EaHTqweVEDxw5rZ/MFG831NdgwiGrm9vwtIw5NBakAkpgWXkrt397yeJUKUI
pEBSJrc51cEHRGRwBougU9r3daYXmOeMzEsWikb43zdD7UtT+JVg/2JHvRUbGauF
+ShZJXuFs2jTMzfnq3MOi3hEYEYQK1Y+ldySyaLRriHPUKsa+Qm45ShnYFrbr8T4
/qY+hezYaCUjQcn4NkT1hrQ67V/RUNmeLEXcOormy4zGasExf/CquhfuhRlkeNfL
a5ry79mZKSl+zZWi9B4B0iXC7UO8LvUmlaSnfxjdK8zaLVL3Q6A4Yk1/5adgwFY9
OgvXdUMIeI2QeLshB4ZNspUMj1amyXN+lzMURgezMhruL4R/AU1RP0kbFcFF/YAk
gUwzas8NyuqcQEqTQ8uiZyelbfIzTiJj6G7pJ24Oq9rHrWOf0fJjzR0510W4tv2z
IlFOG1NfBniFNQTGpQklL2O5DW98PEFps7QoqPA3pf8NO3RUH1l2CAKfUzV+mxhb
IyfmQcy8XT8RPmjKNo9kZJIJXDzI1XOcask0eRrllnzWwaCzxARRzDiog9Ckmc5y
fbXBnc3lFaYjKmjeMqMlBTyiw/eMivtxtGxDfY2wM5qPIvjc6i+FkrJOIie71vVl
d9d8O1gCX6meEIG7AYJMgdHtjI+3Zj1n5uJKdSWMM0CWUI+6q306lsJCCABNMIjK
3yORm2td+Q3La8LUJ/zE66QI0pQHK6gENnEdk8ZvInv5Yn0CRBfZZ8aHuQ9FzGl0
zXl4Ps2CHNSsxS2wEtcy3b/W5RDkpL75DpuqTNZ2tBtb7QCS0BM5P/DsSU2SQ50k
aGhiEPvGnSedYhC28JHyXKsB4WA1f/eg6dGvYiitJopzzgMTo4GfDiFV/xsodvnn
GqMjkLZHd6cx0KCvKvoSwDVjsLu2gAMl7QoMxoAW2YbvQ7IVI98hEKL5EwXx0ZN/
ecTPu0bc2bB2SFfXBVMCrCegwCu9L1tQJ9SH5ReaV296dtRxtDgD2HQnQouncI7i
69NPJVw3QczlcR8ARDb/4l8RT5sLdMzvWsYTvsqzowgAC42qZZLM9QdsVN/aZ6wg
Cf/+vB96aqsnsyiMRiAhLktp0mB9STNwI/RmPLVl5rOVJu0JQLHrmSDDaNrqk+6O
cMnzk6Nn+zhGshssJ/WDqAtrGImFql3JTz8+yn+ntuPXDloL/CadJyKDZ1FEx5vT
1ZTxlWXD8e8J1PbUNZy6zTcRPkqg2mM74QzudUu4I7KF3ZeM7VylG4VC6l8L2y47
yH/hkGC8flPCwJPhUinA3DZf9yTI+9B9MjnQyuy1y9FgNRTAPhBFrLH6HBAqs1we
G8BGODwsZISxTynaUClvye4S7BGxnYSASHwLV+ZYQdmUfet+aMXM4h8hpRbIQvW/
O9pAgPxwMr6F0AEb3Am90G+kaKxtQ5h7JSF6ZN2VvEzreLrz+2QVyWA6Lg8FaPjb
k36q6i5QHa0M/FlYFXU6C+qXNKIETOtG7KP8rCo+aC0TkKSRzVr8Wqrb//f4g6lX
mE+En/HQkIVAIbXIGMAiErtseG/lTKVZKBFAESgPZo6cAAMHvCXeaz5dO8NQaauj
PdbIrZGQ16rAeGhwo0j1BDatObcq7IFnEHVx5Ls2DtSRmLbCLRddK5CU9ctCslRA
J4Q7YGiKYmLeSiKl/9R4FItVvqK+QvI/eBnEXpdtytjtej0kGhZP3ba87R5+i6Wi
OsT3lcKPr8IzEZzd4M38EqGFY1rzvcaCqf3ullN0l5ADQFwuYZtHHt/9PaPueTUZ
pm8cRR+2q4uEs2MrgxhSWPpU12PUoG6zenoR37VKj6WMRiY2GKBHl/hjT6K9iQx0
fdNOlWijHaBb5l5pgiY0gBqWimN76sZrhhaDpxeMoGsouGM0MHA39bHz1Rqivi/b
rBvDjLiKW9SaxqYrxOy/J0SeFe7+RWlWZ+7VBV8oVlxJLVycxbICqV07+KOrKqWn
TNH45hL4Vj6u5N7A5G9bAvNmflBxkLDmPLMSg3NjMR31UYhWawscEiKsgcIgwe/s
xuNqgvlAodwPOeg/qlJup7NGMROy1frdAccqLxiwgvGmAx1u+x7Qg9F1rBXH4Dlk
Ctz9s9ydsLahC8EDhnnD7qgARjA5j6zFtx1fWKXuQuF4/NkBzXwVsHiwuOhVUAaT
eTvTKmTru0XJA1iY+KUlar6TF+wTgx6hF1BTWKHc/VrcnQ2VpjrL4qVwbWaCIRIL
i351LXeNlc6qstb23ok6pGtddvkP+pH6yMzDqLwyQGKxh6p9umOBO8/yLR+eG6Ng
Bkh7DDpmYLtCN9stwGVmrArV379xU1y+wMBUJ6N3+YoOdv1Ef4Y+dIuQsEj1zO9I
RbkeOdanVR0gps5gIbKoAWUvZIUnOpZnxTcSzEBxG9Dwf3ikLY8kzw/lR5ENyEbV
kiEIIG0/5thw5n6Aa0tHSWMdS6mTJVqVH7rQMqJ9fTUU17wPmrfYPqvIME4JlETT
3nzhk9fJN/ROP9PzUHcPjVwvkGqUHoUaNKAujRPBiLUC0w+iBC1clI4pYvaGyRW6
bU0uLQ8TJR3URHW6cZpCpJsYo3Udy/nKt5KFqgNyXJx+jM0snu0cBVcWslEBQuWo
XDR7AnqdJ6V11S84ZM62Kq+ivvvESUAH1e6vSepMiZrj7YpVvSivb/wutbzZM+Lg
bBVRO7CJMOiMlyqfdGNOEfW4Q6utHjmxSplrtaM41x0BmOWK8Y2fPmTIw8h603HW
b5zJVmwlmtrLy62jR6td0jieuAMBFV10Wn6cyBkZd2K+sMAFTPIJTdcgWXUV4pPH
UKkey7n1QDuO3FEfj28C6zvYdUI8GxIpYGAmxJ28Ra9Z7xYFjFE/jYVX0vv7gGhs
Rl+HQ3L6pw2Knz0qgrLNquM/ybzKCP6GGaA6jwqBTwtD66pOoLmkYHTuCruztFll
hgJIGHa5jEUYc15xKK28Q0gZH9Cs3Pr49dEA8wsAi+28RucAlGqISf1flGZ3HIVx
KAT97IIVnzsFWV367Hk1bTredeSEpiPNTc0c6RIDwCsDZjq1+edmnrCzW23NgAIO
WM13SB/ZgwYaqLzqgN+TH0BTl2sU58pRz6xmhse8pLqnU8xLJsHB8NcEtSIVJdEK
VwQaZQwySucLkloNgaMN7uwCk82M5VN8CFrI8w6S7H5sTc9wPNvbjRf4e8ttc8d+
S77zGXCVwwrqni3W64G7EEzNcAsBOxbB0MW7ZNXgpAnFM6kWM+paVEFDb/XHKpAi
MefOR9PlxBpVz2uPNigd/Gvd2lo3pl+Z1n4nG35KD3mqUf6Mm7wA/pjoPG4YC4yc
wdazjWMX+ybJA21xSOW3vG/r7a0wXHY1eJOALOaKNIYgVuwkjCnbGaNzr8qyWYFW
FSWO2SKw6znGDWKWC0orShomVRK0rbJ0mpLxkmxNHQ0GgSsDGLNLOYDxRtWygA8x
oCzEe48CZfmLuHn7iMHvFlsbEKYS9ywgV4vJq+RWxo1byP5Jj5YXqITLhAkKbYBo
VHmUofDcQogddB+c/5E7nGvkfuZO5VQTLBTQGeVznkgB0gW/K30lXvBYAKNd7WL6
fQnEHu0hAqONlO/4AWRB3ZlRZfXk6yx3cN0YnoTc5LpSUVJRUB32IQIDKQzrX5Nj
7slQcDKurQYWNFPjTxficyfPxuy9XTtt5ua1e7w0HYm9R8/ITgPGcdrDk3JLg2sZ
omVO+28uYPdyGfJCiK+ZvEqH81t0/nJxkLZR6Hh1uxX+2vL3IfrPT9PyxajUpQ1D
wNXZNWYk1SmSBWld/PCLr660DmccrTYv75+2e7dfzLvwN0oqxIvWpMirS7UUJvmH
YCKWtHRqZT9lFw27+zfdKHNV5WrYd/9qHMz6ECjdObq1JQ1sEMnFJnrWclRvprPS
ZRyVRtRw2pWAGoc7nF6HfLsoV4Cvrk2W+qismRhtbSeVu7bDqFariPRTfF/mWQZf
b9u8Rp7OibEm0ktTV6t8UyXnyH0IAk88eYr3tRZKWdAYpx+M8cDdpnaCmXJerssL
92whAnUULqCY8xCIx5ybPq1hzy/fssooiARZ+xl3YrvxMbg3A5h7/nCjbBkbDqpY
IVkuuf3/MbH9uhKl1ZLxKPSeu6mPpec5Qsb+rxa8+HTAY5L1k7X3Pqx/Bew4LAsK
tz83rR/bHo+Xs3WTEzF8zQtEX6972hfc70KYExmylakVTwGSUt0ZEFBZjvcWLbiJ
pTfAGJg2GfC04D48Zl9SfMDZyWx9z67H1nfX0Wjbm8DXbXLISboB9HJydbaNAHWf
ub1RMnMh4De8tMHY9nNSU/yAiNVrIaq7aIe3i3/LZKySlZWL+3gfyus1UyrnB4tD
3AImraLXky3jM/0uH9+LEXvEU1m/Ax/S0ocdIWqFJWcujAE2m5O20vDj2kZN24gY
VIjQsKWXKgKA41AJ1vhkPdRszyrozD5dVjZHez4loA4SnNQn2B905n5Q21D4wbBo
YnYP//zy5oAl8swDtlXlOOA8q+52X5E1O+iMWT8LG/BiBwuMna7TVHX6XzZZbOZH
8RT/GYuBbbsC0vfB/j3WxocTf//Ur9QYskZWjVOJhNJ9iwua+SjstZ3dHVpVaJYK
vQF/sLaOH1LCGGfqUvwk1ma4J5OEG4QKbMsNCdtiJGeIhHokFPpbyp2QfZo58UFo
ecUTzKkgIum0doJZ40OGcbGcLxvxilLePpA8EdI/0WXay7pePFhNNvouI01EQejR
Vs53AZOG0/lhg5rZ7woQXWAcbwW4QMNsRidq9k3rvEetJVqVUn77POFIHNu8Z8Bd
X+qn2gNi9XBnE+No6hOHoYJcDJW7Xu2z2Hr6tBO8BswXP7c1kTkl+adVV1Cif1JR
ZKubmUUEafcke49/rAG/LOy5DV6hq3GFLy3MqMXdCjLH1I30vRG5u289a+Cz7y0H
70ClO1Jb1AYIicH4UN1baoPpwcLY4BBirqhZhERpjDRXV8ysStforC/BHCjvNBIY
D/FBIxH00VXExqmsYF815IcFBmAjCpf28u8dMWYbi2gz5US4PfVBZHNXWRcRKN5d
RmIimclgxKBpDlQx78s+DWplAMFOnxS/uxdo9noX6twSmc1xA7q0orowyhWb7GGP
SOErVUJf4pzqZ/rml2lTdk51TMOrmNPRqTuLISH8NfzZe+NRKDnYRJT+9pfPg48y
AXhXoqIgE1ySeRMLG2Mpwlw2omV2X6NVXt15yXRzTmCQNceU11HOw3DVmgKmNMm2
JDoddxwz2S8yNOhf9377XnF03wKheZEBsbfkudHE1osbLWqtWmBANLbj4xxAoc9k
9lLqBaPIqRCAJP8b6JYByAShoXjwsS/TEBQAIfyIYXEUWwJJs13LCwh/jFqEKd0X
zvltbDlI7my/0KS0ZJdsIBruqLUoWD/2PhhIMg09slXatd7aG3Hhp44T7eYaxHvk
T9vdDKt8Q3elpLHwRpGXC98J+tBbwbTI8FeZLBbeLwJXeM1vlY4q6i1sKhdZ0njn
R559hJFFBf7jbLlgUuGtd+Z9Xx0/aJFTwp0ZlvL5HHqfLDsuFkWWImbOap7AUpWZ
C3LZBDnwX83V5t5dTCyFTAOah5vQqwDfWx1VfkSiKuvaKq1WQSml85lxo3eFxygA
l81el28zKEKRqgP7GzmLa/EmcrFEMwfo3nbHT1lb+PNu4wFYAduKMc2YqTQuD9nD
P1G2ymarkqhqsV8GQEJtgvVsAjRPPGccoIAt/LXB5Wn+e5IkYwkZ7qsCpdI6W2vU
3aVA+yMQJTOn4jNRk2OnIEF302sgfUW4VNOGrRR0yCVJF+nh77qRy3oKNTuRLAov
mMUf20vexIJ+XNqbHecwL8lWcEdweBlgaZJFfmyKTyIDxaQ5prWvGsElPC9RM5Zo
66tLMYIQmjf2/5FpszAvtlwKTcTs/Dwz6h58Z+pRRts89CKmWoAD1vo9w3xJGmZC
zC1DFiYQponbOCqjvQZ8dWefIoi8lQNSt6mTLrl3Ac4hW4F88gncjcqjKbs4rINh
ij3MPriD7B8tRtlBCaycpJXHBXRfr5dN+Pry/Ls2mQftNdzngnZ25jV1tM4uEasJ
uy5qJiiHB5+7ZGor4n3mRczzBetbO/mDXtJPAzNpSoJlpcHzLaJdy4WTeqwZnlgE
B/lP8dGwjKdD5aKkUCyfoKcR+SNwX90dpdFb362/5tFyzlu9BcZi5nhQYo0tKCPg
BRQfpLtBOvnvPhxhGHfT6PBVJIMCvRHM5aQNywKLnezSXF2VNm4iDjDvasZpuasS
ixg5ybc6nyivgCsbBsQsxHF+Q8bguE0ammE7IMU+8JT/64rkWoo6smtRxhDTyZ4B
vi6FksG6NJ3n6Y3u1iyJ08GHkvShwu+/vvtONoPFXq400FfEPAT/IbWmejVzWGh8
ctucS5nckryktcl/mUfDXowP7ajQNn7sXPXeDbZmfs7Tve6KvwRjd9frcFZMvRJM
T/KmFqjwBJdyVTrlY0jgC+bfPxuS1v3rJjZkzOKMpw4DjBWi9ayeJ3emzHwXaxdN
nzknWtVoaV1DtilBXKRO5QDckUxr0BMkEDmGQz1+RYxZbKvgVzBplXNi01T9BhBS
b5MbMs96qfUq9a/ImX7F8vrRzXZaCXTDbalOD5d1D7MdUMo4PiZ2pPAa4HbdUKZZ
5Gt42WS6Lq47PsF5WcB9GNPmteSkt+CQIcAttFOwiEjw+u7mjqLzKSiP7zk7Jxk6
kPakHSCbqtKJ8dKGf6DDpw29AJ7XpJwdeq3KmaZkDRo3sHbb81HfJlC+vSvSqRdY
krdcOZ/oOWlckV7iiUwb9eW+QEkRwVbQRAflSRoDwadEwstuN4C0a0PsANmi7zTV
4JuYo8pFWHS+3d4yG0QOccOjeCsvEiFr3a6amxdH2GzsiPPwuLKvhISlI0LnVe93
S+zzpMvpyBLSgm4MXndS+CqKpzkZl/1JXI4uFwE84uAvlhKO9w7a8N3ZFmFIRIWB
BvtUjYIDcK0t5d9oaTgV70DBDwhR31SxVCkD5a61ofuOP/LNPNyidrzVVARvh3er
1GnmQSWtvRTAe9ilFoULTuWOm7M091txivzKrGeYIu4PwjzTiIBa6lU/Oytm/jQP
gMWt1fvi/XP+ArrSA0gVyng+E39cNaxJ4dZkRuW+i3+/M3XexYIbn+cWC+6Ww5xo
dFNJKAcAq68PnrhWR5c1Xg8BxHFHLEf0IgUqAUSJBjomrpMIKnBsPZtY5PKsA2bH
mHaYU66DA7FbC6eLikBU9lt1v4A9oykn1g/KSSK2pA9KQjhYoANp7YAdLDBJftvh
FBhLYJMLAGx5BT7DXiKpYTPe+P34aqYS8OJExUCx/F/oQi4f6MwfiemnUmYuHMz7
Zd+7nCCBBn02joiYrtYMCu6bzTQF94xsXBOMncygtZBLGQppnW2+gY3rfvwaRdR5
mwbql+ZROpgZmfb6gqOr2WQnd7IUxb3Ci7VHmL7Tpt3MPmhYw8yy/Yd3U8X/q4X3
CA2E+DrN70hkY4LxJoBF+wp0gztUItUHnyp8H2yOcCjnKA/F5Rg+HBmITNvXoSFw
5uXT1XGfgLJHgr9xzf81hCkQ3ZQ9J7IC9PxwGGPYEkQCFEdYs6cpypWHIPUWIFOJ
3I/ISsjHOB4zyekQH3iDuYgL0tW8JPGSRBGHkuX6PQNQ/kp07QnL8zEOKfdVlP0m
qs93flvuUxvOnSOLwIyZpkjWzrpU9/9oEvYzRiUEwdwfL/bgWlFVBinaTOQie/cl
nSj8NCVfjhrRZ5cO0JLOGCS1vg7qgTtpwnHueRYKJhCCimkFvqj6ojvV2jyvxaqt
SDXsaxYRq2Z2YZ9ZrXMtn5+N7ZH2QQA/O6oU+3jjmJjdkXVcy0TYBSaxZyF9uuBX
LGypZoqoW38kV9BofaBZRyrCjHTYfkEyRT+q0YJkolkoJ6SQynhgNeCo74+fDoJ4
Mdyv+/XcQekUJfZT//qF5Nk4M+t5iTozL4MzMce0uc0Ox2Gfj2Yg7gos5/MoG0cA
Ekx3mJc09wIhyNRVMqup+ICrqvJf4aTTU3Q63UDUlNyaYAJN16O+n0a97hoo1z+V
xGU89Lk2z/gm9ySM6DyvHmp/a8xoif2xHS2ZUq0mhdMcR3V84MxASSanz1iM6QVw
xM9vGypBm0HsoVpP0Tc24ZV9wj192Ytwv+bpiOPFCuEkJbmsU2CbP9b/WId+v3kb
I08CzqB3KfvjrWMJSMCcGZXrloaYGKJNehd8Wn6IX5rJQx5JvAEpsEoElOEynD/1
pUXIyJvUP8E7SCg6xJNBFBDLrUUAti2bsaSG3WQfvBm6abXn7ol7+1/lbBM2OoPZ
z19PmWfu2bkt+iH0wRpV7f5ASTdKrAdv1F0nX+o6sFtMq1VdnKESXcIh9hW1F35k
h8GGQmu9rzUjvh4+6plW2OHgG5Ezop5XxvgWYB4vTBINovTAfbrXhAYiaZtnjdfL
tTmXnJNzUptEd6J6AIBHW1AU3EQeVHe3TbC1Nbv2ccbodwf9AnXo1srbXl//h5cz
YqfoDVSo6rHJZj6VsPkPnXTLMnCAY2hXbW29+meYFouJh3dc2N2ckICtm0vHjdgv
pCkEZB9qL3+6h5p7Pyhu1wgENHFxgPTTn/Xnooa6BzZnQo6+yqBzVpZfN6tWtbhn
9ehauiBB6AnQV4x1qvE30B9VwLuqDOpEjZWq2j9ZouKkLDUJnp/fJE2fV4NO8x8D
fghHJvfWNAQrMUDrBHmO2O4DNQPdy86UsCCNyw8XEwJ+WNJDhp9h6AwS9LzrHa00
MrPefwYVrSwwT8m/hOYzl8ApkixtSZnO2q0Dm/yf6DJTCheaTtaGu/mJX6buLgHy
cWkNmcGXvJrAJjh1YZLpSvqbeobxaQJhvLcs8LoyVdsDIGi5r4cyG1HRKgkVcBM9
W+IYAV/NjjwOKJSP2EX6igs8SbSsljRDCkPERaN9bvstd5GGvGga1qPBEq3Q2Sbi
hDh9zTdh7r/kPmZUPZ4NooDZfOvymc0KDRX4Vlx8f8Gp2ewodliZcwLtE5vGtYvd
ENb1RmUhbYYtHLl53YNyV2wgcjpwh7qsg3kgkbKfx7YjyuL7LsGaPc3REm7h+aQa
o2sP3izpzWtT7ixK3aNNCePEgcGdGjr+jnJoIi3F1QA3tHFY/IWaZ+FbSUTVe1be
nV6vSwkL196eZM/+Q7An5CHtpHswG2LcEE+KgM+b1vmisYv6+M91sE1eT1dBJQw6
XrZXe6vIhL1OAHTQJAw2al9YZQtc/ahNyFkdeMi/pMBANYqycsleq04Vx5Ieez0M
axCwy3yk3OA2wWskSaB4EYAKwSX0bI+3DKsqjoaKw07i31NA5UGjCiALfuWPh/Ay
wyHqe3KjBQkN9RjWdlLPc2BTeoDzIGZS+AupJqRJX43uFNGLL6JPSaw91NdiSxjj
AbuBD41jeIC2x4IQHgaAKB17Vx6yZwv9ibEPdStcAs0o4wPR8K6+vPtldJnJQJ4g
xWsWxqgQNEImVtC2sO8jAolKJKiHPJPFiza9Fv5aIFC5zay22UI4BrruFseevGSE
W3o6gmxdGvf5FJ24YlbGYbp2wFfNqSL1ZfToIyYlELFuaktfuah1huXisLdajZGu
xT6nrN1sMEciFHqI5MJgtI1Ea5E4d+jRSGi09L7ywr1M28u5wCBzucsRluvRCZMF
ApvKEEoVJFYrEbecSp2LNMZQjGzd3eifJGzGtoQ+2cKRcuLc0VVkajP7PaXRpMwx
tN2gyPzPG0P/XhaFXBZA1hMGV3dQl2ZXv8TPBeUi42spL2UYy0cP5fP/wOVzIQvN
KiOIvQLcFVp7WkVmwoWsC4O9mYlhcBgdUJZ5Vh1ah7XcUOy7/6fDSnp81QYS46FB
hIHMR+M0WjeLxIyF+Y/oVXb2YsMMw1rnDF+j/TpBp5PHecfhl/WnKonT1hyLJ+fs
k5RRL4iPknGqrRTpruJqxMcr+URZCGK0K3K9g5gbFAEbP0g4At2msxqpFYv6gP0q
LPiNmVgWRuZud2QK5PEetKVvWElyD4D24ayJ/EgQu7N+bNi+IPLMMVX0kJgXUE3G
QLnapgGPcByNfV87X2ykDBOknQWza5TfTSEz5KgU1qcd15nUNe8ThYTv0dhHnNCV
/v+EvYMU4kLcc3KJsbRO7YrH0mtTDbkhJiZ1j3aUh2XixOCo7WpQK25WdiVrox76
7PGccR85Ly22MYI9eSqHq6OafwE1vtjo0LKXcORlRHG8jFI16iWMVa3B86od0qpb
nysSE01sttZGe2DqHQeUb7AovbCkiYAGaGnmUww67YvbzFj0FF7QenfXb37knBYD
SIi7oU+afRTiot7PKJlG4WwCphe9cFHXjVjOqWQdAC3fTVVPApyUMnPPfCwgYsEp
6wlwVwTdutkArYUBjSmXlEczTpN3l8nFItYTwqBkGxx70klEOVgYLLpyddzrbciN
mVGlC8/kTFxE6bUiROuSg2Sw9WvHVx+rJmI8OwpQVyhPSGQk+vA4FNGkDjV2bnn/
6T0ZuDN/C7a/r9u8zkWaKx0VwKNf1+d+fp4YfuJwVlH2U4YR0pAhzWo2FrQRwB5q
FowwDzNxmi9+FWQnokDO/kNl7+rOVKL7e1HNxLOHj25UMtOg66Op2QBqkmm3RVH+
mCzvc6ZKuFAemxYP04RufrjEURf1tJ/BTqmszKd996F/ozrQhc3hwp0C0quExfsU
jAIBECqHEOp4NlNh/YbYzPh0yjcFI5UxFTbW1AshTd9WIhLQ83cX5eWFZAfsSXpe
HEu/tpl47ZMpsTewkg6IAQed4i8/5pNLhwCH3X9scV1gqyGOd0n7kdgfktA2xFLc
VpviNP0MBDl9lXvspAG4YDMlHT6ouwKR7+/l+DaS17CMBOYaCMMZWTQteDK6u4vS
V58iPKGmtrm2TyVE2XXA8th+/2KFI8BVmIQCU2CPP+b+3ILJtBIpStNw23YTm1tX
Pyy9WgAlpkD2XkxKzf0PUJ0yF5w7Jb288gs2EiuHHbTsiTRdRgjIe5EV9tfVPYGz
MeA/rcmZYm5y2V7xvEPsrtELZMDbfwLua/MvjYNia6wP2ypM4LcBkTAhA+z6kSM7
MKJbTP/qiKOV03SggxwgIvLLUXMDA19JyxfAc8q/UnGtsrP4SvplXbQwfvdXnh2g
BAV56BqKlU6bgQ1wsUxu+Po34GWTsX5mLDU0UMHkOOa/7K2wKWWC5GMCdBbroEBR
ySySmsKkwmor+n0ACWhuMxt4NpGLES6qo95Uuq1Y8Tp7zundf5pTGuOcU7D84fgs
3fOoPS1HYM9t5vH85f911anG+wf00nt9Go2CS+9KV6vQwtTcXMla44XiAxeEYN4H
C6dgRILsX8R0tmxYLnew+O2NzfZN6pEQxn9+41+PVcCfdZraVY2eIXP6h5ogNemP
l4yy+vHbPIszzBJ3Tw2nYMyvO2O9quO+i83qNPSwScgohPc9HP79wTUf4irUnXRY
zB5jlVDo9qGWItt/OzMC/JgaHR2fX1bpdDwrNYZDoE1lKOyznMF7jGB2yvbtznjv
YwX4AFZmvaPeg7+vooVVpJRv0HMQxKqRwDhn/81xe9NzdEumx0Kjlz1JVi5IMYFO
dyBvjkn4RBg9SSkdtjV2zBoC3OrkModd6h7HixUKWiK4C4etdGVxSAsGNkI6+siF
Sal74mSHSOtUTa7MjuF5zkjwXuUqYYkQZ95kj0v1/WJhtR/PAG0oQVpO9gBaMo2b
5/4IEesA+S1jGxu17U9/LLbPDByvLmMyMBYs7+dgbc4XmjMsCH8CPTfO5q87ayLX
St5TToqk4OuY0fLs5IO4nz4+0+UG0YndzZ34H5BWDPBLxKD7wgGInCYG7jxwHt2K
EyGG490JFBUbsC7J1LZWJtBEWFCn7aywJi+5ykx9HQTvw9ZiIxmm4I20iPzYISOv
+CZgmg/oN5GQ15EwD8z++ZhItNw+gJDV4LYOcUI/R9pndDLzLBZdiOLjLDIXvIHV
hwcLICsSbD1eJJ5miJAIUII2HD9dMUOivC36FwrwQjDYlHIoe2H7Vr7YWHQMU4B5
LVruWLdpGu1ZorT/uxNGnzBpF/zhK4J0gUYtIMlVzenVW1zvJ7Glx2bqa6ztbdj4
icDfax1wMFqgf/MKmEPQJEPSAnObvsConwnPZzpkIw1qJJ/te62f2IGULAu6lqhf
KU0yJN4B2S9hbWl7qfWYeGVeAcPfAfL6/sOacycW8ECpI2nUQ9MFEIWn6qUK3qe3
deFGF+5wQcuGrdM28fIm6FFcGZh0QhcpZ+DlXjv3dxck7Nj8u20adhNCaRk5QbAk
ENkDEP8Bbxgf0xc2K0Sz9h11I+cFn902A9E6337N0t8VsEx9udehy69RJqpqnHlu
u9IwwuJJVTYkQhN3BX9XW+HAKVNkAoVjxwVLtO4nVPwhIwdvkwtt0pFmbjl08CXe
MejvEgvG3W8kb5+QsDo5w70MEq2F+9g/AYx2xP1sVCPvUqcHF3hJnkuce+0TsKko
ycglBYM9m1rfPH/cq+Z5bXVXjwkLWTYkMYRh119RENKa3rzkaV6Vsu8wfjUIZAP6
9qmLCQCNRWE944upF8KmqF7y59RoYXBY3qC1+qLrQRWkUy5N/uxgA4F2dKn2xGTq
jwLDhE20yjnSqeuhktmG5f4VuuX75sImyEcHtJafxPB7+Z26Hs3hnZZaRrtys30r
TlPrVGiPUBBkiwEfkAXZ4yMTUO7tVzGrGSodA+EAd2AG8HCsZgoyVu+uJsbfveER
GdPSgKZMmDqgr9KCoBKCoGW+JfvYcGgYyAZtwZcPMnbVdBwirmTuZGXkOlkphdgL
WXoUzQPagWI6i+2Vgg6gQB1xJEXSvMRZRr2QOki9QQKXedHlgBQbrtJtkqTjGkki
s0LkeMh+54jjBKVUnPiJ56al9JCqrUFYTAB7KRvR5yGB0QWkgfNap7Vp//JcZs0d
bFAvcc7xKB34Qp70qyNrVlbKBCwxBNYFutBN+SZY7lq0vbh9X5nZR2Vz3nxz807i
zk+8DxG7GZlKg5fYnZvJByGOgBJYaQzSOvLyptPHSL4CLmZMuhrPfueP0DmumxMm
EFsu289NS+vWf6D4ja/QhVpmXlPUgLlDCLdq9919wUEM1s5ewcuQIaOzPMhC2bjl
Z2n38GlEHtckth3HKFKsgQzpuWKw55KaHHF7T36NskuI4qnbccVWmkNPyDQerLfz
LaRlclB3KYCUr2j9X+PS7ZK8VcSzxah32ikIN4VFL25VZoK4cBBvrChFCy/HsgIt
MWSBWXk2VagvZlkAtK3UDOy4S8OMXCQhTCre6ZYYDmdEe21sCisZyZiC4ObXt8Yo
dSNNJgDt7UyDQ4MPrTHPrIngJ7LvNNfeUOuinbKkK9P6jjT1I2ikH5tuqtxsUPQF
oJIlIUf4ie2Wg4ItjfRcQr98ZSvz9qDEY8zFa9SBkmXXD7/wBXpzyj47l+Vwpf/o
wF6b9UXltvjq4lxzK43qZQgWnstgFIxHmgZU1/G5D1HhhbmUGZF6q/YkjaR/6uW4
WvS1XyMujVnWviScgVfDRiWGvgb2BsSqluMecYbmZ+6E3jFN5MKZhU3ZrScq31W0
ecbTVLavV6XgKl+U49s/p8KA30ER8Nil3DjR/Mk4FAbwJJEJ9zFKCA0lu66WKcpJ
nsfTUquJgA2ml73GO5xx4kzCaDE2IwbI53OpZRDf3td61qSFnx4NWwgM9QeXVZz4
H1KB6YpbuQFxzfYTdP12c6L9YyuW+3ccvM9BTRUZxDsXdRDqJlLl+JxJPtVpUTD5
6qt684kY/xD3xhRtK9dem5UlnRYiJz3wCtPLvCVSgJbyniFvWXEX1FAArUjaainE
2XhLPm36/g8O5YYWla397DsCW4uL/y8cFE2dgjZyads9foG72ntVaQ2nthqFF11K
rqIvAITMyeqoDEG7Y8kdiQSnTC6Ofmxq+5FHWTolR6vkrxHWVm6jibBn+dg62hgN
U0HEDhqFWr9PzXXKHZfYxPuBJYSFde2ex1Pia3z+PfOSZSG+BaDlbLRJ5evQV8WV
hl6oDmgfdx/kOglHhLHcaSbykzEmyoY8j8OeKpH+PYE/mCBtXm30kJyCPb0qZH8m
dxg/w00FbgzGOYK3yxrPFJjMp70Gk15uKgrmcovIC3LgM/uN0s9+F8jytKMOC74+
86YBFrCEOniQSIQrjVtfA0WsRXYITirCR35YDr9vmEWqhkcho0miHL46SYlsV2k6
Rs7dN8xyVYWhgYrsl73x/VyJZMbXNAKWhh+OYoBEiK4TtvAMSpv3Va5Ak4dekFUv
4gzMGfSNJ+cVjOyXRsdFjxHq417fKvM2q44tS3XxpU1wup39+WPdx6hB2oXH3C3o
au7Y+RQc6nfXNws9QS69xsRfxSPPJIlaD1zDPHtQRpP1A+4gBsYFt1CwuCEz4H8W
NG1H3Kls3/D2d2pbeXPm+ywvkCPLTiQBJ6QrMOCKAObwPxNLCzG61uBKsiAN6ecH
AZmCc1xPMgVGC5ys0AHes1uE5tFW+GTqLlHHO/esl4sSAt25sBktyLbIEwkMgkby
aYezg0ddSxZK95ReDHYFoGHrPJn9Jt1IHBfCT/JeGxTq4o7IraskUKF8j1f/tPbZ
OtuMBRe+ukExd2Kb0HDNkLrpjLWfDovrYNf4b1n5s4H3fncsNiCIaVmacvNliOyi
fv7gH4pQ7I6SQQuQJZPxdR3b0sNuU8m4rLNQEkEI2QTlVhKbLKsTS/YJkW6jA4Wa
R6LVOXY0KqcdF0AJCbqVGOIYYcSYMeplXE+UEQyETDQDn2uOvpwhJbkL80YEOH9b
JjAdQBMjzKbOCSwqKu+vXUR/TllDI/9P1U/lX1W7c1def+PaZr0hj/+MCR11+nPI
oLER4sYKPD16YQ8Wm5iozVFqUYTQ3qRAr/T/OH0xNkNEZJBKPeA6tCiDi96cYdG+
ZS28FImD8OeKWVkgj/0ldDtzxDEg9FMoWcVngjgLldnC6a5QKkFeiN2fC36jXjGZ
LjkJ6pja+ePOnZatPlk7gcei0L49Z4rDAZWmydZTL3je1m+NWDobd60k5/YdZRok
oTADNs5c0I91FwKCeox7eMoC1XkIIPcveJxYR6j4pi5/SHvmYHW8UD0PWMXeuSx8
a2ZyxShu5iPiG+wHTchbC+zfDkJdVlom2SeU8hyqhEL27X0jjdRzARDlzXeRn+6S
YfYbF1l16ZP2IPieUbH6gjIE2cbcml63DetwMWKQJvOT1/mo+gHlP+0sMFzHaNoi
ZsLaobYW28g9pQes3pB7c5m5Eo7XrsbGBxtZ2p+WJ6+azuWIx6iZ1wkueHEIY87O
8e7mIY6gSbn6c62FY8Yp3i51KShsFReeLeNOZ0ZiZy9uEZoJuOJl2ayk6w9dGtIk
aDN5FIA1CnbsTkCPSrVVj7mc3udGgxTCmLp6cJGXXvbdNKA7NtU6WgIKwylzREQ+
WSCmz6JPF84ukT5h5zwqThwF9/iKmuqCMK6gIOuslHK8BHCBY294E1bbTq9bDtcj
n+nn9qLv7HlFK3X/8ZTg0DQYj8yrjd+00mMSwAy4GUq28SWwlF8S9sHOTEkX1xN4
fAzLFrmyI483sL0f4FaGJDqFeso65V9FEXa3tXsSNUnqa/YOLeywHK1zMagx3an9
v149RZX5I9eXqr+Hk94UuYIOXGBhxXfMp3Syhz/iTGRo/ySRR6r8Y9rnTbTRoGzq
1mDMOi5SKe4gL+yCDMElwP2gEcb4MsxrhaebszC+CxG+wlk/ZKYkuDW9NnPp6SQh
TqSQ1n1mTjKgRUbqIruwfO4zPw6TCeA+U6Dt/C9yu0NFJNgogUchkm1pfmW8d9yn
kA/UC5RgonqUYw36T2wYK6Xrv97nH8r5pzJGuOft1QORwLuexwZ2qlPQEk1GE3Uc
k8RpY7Qun7cXiVHycYa/XlqXt2SjNNq+RD5z+wUXJZRoWPdvaczMLSQruLjbKF4O
6QEKGg7kUWaNuhzZ2ByNW8PKYwPOLqVhZi/WzXb8FmYfT/I/wkHXZk1uCqMjayCq
w1StQc/j4RSsc6nxAuzhagNr2AQxRxUxFCfuVBI9ylfp65keL5G5Ci+vbKpzllvp
WtRLAq0LC93XuqxEfeHH95RMXzL9fQzBVGQpdUBCr8RIUd8x0rMnXgfreg2M5+oi
Rz8jtFcqIhDwqo8lbnSL8W0o6SE6I83IecvpwIyzW9DB+0dDJKk85gvHcwvGukpp
6DX49cOnjGjiV6doDZ9HBw0d0Rlrr75Wb8WbUQi44Uo3/Y5mrlmG8wpceSDw1Cjl
LFPMI2mMeoiybQRUBOzVJRFxk30dBxW5ILXkSP9z9VCj0bCHGiswpkJRt1j6Y+wv
esW6PQAOfjVw7h+dbdkAkxuZ+1Yx1Zx4bZ7TaC4NOSp8QKoroxO+b5WpkEQ1vfTV
zwZP1IF2azOGrlSWXGI08W/Onu+ABcJSZ+7yw5s5uA5yV0fK58jkgzZ1mX64smdC
TbLaqtOBPzv1f7XNtHnVsvSUxW/7Ygkl9FzNFEitSlYrfAFUh7mo8ybikoSgUrb6
K69xZS6J4gS/ixK5K+zIbUYVgReOkISW+VYk7QBz3BGLQCnsYs8da+q0bty8+Grv
mTPrNaAusAVdHJyL/sMC1tTh3ENnww8s0AVEjxWlnw8WlrU20bEQudq/JOcXEyUv
5+Ec/+cbhvYe0lR2qiejmupcm9mDHfJJnHx5UlN1Emq2oW9JzxK0FsODQRYIjHaA
3cX3urw+qEJP1Cn/0DTk6eg4Njl7Iy5A7rhLbR/qP6Kc+5fEYyjtcha/mCfH+cHI
ISFFV1F7+iLlZDPRyt+oaigoZnA6yXjUcixkVMuMY+QhxQ4hZOykNPFLKDpKyTRv
F3Mf5SBt/W6+tdqDI9zqsSQ42Wm8D27cMvYrj+voSYknACP39PesjKjo733mc9sR
PpLEDiUCNpN0k1rs7UaxspRbIGEEoiOLemZ4chjD/gJ+zf8wRohWyaLa/ESTwzj/
0N3LVduJrVIS5hAv9ITo+ZXO4j2G2Dr21vvOK2ZN/or3N6Pg1GXkm2j1nd9LGpPd
rEP9xO6sVaNmgohathbkLjYsZqAJ9Pe08rRbmB7/O44U5imxCVoJt71O30PNpXDb
VuIIJcSmneSQMSLD+fcTy7H514ybd6X6139i3XOWlPFdEjnpv0lMeQyPvRBLnJ1w
ENB/wCS0UtO8ShR6pdm2T8rW7AvuE5b6Bjl4AE2v/nVuHh5u802c3Yed2TDX0HYg
Kmac9/SK05sjRISBHsFAuz8AUdwJZY9fe9ASv8K1najX/GxC01gtRVFYh0ZqcpWH
Qw4Lpf7DEYcaP+CW27e/ds3spwd8D2hFXaEaiDiVsoxZE0jxUP13O6U1auvY9nT+
u3vX3EUZskzuxEevD83AKH45/Kd6uEUml8A71XxOAOy3FHhfBUIvfg7CGYbmeyvm
ToXXn+FjlBy9fUSab8n8cgcFCuSJYjdcvdQB5uEU+4GBmPVp+LV7euV6yuuahpzj
mdeDbDQlKjTgYzL8LuXcgH7t4IA6GnEfpEKoAzRThfYxvYSPgEazQl3Fd0SNdfDX
jyC33D1pSjO13Vu4C/FYh3xInjNuV4mDx2JuTpaqQUPoIqTrLE3VZNsWuCxV4MxK
PSyQ8KiFIbyzCAdcBrbblgrD0HVu9IxUUS4roRAgXhiuhXjXgWlqIiB5ESX8ez3o
fbiEwDPR9BPbhNIPIxXsa8Kg3jRGfoptL/+Vj25r5qI/1r1DNjDaRlJJ+i9YH37i
t9/sF25mvMHZ7WJCH+U9biXG7CbuIez1R5I7NybOOB/FjMRnd6VbTxoGxNk0CPGr
KG+0Gu0ipp1IKpr+iWHaWWCLvPmveyxRZ9SH5WG9OabjFi/sgn2MUv2zeyZdbLNS
4VjvOZ5w3fx27w4EKedxzRnXTtg6so8SNGjlRwbvdYkZZkMUUYwuQn+9bpXtlZh1
odhDXFw6jzajw1ZMFAKuuFTLZqA7EbSNIpfsv0cu+Xxrl+M8kosTswdi6Il6ow32
DQ/4SzMG67wYsnPZqD3IH7IuYfRQFJF2yq2njoHXtasx674q+p8lSA+xo/y+8zTO
WivrN9sC5cabLXy1D9J0vVjg8c7iObq/XEMNGx2z/kIc3xTT/ciL33LjmlXbZ485
mm/HeE0W0Q4+XxDsp909PFQ0Ny3khxRGSrW84Ufs9++iofDGXBj3AEo+dfW+kQx7
AsICvZHMds48JPvvJgQdSA0JbQAtLB46n0jiDaS6B92HGdhcBlUppS0Qcejs7V6O
jicpHdILEe9aA1Tp9ShsdTMw9MFhI+vyuPN1UJQWzBULs59LV22PBKlMLv5P1MvI
77y2tLyzWPERyUsy5SBUDUVmCoPxhsGiA8bawKJ9My5hKL6tSCtClIfsrIgjSEkV
RC00F5alZ3IAIVSghbwjZDq1V9LwPmsX6arEpYqgfdIK71RHSonQv+ErNy0HZShN
njR/KzaXbRUkA5NUM4DgcJZpvfTr2IRZrNd+HQg64yZHo0DJayV+XVhvAlrqXB9J
5mqhVkbXkYvaBBv3+NEHXts37Ec54evH37PRvswtyJXwlMcQm2jPsK/bb7GVfr89
K08iAMECqaKUR8DWOdjE+f2JRQsa5ACETyBPVMFbF/S67OrocenyAmcpyU6yWlYo
hggeyLS7SHGj1fRtb6BHm6115V8+RRhcGiDrMTcUT/7szpKGLl9Qps1wjK93WYbB
SoK2zV+rvWhGdLoLt7+UjCEnYo++DObvH523EGdfZrsf2rC0xIKJq2qBMNgy6FUS
QIk/Oht4Aw4aNRFy355prPfIyeW8KXnJYft/v4NtcohhoqCDZRP0L3HVmOxIU8dp
joLEzrDERos0x9TTBtMrle2SSGhMvgLdQVW4z2WGfR9bsCmxOmnzNXZHm/GhWYV9
pTES+4HYkennLWbOF2xvv/qARC26AXhHEJpcL3q97D/m5/fHx1G0gVeq3Nc8NKWn
j0wjvbSIsmvWh3XRZzfQdLynxoRqqtw2pkuUxPJYmQDG0t/yaHOaylNylJseSQKr
5iPMssIIBCAkfudnqiLLnblKkMbJQ+zHLc5kzAhJmTECzK3yu1fjQLXMScQiSC8h
sgbBeWCPKipsHk9TI47ejczx5sXiQqIugiGzm/QYOf2OKsd+fBvO68JCtckdlk70
sAFYhylePgb/rx4ennDq0sy/7NP9KZQhase/EU2PZwUu358JKXJ/oZ/1SlIO/xxd
4bM/SGYC3IkggzE0S5jx2r5sg5A0bE3RzgV3iIfBbGpNezQkKMvnGmoTT7ZqpQGD
O96i5Bz6gDzgfEbRv6hudh064KTS4rhyH3+oTovs6LxqTBRlng7FshioqAejf8zv
tyEUNQG5gOLYMJ+IkJB2emmEpIqp+/wI2+AVkhzYJoBUeIM2f7f5VJCA6Sd1f5Li
Xix1bRBbutJitC0Mqm3chfRKdxdlY4xuC6S5yEC3LfYJeHpbyd94ZcIV05fQ0Tga
S8JCOhNli1mXzthZvK9cQZo8VBChTpolwt6uK206aR2atleJj2emPh2fH6EWkn2x
JvvNPTkB0GyzUfF/PeDRoNqB3QtiCSJE7+uKHz9zoICRkYXUddbiUrCvlc0yKQAj
rJPTeMElCQW928yBuQQJTDzKmPGteZEe4VZ0T4MPhKRSxWP6tLcanIXhivqs/le7
U0fhEJ34eqzOFgOhpPjR+8VdwcaAlCSHamBz0F9EJlSi0EuYZSyvVPSUXQxKXVcM
6iT8Y2X+uewsWByQ0JmNMLf6iPFnsUmo3hsb48SkJ0k4OabtN1ts+HvJIuHaN2id
nT3PcTdoQzbFzNaSsva3LiY7rjowKRnEC6SY7deDhW1AptBEh5TPdWEzdgTqxO5W
bl1McXLyBcmUk3CUH/EecXAPeMSfkKGZRsz1SklPzmOQG511KjnlsuTWVjHeo51I
jmDk5nogke9pw2HnUu6RcnJIkgriGGsw1FQvZUC1QieClQBMutTte06I+X4T8TWs
Eugxolaj5+g1v1cJe79wyUpsJlvtOT99L+JuxMhoDv0XmtLGrM/UW08Hv23pTH0a
5iqmsYKMYBxdOeSyETDmwqGx9uf0u1gYcJunGhFy3jSNC1rgXK3FoMwyvi9uEWRT
Jby1xwNRIBeVLzF/rYLK3dv+zIwdcrp/epXxEISpab2Ie6c0r8jWcUHusrpYZTRb
OytOVmOV5sug2A+c/YS3tLK0XhB3eS3EFEEmeZ1++DDbXHyv3Br4+ST4RlU8PAZ9
hdtmY6hU2XjJmKXS21G9zfZinn2IQy5YOys31/ijGJNg+oOwUVS/1O+lXP8VTgP8
ugH9EF8++OoTuW/t4CwXylTjR9WX9d9eiPRIyWcESr9UMXgpFeFrdKHEIBgYmaE/
9ATlEl/wOxLPjJJR3uFu1TGkKPv/R8de9fWUiLtHhScJcnYy1s+ZRXJwBFNlVXLF
t7X9c+u3l62H4WdA4eW2+FbwdBHh+/c6h29AeWSGSyjsW6VWVxerKEO6C4Rqye0x
ZaZgl/3MQhhCFMedtPgFmWsqGtqXt9/re+62wE8ba3b3kqqDdBEBG+cknvHj/nrt
O9J02oc3+e/zwA2eq/fp7hx4uI5o6OryN5fucS3tj4t9ZhAwActa5AOhSq9pRZVM
xhRtUw53TD2L6c6DPTtWSpSf6aDHTj4A4z/1Qg4IiCnS1KC9otmNj89xe56RgzCt
5ojeEJuk1SEDhXk2TJDkOP4+LwDQHWOw44mYItvzUZHYRTZRlBRZlpa2V1fZSRf6
W+ObUwl+Ptwm2CIx7c4wFJyUa9hHFMWiRBIUxYqY9cI8gFa0EfiF80tXjykIVWpS
pdURYJrrKP0/HHkxwPmdbfGTxkdkd8K8SLughC/0a9yN+2gYuIoTkk1GmPwtkTiA
a5UimiMeWnPNYXqPjR/si/vD3xUl7dTgjn3pDoOvKJcYtppfS0HvJ63vSIzIGcMQ
IKmTJ52vgC/cXVUXpVKj+Xd2nGXlbQQWBZYXk4hanlPVTHUNrUs223j6UyjGCGYe
Hk3rGQn0PFvUwmrtG/VI3LISnTPz3lzBkGVOgObmIn8a31Yib6Fd2gJF2cuISjwt
Z6rFw+FzUd2XFYm6oI3KxAQ1br5Hj1RHC1N/QcocRw8appTWmnoNe1WFkCxaWF3/
7Dk+Vm3rJ7kDdLRopTLAOERFUcGKRAuZlJ4UD+TUvVTjSrPkYKAbU9LXW3gsa1L3
HURN1AQBOVocR8wjr3DpiL+9mEne2prLn3+LyTAoDR//kvQEjtp9OOeOlVaNNPSt
M8vE+G2Lp6qyngi0CRgz99aPppcOKW376wTGpBWdcx4F+SdiBcU3Haj1RKjZycPX
q4Bj81+5IpeYn0zrGHqhZYRAS8xfR4iwFZozGRbs7z82PRggHF/Hnu51O943bImz
TTB/3DDAWUH/FVKq69NH17M2H9HYPRT2Mmr6bisOmJMy+iKpJmOIsG3T921/HfZI
EaUrzqJvwZpFyF11UPzgVBtvp3gD5ZdvoyUPzY1uQ/ZIiOH+MXySRwcY8mhxc5/x
3r0/u7DejqwJekAi4YQhJW3wnmxH3qPLtmcf0WnzqSiO8FEF/yTFC6M1bzzlZ8iv
azNzYk7x9peZ3oUHdv1bOPDzKQt9MWzYkfO75NmdWUz/NKeT/ZIBEHJLIHPMgoWl
Ro52UR8GWsI1v335WLxeFElSYGx+0glsegkQ6ykXvPtQzjfkXnj7keJstJuImW25
QS4YyEQ5GKMqNoGgVSMCcNzuhPzNyDJStOAd7Jmu9zwuo1WdM6o892amJdhx0/6Y
U4RxMG/eRNbdPCanA4pgAQPVJk/Z7FvRarlm2Wy6/RG2yVwMkWryh4E4nZkgoI4S
ATGyzXrE0GRsMW4BjDLZId/cs+vB7co10WisyzCx/dO5RjCB00UV8Eo9bL4eboOD
TRqIcKl8xmkMjNU41Eo8nzLj1cT9d6toqhZvqZqms6+dT+FZ5h08145aBXoqyP9X
Ez3KtXYyS5k06EVr229TfcXoDgTRu1HkIonmLeo0kh1MzEIQPjtr974cFfP9OL0Y
yTnII4kyIKDOh/8st+xHMgaHJApKIPTK1j5v+oKH+QTwS7VbtxfBtxVwRghQFsbn
fD43R9/2jcWlww4rHK64JibTR9+67wLgP13IJTkAhVgT7VZABk9IeJ4SNKxHC6Vi
VAOwTdFZogsLGdUgaJmxAz4bNWGCgH8XpK/hI4adfw54i1WPu9Ix3+nSsIzsw0hV
B8bI1GkehuhzDShotdIfb2yOnXCad9m0Tbt/+vKj/dibPeZSfmhg6/2aQjsC81xX
0OXiL6jZGXKp8b5p9B0LWyjGZUwo9Z1tu9mTNnGx5LirYLW+OW3J8Hne0LLc+3Zf
Wsabfym6PP6JwMoiAD4ScKV++AvZbw7Ys6OwaoFgAkRmFc1sFZFEZhgrPpx9hShD
XrLTsA4AXWg0ItJT/9FC1C42k8Ps0lDirbHtHYY1nUAUWxhzynIF2TaBkv4l5J0p
+87ScYFnEqz4Ply14Ap2WiviPce4czOQJbra2oCuvlQ45f/KH0Uorn/1sLYrEsc6
ghPyxH5pOWgmRTBqIbRkoKK2dhdqQaXdXfmu90tvJVAEnCbd7QMmjgxXHn5EzpJf
Jh+gGxKosd8NKjuBciQ1P8mt9CtLs1r11qm0MtusA0nec2yuSHDGiKYS+iQcbI9z
9lQ+n+iEFG5CcDz7W/5W3S6+L0K5Xf95C6705T72PpRsJjObtHa5ba7mJvpGbRI6
1qXRhP9WhYR6496b3UWL5eFou+xwmu2UTe2c3Ok27uAD/AMi17gx26BSK2qe6xyW
DMC+yr7pNiiCEcPhWb1NECf0tuQDcWtFRIyNd1D7ymGo6TCSmRy7lX3n9V3K7vlx
spIEhcu2SfNyR1fNDSXB9+KEFvJuUav6kTd1T9as8HFip0BjVPc7WyHQikfIJyw+
qHd/vWdtTKIhFD0SHViZHR7wxJyNhfblMyt5jFyh7yhJc7VEV0u/xbHpJliZ1d7c
uUwKAqASaU6BRDZjOhFgT2OOjrx5FM56bqz1JeORpOErqJ7laZqv/3IE+dJR49Mv
dIw56ImF/qF0dxuQmu6fcsRNLxZX+dKfsT5fyZ3VhUfomWZU7P9qjsycGH+6oKKb
lw05v1kPa1tWwm6xi2yY4lEXnlNGYok240sJ8dQGjZoc4rA88VSA5XaLcizV0v5g
FXoKoDuBxjehGJ9Ukr/2f4DrNdL0hyK749+d0mvdY26atLodq9q7lyfSzWhLHo1j
YBjk6KFCcIdcDrlIuR3rBVlQMVgwTXnfbaML6mEzpDqz8doyI2OPMElhDNVbEn1z
mqcvW1rCJpHNojuJubHOc3SViVJ1xB/QkUhEWxTEDkiN9vh4bXZtd7kszzgyiUJF
RskHfOn102JRUmcrvIzuFYgHSLLh940Vrtpy7Z2bPcaGclR1Z1/qiI+iqIfSjv0P
c9HzO4/zNB9CPEeU/tRj+mLELwvzoNK01BakCL6FhLcGbV6owCljFpp4Ad1g/DEg
KyuDMy776kW3ya9w/0cFq5Sa+lHWUWnHqMwV6SuEzY8ALhUSHtJIMS5cSxHVwMCX
9QSjKvK0xQkOH7yZ5NnX89NGsMUeYCeijUQAUw/QuTRTGrg2GXrNG/zvocMLLv2b
k4KgFbYYVFCPCfWtFuVOgzQdmlsV/yEIt3y4+bsUVDsiHncy+zv4ygAk77yhtq0s
Yn7lv+VrGpdL0YXMi+xyDpwrdc/erUGt3XGFfm2be3maCTOU3ExpITOpaNu3WbBf
mLIYQmorY/sFpBA0Tjd8l1nQ0TMaMYasUC+dCKDfTGRVknR/vrbynlI/GWX4qjvl
tcHa/vzY+/C0Jk81nqbtPV+ouTFIleqTU40Nw90lr1FUwapOuWLQvC0lKUCwgC+b
G0YjjMUM7sfbpQm6cIYqO4tDghI3NYr/TQgIlJ6quZe5B4eg0S8Sa8rSrEoFapZp
+Q2gq2jY1gdrm9BoelAUEeDLcMNTFbQ1RcfA6gSZfyWGEn5R/UW/9b/VGlDyfVER
JNRboHtHpNjS+htZoEsDcI8WcqIIypAxzeP4fmPKG38uEGNjJz1vnDQQaSLBJPC4
1pvovOj7nI1oAS4rWSAkwEJiHMQun06cSRhKCGonRHRgEquR+n/xgs1STtj/1EnG
Ew3wq7v6tg4Zu8RTI9gi1EedCYJt6bXXm5SVlapuEGK39rVsqN4iPdducKNE59iV
nhZBXYuKyGw8j9e0hkycvP8DmW9qEnrwcJ5zXV1858H3GvoKzYts1tt6TOEDIr8Y
rsqgL8l5+59UjvyrxL5BrLhF8ZnDT4AW8kfHm33bcH7j24NR3LsBhMMFFe1otP0a
H0HtOxVFh4X2WD0WfQ5gLn+AlABv1atebWPRptV2uRuaUao63NR22KZmXZ35rMBA
YPZ7rNKABAuiVSKHMp3LrD3ZZDmIir7tw5R6MaaaqC3z3i4zV/FwAIH9I7t7ZLbt
OAdePVciMB6KZMtUHuMBmkVFPcHdmCAxL0Hb+QNDF/3UUvDUpWXVWBciZ2X8k2s4
WehBQNMmC+xqjxvXlmgJe4dq8er82yztw2J1nxEHIpe1uhg3kcf0fhlx0gOXkYSd
bs2dJax6KMG4NJKJ2LL/gpOAdYqrysBOv4T8vG8zhnW4d3MHw3kBbht3P0sQwRIV
FJpH/SlG0vsACHMRqVl41IKXFljVhz7KBBLXYmchjMVdmpInr5DiHA+fr4GcMhSx
u/vw4TTMQCXc3eSQpHUpXW+IRsxuZZRGnE3EoA5Fbdh9YWDc9KoQdHAFm9B6WP1f
cnNNHhlHG++4EvmN/TE6l1ytyr7c/NLa+f6vtlvQVua4ZEwwHq3Smzt7+ScIh9eq
VZiQwsarKyFFmbnSNBdR+QT763kmjg18b1eb8Uer/v+pikD9DIR3dQlbDN5iAkaq
r6IZKlmMAQ1BZ1sLxZrfyq9pI8gCA642sqUC52cLJgN/RQKj7eVqR+o0HD6Qfiqg
RmWCw3x7XHtTyHUvawuAi+qd5olUvKSi953/Laz1FitYXSQ8SzO6gKgT7aDBJSxX
K7unFGzydMLp2Nc/9tTQi9V95ZIh08WwvzVUBYV3ZZ5jqZAhA2giagpqvBZqb3vi
KOStC58uyA2MWXcZd8Md2ImzRaAt4qAsPP3a7TDMUjromkXoTD2nnC5iYKOGey/P
YgXeHK0GiVpiClSRNJuTaTtEju1C2usO6io/UaL7jbbLlUHYLSuM+HH62O08ev/u
9LiduQ2je2eCJTPS51fz5Bik4KUSabtyuUfNm8ZYt0Yin++EhWwq9N+m9DXaMDRG
VGucmdc8JCSxRZBjUTVk+QX8WEOhYlweHORAm9zaWX4HQX5pRrVOPmdIpC7v/uTP
WJrBE1qIHK4t46dT9/jruYse7U2B5vj212z/yDrHX/nT0xaG2gOUpRinU1EYFd9P
vstfJVkmURdZyTbqhnMRLRtkMoDaEyaNSEcNwuhW9MV5haz5LEIZ+BeHHkgwlSkt
ow3I2hRjmFSDZrA/I10OEmsnJ/0Iibm0Kgmvp2zhrsEiOrg5J/fgRqQqYh70IZOO
NzfBWsxBl6M9Flcvsg/+t7Ir1ro5lp+lDZuzQXzh8Ht8ERWFd3eMzRrvTAzmggqD
We7XDDuqBcNvrqrIx33LjrN7puRxQFuFY/2phBxD4CevkyWEMS/4cyE9u6mEEVPo
v8ZNMB+fJvPjb7HuK6yoRJXG3LrwkibpTPmFQaOsRf/ektVPQNIPg4U7OCxeyWkF
89KkHBAG25lc1jgeir1/H/0k+nUvhoHZ/+oNcAisIBCWTexzE2ftNkWT8Ma48yif
Nmp/LkXisSXjOeU/aG98kUA1xmRYj2i23LFI6+MauXtFqiHAuAA3VAFcVZX4fFL9
cNKNl4bcLJNegWIPZl1BdZOmx9bhi/C5fir8RxtlAWvroyImqyZwLnA4+/BI99l3
B0u9OBSasdpir/EPhTLu6/THWSO8HByaMuz0uxrvrTeg52rrRHkGve0eohMwUb7r
tv5b7kFjfm4/wlSaxjVs5mEt9sTtOMai8yldGO9sh/9Rd4tYgxyL7N6VdqCsmMrx
4IQoVXa5HWhBELkeXI/O8EFco9TiUvSNcZ8mc96jnt6ijHyRW7Df5tLF+eV0eqmM
Tr5Lw69oRXwROio6i0bcXFlgEHxKmqjES64WQRISwKHcf2PE0OlZJGFln1NgeCZd
XMn85lV4r17XNjCo31YHpfEdEpYbrd1cZAZBhXw47NMYlR5LjC79QK+LzQTk17w0
WBeBFzCqDxmZmY/Qdp5chTDXcgDwJIxt91tFDIk7OWJ7447/SpRrqT5nsMfHNtVm
oDkylKslVRZrq0Ap2ie41OgSBsZ2ERiNypt8a7WMxCWmr9XCFxtYuSx9WmymY6lh
Ok6TYtSfHg+yYS/I2Mo7FB+KovxWo5+B3MFOUN2KcWrZpJyXxWv0KMNsVX4G239N
ABZ98thu8siEE0C3PZDB7nx4kRluut7nlhSisSO+j83XXRnfRVA6vdw7uCWWTXgg
nPJNCsQRPtYKslED1oU++eie2CtNvDG3xTRtufjhrpplSEsUBB/Zv6cTHHAPnzzu
cwwoRjKu+e0TQkuqMiSVFQU1M0qS1pKftL+wvM9KKyafPz3zoXSTA9FwDvQdBCL8
7Tp5Mro/9PFUo3g57F8RSxLDpg6BYrmGH180fhV90fc2Xr/mlhqHngN7ETnpKh9Z
MlmU4tI/M+NO4xGDAXjmyZgGoTWBoWjODSLkh0Q1Dnz8BWlRxQBoztzJxY8SjoxQ
gIX5m/ackNOgbwAqF1cADzRIsbURTHvxcldWoPah4ZGdLr6rIcC9ZnbTYdUaCQqX
e1CSmDXpMRgLztGQvezShvUccALKV0cDsbDDRFUSOL4+rED0OUzPI7IX2oO+Q16X
2WgIoen4kEqpZwZL29SARh379ntES8h4slHTMq2IakGuyoRohr9KTtaGXKTmyUjz
5HaFfEqbBLtAXL45hjHNZW4k2Kekw7Mnb3ARmtVsvdkgPNqA+cqEbZOVdyXeifdL
qrYe4NOS0S5iRv3gkm1l3buu8C/X69iN/0F9Zm2rUq46zQS/uPAHi66WQEMDia0S
27NGeCi+lbOO2HpjKi/bP3L01LEpICDMQCMDcyvTy5+J2KSwIh2W2P8k3pNb3UjM
Whv5BanLq5DUudXHbpUnp9a9UITY7aUk5DgXO7ybbu18Bm8h5Jg+7RWhGkvQLbT+
6K00cQBfQP11Dw24O65joCeA8uIEwiHbh/QTzvf7DmF3b+NErjC84nye8Cv9eFbj
qKP4XxlwiWddinhddwSHSbKW5QAfcyuc4O3UPNA5kNuNQDtc6SFhGnf2CIfjlGJ3
TcNNHUDI02EDNhFKjCwuIpzTnn2CJoikuwUiUlPCFZA5UFi24Iza2LnIfMg6GNsF
7Kiva6wTQv+7breVbCd36UZ8SFeLLotisE2hV573VOdBdfm0yd18e+WlNzbKj7Tj
DEu2P94ouK+amoC4WwfZ53F1HzaXnMyFKN7D83+o5Y/kJ2KMRf3EWJ+ucxVbK1RD
amZYilQvUdcn77Cn0h1aII1gEuOhkEUx76qNU7UjG8XHCNpPOZsTBkMJhXXe/hP5
du4JukEb6GLpKTOSuhG/Ss9KzTJvEW5MO7bYGxgmI08NDKrRd0j0LBM7S+LBMnBM
+WR228FVgnPRzrA1kbcYQkFRRDPUUPJ3MfJtj0+eHxwc62uHXWqpd1MLt9rTFTOD
Ucv13POmIMdNStJm3D8DFgweIa6hl3abUjga2DtrUyuyPML74XDS1QXniwg7t0Wn
Y6uCzNzAhcEr6M08ojqnejGYIO11MFvGmWUptqZV36p9qQ3wFKTG08H5EaKx11m9
06bMkaaDsjSWNN5Gc7YqSC5XsNupzXs9oQJRaP3cKvzE4QHiEYPDse7g/NBE3fQc
qgm/dJu1llP/h7e6foEBO56GxaUu7BCeI0e0XHPSjyhqXdmhD+fu2Qgs1/IM32gj
cEO76XBzhJPeLmiyOo0ja7FBt4EgoM0aKu3W7ss8o0aK7NpiHAFfpIeyBfDqPbsm
XrQrQUh79VzGBseNZojMuo+V1yaCrubujXCJJ6tAsMiEdspyn6mxuDTdTQT55aN7
5jA1xYVwNITRpFS4/23jyUHnuqT9/KRaaWL+cIhRcRlyQxSheQ54Mmureyv+iyOT
MyuZBd2QawJJmDNBfgwzw4VzaIpWMYh5d/L/pQrw4Iy8cf5y5OZuK+CezNFWbYkL
hpA3zv+TbNEg/0i+03SOwhqiFcdmvwutX2uso07BUKr4VogOg1HTsd4Af0a1d9Qp
CCd/sUZNiv3ycSBCPT5aZ2g+Z4Qwk5uYoPWMShVHoipAAl+mBU5uw9vr824LpnF4
NJmGEVgwYmuLgmD/tUuiyVnJn1/tC9tPq5x/HWT3t2shWyYd6CeRYGh7UIKfUOaa
eIkTD0siXs9RvrqnJXLbfo3TM/igw5hnEFfdN2m0BZ1FNovkuk8RoKyqsJiguNo9
mhiaIopnpRQ7l9Ac6TmnKfRUmHn163nePrIwUJ0o5lyUaEZ8yY/LaoO6EHJML1zD
5oI1jskH7PxeM85XVQD0GlMgcavk0Lbyu8QDzlPhFsBY/EvgTVLIM1F+fWMWv5lp
F9KrGIXIobTxcclz0C4uBKu6VFYzxZbJzDheiWqcVzEGbgNnmEnLWfN79lR4dAFD
Va35ZaCzYSD+X4KD6mJFtYg1ylrJTCzrKomSn4pXv/8te5lDexeV9/uZSPBjGKNh
0G7feM4BghOUXrgTBcTfv31Rn7LRWq9qE/zVLQEK1h+c90/IF6F5BBV7H7PcZxuQ
YTvqzpJcOaervBktxJwNBfKlbBBwYfymqTzKHGBMZQqbjr3cesTpYrVWt8FEygrZ
IU+sM7oGYfck41urAxIbcNLSMxwTGm1EwbVCb5USurQmP6qGInkpBe47vkHHFH9O
jCb90A4wPNFiBENGAA28ajycATR3N6UVRttSZBFckEYhbxzZBo+ONaazZOtnQRu3
PtRQz3nvSze/dw2bdaXinu/BfPFWja0oaTXW11K8J17Zk3vn+rwRW70ObxBxdfTZ
jxYFl+Zr5lAWKdFvv1F0EwVWN0VIhbUgN0Aln4GI5Kh+Y4AbeYXmTBr2G/oXsDMD
5pN3S4CBM+YUuf2DU6NGPN4+yhjZCEEBIHVErzUQhE7HLMWLzq12aHiu4495JR9R
Smv4kyRiMGKk96CtPXeSrzpZ1dYswx/agHzy45XdKykqp1Pnbt+F48ZNQoeZEifC
T6MfUGxl61sS3oeD6Z7v+Wj8T6NrkQSwbwbEuN1OtELQKiWxD3xYnE35stPfS3ET
/gQ9dMY0EfY6qBAC1NnEuTQMy/XAaoxS9vpkNv35u3DuW1g5NI2DPrQmQ3nNTwF1
q1iio16hikIshC2O05tDjSBRT6hLsKQelFi/IXE/WAv08HYq8uQ6p0RQpfkG1ht6
xevS5zpxJ2oleVVPMmm4pybMSWI9h75pB2BG/TlY+j89MXVz7py58Brh3+Z5fzmB
FNeTuNYL4d7d2VDpVwicg4/dKRVk/dldNDa3Kv+czULH5rT6NRSJ8WIR7fuSBtns
9IDNgtLkfLcgf4SNJ9DN+PHe8KkbS6ipo4p0SFRyeXf1H00zyoISIPT3vpMe+jjg
Eq4a7vzwYP/umVJCTYvUvAfl993llMefxpkF9tyKmnlYGdr+QjoADpKhdsYUDreE
9guYcMPr0f9OpwJaJiYlW68gnOYbuD9Oeyjakkk1S7gRMsjacVr1DIRgaMxedDVo
1kcTzLx1u2Bw+MHDeCD+klD1oeJ0NEc4zrfyaodRVCNWWNZ68+I+3fWKRk0nqncH
uoPnkX2mPxJ2Pi6LMBYKDKCh2D9zDlJsNWVi0VCby6ZYNm4ktpFOam9UhW7exGmR
ICwJ/oxkEps7Hq10RHs2FxY7GEz0Odm8ojgcok31AvLIyzva5w/057rYDXsKJHcp
NRjjzVWyouqhtR85bSpOavISp7hbHSeOWYHJ5DmnW9wUQLQNjmqg6u73WR76T0eb
DdqOjlhcPOrl2vUV7GYawLHMd3vcx8VXBBRJPISmLgJkzj76t380/2d6KgjgYDve
AAhwhtmyHnQmVHfE0tBLfSoJEVaq2K4h2EBOvh1Ok5B3dj1PWSk/tmK0HMBTrUdr
OUgHTMOq66EsMCOmUsAfjyyqGXpzXFSP31mRvCTYDjrzY6UUpG43ldS9F83MULam
tQm9KWPBGvfaUeggX1+AUDXKzc1U7aXqFYawuOUma+ZbpT8e2miftI65WBucDpyn
Ec2vE8cyLZHkprNm+wJ/G0g8iwuQtYGC04Szp8MTm1/AEsIxLe2c+uTNHVB7MZ2E
1m6QVgbURm2lqC2MDWGOYuLUfGAs5/GgRUU3rBkaGPO5WHAQM2D2Gp43g4zqHtvM
TltYM4+Vx9I9qRDfqxmvGPBufMK8zo3eLTMqYzDPwoUnSsKda45pypsmLEym/16r
tF1jIrnulfk+tjV+LInE4aAYVptj4j7yhZVhNgAvmDuVzpP8AgFUtaWkWpTxOnm+
AZub4CPPQEB1ATMWpYuxAAhTkoOCLYTQkpffS5x91Zfl9+gaGvRyyPMKwzbWRW4a
xQNFYbBgzZHhvDyziOpMob+rSveoDO6fu5L6lOfNNxKUshPhj3bpi3FCAaa1gIP+
R6/VMG6D570gI1p3g0ITj2NPkVj4OZjpcI6I/bWtrfJBXoPPNxDx/nZ3Jw8owonB
MpiD4LsPlmlXR6k9igiWFvHyQuI8PR0k4129ZoZK3p27PWIeDX+R7PHpIRGXlAxM
afcmpuQnHhRaIUHmlz7UWD+iXoDgF4y8hS8qTgiUMpKx1HGpDxxwkORLGptZawgD
LwJtJdk9S3RNmw4nmP5cVr4xjCLowDbbdQ9+cRCTdDk5cPOf/anClFBJ+lVlv2pF
COtUuzfXVnAFNM6EjWL4uWZRALdCgc23SK3WfAS0Nh92s1/x0NKlP60oMx/oc9vC
BpV2r9/8xZsyBnSZzslckroTbSNV3WxV8lBwcPo5RaQ1RnPTeokCsKEZIJhIM1II
Jzq7OpAkSELEVSe8xGvQkL2+3DPrVAI4zQqDl2KAd+NyxGBcMtqvzgyv1F+4CM4Y
Zno2tTnhkTEQNLpm6D7TIsLPJ5wbgtQPBS0Lnwzte1vA5cBjpCmrxSes+Jiw1IIn
nEmUtzav+LKyiMoAfFqWZFO8Nn+p/O+Mw+jN9YnHtyJ+P1qn6bRKFnAkunj9lLaz
Rt+KmroaA4q1zm8/xUUXF3DyT+gTeL7g1iRnnhAYEtZ3YxBoeaz0Wefj2N9LI2fH
yjVz1GkOUoKQR5qV1EKFyUT8gTkqICRZkMBjvAfvjE4o43c0jXQSnX3TC8GHZ66u
g2y3hrcnR1g6MLN1UiwRvQLEJVup0iYfnIO7/wfm0nSNifNtpZpSPCZAtmVOokOS
EAO/slA/EMI72WLj3gOgIaU8mLjznJsQBI6/IRr/UxGqHoU3ljuCNvbmv61vKUsp
MnZ2yZGGGWzCCg9M1yv/tLFjzkMmg2q9UJKt6fnSfDJXmijQlFmmx4P1wYN/A4G0
AnM5tJlDHayrC7kk795I3PvCw+I8nQt58Iv822MbylNXLcBW0YkQ3JVHulbNrxO3
bOTwYP4RkiuWf2BEBP5SKcsfX0lyNK5man0g6WEMh4F6vFXfls8g9t4lazuiXQn+
OPLie/3UZKwENXfY75bx+VZvg+skLitLpJtnlmSQs2z9KmNBT+VU0u4ULrTi3v+I
UDeHBxdp3FDR7Bb2CrAC1HzZMATBJ9SRPKTWtt/ZZqTgBu+PXMnzJC8gm0X9hpRr
Un+xvDlZsgq/YxilOO6suFOf7tUOyCkznN4vWJAqOGz3QAgAQltW1dCqe0ABhvhW
eS/XOYXHczOdaEOcmLmt5N4QKQjL42Y8sUKobUKLQW4eaYdoelzKYCNpCDtMx6Ca
TQnvQh8MwDFHQPAeE/sUq7puWbzoVKvHQZFy4C8MMl+CHFTWHGmu7D5pp8YAyouP
Gj0dx8Ew/hmvJ8kj8hLERaD4nVTQCO1bbj8/yHsAXPby1ao9LyGLwInIK0ZeO1dK
XWe0wRXF/H74SbiwoamqBtpvHIBTjqjRsUbm3PeNcTY86XzUCoK13otsvL7RieAK
SLJqPR5YnxOkERVvxYvZ6/NMmuVgb8AmLv/jfmdPh/jbZtp3FjVOzw7Sa0qwqFBh
LpQPZLXm2rkTvs72tRw+TEz3e6dOZ4agDk0td3zkUYi2ujl0ChtRKMdJCgzXCxYK
kdqNTS9PvX8vwAztPdsgUHZJs5YSqKnQquU6JNzSQ6B0l2wRrByStP3hki95A28u
cL6ZcV1/G1ZqPnxQcW96kF5y9z23DhcIq+1bcwrz7VIVBvwvEsLzGCmsyKkmn0bP
XAxdT+Ur3DeNLJz1CkGNbEcd18FP6l95VA5kQI1pc5zq7zQEerQLiZgfDny04csV
IAsTqHa4Y9PuYQMERAcxRZLo+v2x53FRUsDPLy6gAoaP85L575UFNow/c5NrGcGr
DEvWaRBC76mJt94UHRLmcCUzvETXCf9fEypYm8nt2sk9TkG7ogjrWA0ThzkWqPDh
W8VPeAlcHKHuZALJIrL0y1+24VJMkmo4VS8HrBhn1n9orZf7kiyJ3M8uC6nItqzJ
JyjCVpm1Yp3KZpuWjB7RvEDm8tqZqy1NcIZFIvWZyvIlY3WF6iP6vIpL4FBTmbik
H9Sspa7XkSSmcS7BDT0V5HZ4r/S/YmKlbG1SF4n/qrELSMVUGnf/hk7j1iNizsJv
V38JSVHe8uGjhZAYQYKd7Tr52CILFlybpFu4m0gP7siIWpzwEJZYClZShO6sSnJz
mmLbNSb/sUjmkhTcKod90sujxlzxvOSzF+mYLxP0CfGtcAMyS8eU9OLM+AXZbkEq
Hx8frrSP5qUSuC1NJiAqS0ejzmFMkupiJI8CapW6hKk3UjvLDwNCFFpBwpJME3Fw
ixJemiVIpUve6RuVaUh5+Dnu+SFUFjuVF55ThieQt/mLlzGgFGv9v7/WYwO00Mpj
BtR1eCS1ps30s0juCNgAOqAm0k+kgppi8GWstJI085mtDeJ1XJcBQgRw+3xCepVH
evdptb+PWpvVbIvPMZghrmuDzMuYq91d8U0y1u2oqsizuT33Zp2v/Y87uvVoYkUj
mql+NyVwBOqDT94CQsbS0IspfHaXKfRUw3Uz7eT4PBAUsl3e30nGCcPCmSUPLKUl
qhqEOmHJE4RWB1FWyhyk1qLQ2TXzfQ2c5Wqsgyf9PqJaWKSEAxOMndCJ/QhaWM0Z
By++lleWFt4jGRsS/HO7bCLa4OoxJAEIC/gDqm64vPWEcEv1srRsgcGZmUnQKCvV
L68vjPf54zMIXua25XoHho++7IDH26lzgT0pxIZ/QxYNh6p0XNrRCw2xRE/7VfQz
KOPvkzmnC62xhUrJ20KIZgIQ5ve6V7Bld2AknKzC4YumGD/WW1ZoiyXpjUokLv1s
1fifjCRSal8KlHr9wq7EnZmMjZyvlMI+C90yDY2kFqRAPBwtAvhh94qREObEOyNC
LM53LSS8CFjBBGDfEF0sWc/1vqBW0oN1dJ5iiul0X9VU37wmINE1zDWgFnpMFtEI
E0IdERCPDbMFDgEg5c8bzhXuHvVO55+RpZgzKowdyQ1XFpOsLUBfACF3okBOTZ+g
w/gXOflTr27S7+OGFoAcwcCyrmaCkdLqk0d6mK6avsnOAUe2Lob5LOsV59vh67Gm
q88adeSH0Qd5m97Ul3LzhQ2BRfkR0DXtFPR7BnmMLEDT2Nn1u1DyfsqfQs6nxjbn
DsZHV4PoTzAazS1fQ0gdRtI6cydNeNZAQPAzJaBKujComPTN/hKsMgXtxwcV8XI3
k5IJai9fm4OWDsv9/BSyyIiDF03mjs5o1y6/ZNvPyUkps8jCuBv7gVwvt1Han88P
tf0u4DEEH8XlGRrtb/74EPlPlpeuJOpPOreUKsjGIOQQSB5n+bnHPuWlV9Ic4CrY
FeLMpK5gmneYmZU+QoEKbKHbw2VKTK9yrOXqUOWTHUJHtpuuU/u65EWJEn6HQkVE
L/syxsPpsbOUCMm7dsjk09A6Bjb3qkjC1a9LMUdwSKDnDnnmLSFUnsvBscNoYlkf
a91Fb+sGyWDIZyxjgFsZisF36/uSl09ZwlJ292G2EBjFkgdLT2kGW3KaEZS9kB4N
PmmvF9POvNP6ij9dYKOwVOEXoEeiFfbfEX+OyIxhEv6z+kpXXGhkO9yZJTeV0iq0
3CJMTEpRyNO73Gt+M8Dx4Z9/AhiqmKjdG24FAu+Aah3CARi89IsdviAxcDLKvba9
xLo5id/YAckR2IhZFSlZiayy9TvFbAAj8PqUkbwjNfL+VytfiNqJblhBgH1dVPV9
UntM3iwdJaMXDupyt78FE9iMN6bl8v2LrIVd04qWtMvmOthMZhuAl2j2Dfwfw7dO
oweFB8KAMpfew9lHChp2M3HrKeSq28/o4d2OkJQwuaOGF0diCK2aUdLbkS0Lxh0b
1zMMXvcR5zDM31bCjSd0YYDNdUpMj8ADip1UtrCu5kA+Cr9NyI3StAnEXWuC+rAI
fztbIV9GEPWu1nFPQn4iN7WoCMb68zEhylgBPo5jYddZtG5HKLL3VexjbJFKeWbM
j23oSgm8qNUjfGcoLSkxG35XOxkOsY5SPuq0JSK6NSAzi0y9mUWY7EAkeK/o7nSG
KYsprVwuRbtZwwcIPBB/oPlLWFZvQpLpzraQdwoxDCJEbicLzSnSOu/fi2hCsvbF
XdLrxCb2XnT7EsUgZQLOiPe6g2cxKzVTheqzeUi004J5YqBoIe7pFyMyVeP9u79C
uBCkccb73LGU/f2yZy22O7xsfaksXUzgpuia54CWqY3CjPqw3HtFyrznUM7S5Oq9
WGEql3IHE/dMBcnXtT/WAnNhsqc20OXipUZVAgTxCQ2lmhfzqLvo6NnOmutUvkNK
9ONUIqFbGa/qZnhpZo5SgQ0/e41lKwKPOmwEZWM0gc2c6PQmNRf3kNXME645QMyh
N703FbIUlXWvKgwihju2rFnx6+QGhjj0z8VqS/cV7spsH4uai0hdjs77qpDxEAJ8
qrbx7Ak/pQvVwIGz4yFR2gIvw482kwinSN87Y6LyRNmfRDb3lqmAXH2No0UXWUl6
td39EQi6MEtLomPsqLaj2Czt6b72YHW7+KI8cvNqMDGTEqKAH64IR4FnzQ8CJXaz
aRUL88kIzq2zFy+lET/w6Gion1RfvDqOX3rjXtyA/CJP03ia7XVTc0y1+BoaxQQp
9EqsPRTNlDAoIyKIeuksQWkDdm9SB9MRLBteRkSf9I22axRVas9+XfF15+3dAymK
8W7xNTR/lUcO2nvJn+MX4QMHom7hqVZMkdA5v2va+BG4Ku/Rj7HvjBuc47hkuwcY
y66nr78beEbU+sgMgwU5oj31i3AsO3wqEhOpGFn+V8GqXM9DoB9u+jy3jNkVoGBQ
n6K0MLrkr36tziE4MWy7rizRUSTq7GtZzdy4igxwq7qsPbzHR0ri9RVYwKXa955A
5iQO396sJsg3/WfO/JoaI8/XSUamhjHEgK/4kH3ChWaqaILiy1R+hMUZxYHlTYZc
qm5dtwTfbhF2vvSX0+6yVFPTJ4jRKpY7qE2TBJYB/eAn3TMgjweqMaOd0VQjEJhM
zZ3M1Zg67J/igsTl/qw9WrDM30lNkbepu5MyGxJOoizPFYfjQiLD+WIQHpiKC9rf
Yv6QatTt01kmSFJPWRP0xCQqfjI5vbVJcxSppOKz8I33OfklcIFwT3Z4AXlgfcCR
nc+87Z3uAQctWBSJk7YMyne2Tf+T8/lYGaP3jrbrH9KaBvNxuVXKm3J4HiAcRVL8
gX2IMHrbXR/FJll9A2YLzjSd6CGvc9Ui9R8geCv04KxMgSJ1JcVKC4FUl0Rsx2SA
vuGs4Js3S52e08UULwSuMrPFmleyYGOOeIkTv9cRS69K1oKQ6qoh+PwlQBfCHUtI
rEqVdTWPn07rKwpuoikoZCTmi977axo1301AH58KuD4jo3KHgT1ul+rMDtYxbVk7
qrXOoW53HoeeX33MqRvow1d78qfejOXEtwloQ7CjgZw63qh5pk1DwbUZb+cqDL++
4wZghlv4EX18DQHw26QkNIwOA5VI7EkejKXdnJOdXnKGXOtY3nLeDbBkZ+nqFwut
KWyzStVn5qwTr2ji2NbFZmmdfPPAyaLoyFuRzrzzFsz6rsXYIlPpXjK+6MoyZHKy
TgT21Jyl9cr6vHAy0QizRsRhFInAYyjCZVEtbEN8GR1v/OOXqCy/lj7t3vb2gqpW
HcY/TgADU8d8B5I9B4GNaj798I4xCU2mb7Gpl3flHR6OsB7i9pVcxlsrWH3nAvW4
r4NwjBEsmKoO06SZ7RNuE+1XQNnccGYlOkrW6/CLR3LQ2sFscAy3q/lum/kznsWa
XslqQxZbemEj2jayIzeL/N0B6tGNUkz9UWxjfkxsTLchIMthQkk9bdEEw7CdtU9B
Om/iSfb4p9fSrhV9i2glMjl2hnv7rJkfXGuo9yZulxL3eZan8sv1HDR3t8xar9Yl
3tS1cJRDMm/5N1zyeulpmpR4xBkI23o4g2NHhwOdxUaDwK/ULL75AgdAhtUoJ4Q1
VlR27IiZCheFyDdTrK2CM8UMnxOafHd0uEgktU5mE6bE/4tPIpqgUzAvx2a1RerY
EhuXcfyJuBr2HRZdWzNUIUTbxhHwPN1GkRdLWOrorxQSj8GFQpy4XafnwCbEzYmX
duDnyXfX6cSMVJto58YeLdoBf9d5LRDOwmZYcnzgRB0iDnEDlgQ5IM+zzPpFE2ZK
l7WUFrY92ipoqC0DOopU3ArkW56NOxNNknn6PTLTuQdclRVulGqaJNepjRLn4hgw
6VGojLo8Wqh8jFvYsS9dsolp97lVmiVDTur6e4hBtz7BgjhYioc8+MZLmy+XuW1M
8yFZSJS580K6foIJoCX5EJyimdrJF73aSkykCEb+lEUnWXPQ7kyJdigSDzqm3i4o
wlpiXQCFVIxnW78vuzOH9mbmsYUZaGz3nmDMKceDnJWHvQT8nh8y0XC2dtUhPIfH
RjW/E5WrP0D7LPXxepQv40gp6uFIXbo/F2u6AdSao2jkXfH5NFSpNOlJJ4zQheoo
MtXsuK8aKRPMQqyZvsG4osZM89dHA+3quUvUdFXDNpm8Tw5z7Ya2i++AGgzAZFlH
HUGMlLAGTxF/CSE2DKEJ3wIx71Il4zXvLvGLniOcHfv+gZvb80sE7QJ5UsUXCHJt
WQyLONktOd4Zr5aI3k6XAhglPSXJKSHMgNMjTZogPa7nk140GN+xYKzGEoNqh+L8
u4of651rh60fcg0xNgOWf/P5AankC6fX6RPyMIUJHMPGdaSpa+SMsrMsMO1fuFOs
4iJGNYWrf5kpm8XDPMhIOuSRWiofkYPM6eAULBUgBEj0NddT3DqS99qve1Ss5Pc8
gCO7fUyajZ3iY12n674k1AavWE436SIeNXV1TwB/zkteb1udIDjLX4enK0vmsx09
javk/H7pl+KoH0ZJxQuEYuDiiBQcSmS37OTtRykdPtqvccCiRKg2q7M0NmXI7yF1
kvA7yhtaPZU73OARwAyDl/FHioqayx7KEr0tBffb3+2Az5SWXmvR1uvct7pNP7Ff
m7h402Y2iOThDCA5hi0vhK/TMoBVOnetZE+5X+edzP+FlDyQn2XTsdrMnykUh+94
lQNUijQIAndSffgdEfa4oUoyUNrLJRGgziwxH1TbvJRtNj9H56IQYDJxUMNRYOm5
2tqtbBocCbcvImOvCtHKt6RxnigQIHybzYm4rIkQCE4199YCZYsvjBklW6zEVPsy
5Hy4x+Xe6SeSbd4aNTO8ziolxfOXREZTKcilPxD7Qg2XUujPzukXjd1I+NCzvVRh
awaL3G9rl7hf/yjMOtNTYOdl7zQwUY+4Y//7vkKYebbrr5/KfgbAUAva5jxFQ5ZK
VnQkM/0rbxQls2VvN0OvoCrmMNFX3BPGENuSEysJ8Pkhpl7itXgQprViTakUHM54
1Zs4UClg9SKZyfZdF20GZv/YHn/Te9rVecGcKiuDJL3I70dLP3PeRgZ70/X/wMTw
Xdt8PNGaiM32uScPVJV9zPgZ+HnR6BPvh1EWPAtqrEuRSH1IlLqj9ac0CrF1a4jY
YDyPxjLZaT5CXWerKSouc1fv2mCGGNvPQ9RmO7WvCm5uuGmwJLc00z/WL1JUgs0w
1ZDidU80S6GECFK7a1guhibRFp+Zcvpiiyi88qG4wA681AZEwuI/QtKIvtWFtySb
Jgvl2a7Ps8RUNDhH264qNG8k2lJv+IVHC7Nsg2nZS/8omYa6k7KiksYQB7tCf5ts
AafMibCpDhd6RDeWBIySF3R74rHMxKegswDUGYNPGPntbcAXkC9McCXXs9zFP/cE
1zdoCeFhuCn5vZntg/hvdVQWux8WYeqdwfhxaRih0/g5sREKG3D2G8/dIWB/opf3
W+9yHYeWuFG+NhjoVvAVxWDH99O4n0bUps7sr+6QoOEyTRqP1czvF4UccaP2zC3b
oiv6LPpdx2G2BWnzCsdiaSUnt0uQiXBwg0a2k/DSNGURbZe1HFgnmZI/c9AXuoOy
tyzb1hn1peWsZ1daehy08wdwzVgjA1nKTJY6FrcqiFFiVrEbygX/zGh8+6rKl7cs
TnyyzMqfydgc6Pxaj63G7K4LcW9Z3nvUdwTTcnMn0Eto/qkcoeBKwgikTxF3oHSF
dLGh82FgR5XXK4bhbwzXlOVi5Qzp2Wi5LgBkbLbhnhM48NgTRv2Bu1Pa1Wrms57G
NrreNzq4eRLqsxupkais9qYT01duSyUlqRAvtaQ5Q0nS52srsM5y7HHj8/Rv/cZU
6XZ0hSvo90YaEsk+JqABADl2118HyXUQHPGvyBNkJLFFDi0IkwgnoL6I3+4W8IGL
GC48YxxS38abFS+ixmCaNDkig56U3ao2OR5kEYJNhSXRiA2R2611aZjlhlyyC5up
wSrRDRuKiGXeRN/4UnhUte19qnGRjK+0xsz5zEFVhuCXpYSk2TxbY1cAXhW3m9ZA
g3J3q7gYT558nHwg2yUsrrKNlMfVye9mBD6SVKRiQQ3zJFrEjXCsLHmc4x9lZy0h
ysuMoxhF9oNs6bMSYD9AdnCbkLewyCiA3RxKIInxbW/jMlDnuiqC5ia9hqCaUNZx
lYOcBjSrYtW/Tmo60JPy3ombLIT+/tz9dOEA0ND50x9pp2rSUNXvaIyYlHovw48T
ZR8pK942AGq4MucJ7acVZpOpUik/t+96egHvkHD+VsSLFHKgDREMo78u/PZCROJL
kBV/B/Zk1WEBjWQ663GmiVFEA9EgjWh+7FnKtemGMA+VXBHig89h80a5vlGo4+PC
08Tw+O1GiGkzYchll/Yim6bWix7tMvbR4vR3nvPz7MSi66q8477hB0GF9+uqGl5N
Ja7DPzh64bm21390Uq++6/+NtMJ6Ws1hhCE5gb27f9VsB2UhGI2UF95TRoqwNsgb
9E4ZCL/n3KubLdkIaFknygQeV7f1vk3a4T7jS451qsOPtbigLC8s/d5Y9DAPEva4
xYglozkbGBnxYpdVoBoIMboFW+uKGRHHJpbd4xjVUSh0A3QUOsc/9a/dbJMFa/Fd
450Q72zHr+ZQ6sWi+8KgmMQobhrL6G3PoAL57SfpF37OV96Mopa76hpVo0iXr1aR
Apw9fbky4Zl66cSYGHG+uzNv0ySgNF6A5Im9aHTtuX9JfcactFyHSMFsJYtcfuYS
TnsGsYvRUX0SD8/8h+EPy6fszF9LbTz0AHQD/ZN5WJ4pbkpjNHidm1LYbGFxpZqX
ALrGA9zqndhLT9P2OqtoQAnApKv1ldQm+fXi+iHkeWMoVidJXMQv/ncMneOK/jiG
rmHSCZNF+WPd5EEMnOSjgKdOY5ioU7DswVE0SDoFH8IXRa39LQXiV1eufLyjpuR/
fR8qDJKTY7CMksG47raNVwgxPZ3Hec1AKWPN/1ms6U5xHyca2y3/3KQZHBDW0QDt
Oi89448iDzC08tJ84VsJvFyWnk19px8BKcXTzsjWr4g3Y5KMJ+sHNAPYseLKIt0j
WLi+RxEY+ouA6ES2a9qm2ku8DSHETH8gI3TxyefrGjmN87pkI/Vc+4Wi6uSJeKEo
AIiH76wBP3PTw1uu4JpZA0H77kiOYj7T3oppUviigGx8azbE4Q/o9nMstBE9FCkw
1pTohm4xDunQwqwnjtA0ZXRk4mB3JSjsbB0M1UMfAyEqkZrNnbjXdCXEK0Kzbdfx
4Yf+rr8Mh2XSszsqG3xkhfW3uuepZLPVXzeUYOALLQPeCiBaRjIFHPUIZZMN63qc
XKUDiXF1W79z4gz2tH6ssbPziAyHtp4/agtUMiJUnAsf88bLgHwFQ4/GUq73/oBv
6UFBwKJ3xR8TQd20UkKp0EXjdhtW53Hkg2MOqRPTfKyEU/cjc5e2VtHUK+Zrtzv/
xirGQLUoeVvoq9oxKX5H05XtYdOQeFadt6kdffzA154ipY8fnUxOo4L3muEACCU9
KG5ou5yw7fsNjdhdFkkp9K8Ml0lGYiHqCWexM4yAUJXJRvcLsLVWLTDgj0EImmF/
Cuf6OWqZrLEeUIqKENulgIJGCOlpxKU49VuTRABx68GnBHo5VbplBYGzdqEY61Jg
M35o1QO6VFY+PkqJcMr/UyUQGgEtRhrnhn7Q4URrtfGPpOpEy6V0/WmLuVb1JcpF
PBmCIOqhqCta83P2ehMNT4ZMNn/5xnNavn/uZVs7rrcOdc5dWh6nROF0Sah0NH3x
Ll3YqSD8FSexGwDjZvwPOUVagus0g5wCoUJjvUYSgFgZYQ93SxQZ0avO53Md7B3l
GEE+HpNxVSbNdYSq9YgBEome8AFSMzQl8z6yASA8YDsuQjwY4kE365n9lE4w2Msy
B6olnkgj3NsQH62qHhzN4DDITzRqas5xistfmUg+HtR2u+E3HC8FMa7Kw6yBK2uc
NA4fyJnUr4Yxmx5VMwm2m5pI4/SSLgcOycJ95249KawyEnCJPTXfuf6+kmq+nU8U
PmGNVps+nZkR2yBKsMLUQH2SoesaYTbYCYjOrbLX6o5JG73t8/PAy/hygTL+rMH4
X6iSJ8f4upbIxQIhWJuqU1XgOZIibD8Xfq52PqHZiCdNOgphSBEnxGaoqAB+/f8/
mmFtD8Jpg7EgUmrszrS/adrgX1iLJevtspYg+Ti4khgw63SWn4LrN0PQUrOCFNEQ
P9wsm9rHK2yEalwBdWlZRFqgVvbzUVl/Kuf1cLw73yO2NOg5zNqiMM8BPK0haShZ
w7UFZMKSGjPsMkfIDGPUkzvwxR8WE3njgbs2fRX7WXS+wYMKwHV5y4vjdng2nRKb
5hE3CUEKhN+u8rUvaciX4cqZk2HcQaPaZ9uMIbUKZ5GfDUmf/u5mfZiMBQD/CzRn
RAHbveZWvu4RdalG/nbRuMXL4FY/bjcW1nIi2NlBfPpBvH8YHAi1631gaqPQUdOH
4Wu9irII3sdZOBPNcqeamcADbk7kmOabecbjr0i8wmVWdKV6DVxietl7VboZL5rx
4dsUTm573/KGRPGLlL1/a//mn04m0Djx55wYow0NuS6sVyoHNmwsZOy4XECMEUTI
dkRwZspxOpOMprns0SF28UhKP+0cq0Tqia+GDPdi0Kjmstonx1QfNv/YA3Xij6mj
F/xAHypVece70uhe/F5YM7AvZRSjBrn7dbJbQxm318YnjzKJXOaoUzNKPVGH+6MO
egD53jrcHeEvGnylD+19DXo+FIbrHkGoKWFxvatU8bYlCEC3Bxf1BPOuzXSgmZ5K
HCx0i+Y9pS3Yq/pZFeg/9BYazKbcTx2J9g+L7aGZ3ZFu/TaA7JJwwRrcE/DPUlcl
eio3P7SavJ8y0cAQZMp21HH70pYfuwEpj43dg2vHAnOjyUULrkbQBwXuoHywB3wB
ETPVuQQIcUg9g6sjvkKIb392K0JiMzZ+VzyV0FMh4Q8Y+NDGuwquCTwh+TM4I/Iv
jF4rp3bWiqGvUKsprP6zAcczDZyoSpjoV+pCR/4vEh+Cq8NEqUP7gGUhM7VG1fzw
MiQ7CO/PAJk+0affqbB2h3bWAWzgj3edunBJWd5RQiSknCuw5nUYZxfyHGDv3szp
pJv9kkqtK8x4Fwg64J1kyDcwzvvW7gYh613JPJRknlD/OgGF3W3kwt8nLFwYXdec
ARfhm3q7y293aF+4uMbQGduPFD5ITBGTQ42JYl3QA/jiXS+yQCMgOGX2A5ZN5pnZ
A6UAnmiSeWkvwz81c1TS7VUgv6BD72aLKdHr6k+uc1D41J+SLNVjoo/QfXvll5Kf
JDG1QrPmsLDB5waSgjJXiPWtQGVvYdxzkzxH4CD+rs7qopbFVS+829wO0+vWpPaH
6l7lzP+gYSBisOymIVAalu+C5Wu4oDTgU9q5pENFBNBtfdP8aBp9gHEowAYrE9Eg
em6YHbiU0bGw9RHf5tdZyzaqmdg6DWj68rTDb3mA5HNTX+uSmBHTuq5OQNRz+sPr
qZjCnvr3rkJDfK0AhATGONG/mIkANCmQgOvu6MTmb5xva0CX6OH+SMGMF1ouPgSG
bQ7m7uvdSl2JdOgtEyVaWdMwD8cwEUYEVSYcR31rqw66DU3ejk4jKlLAiwslvvny
MFljgApKC9FtcA82qCAv+vbKV5XN6iTUfvDOfIpByzJZHQQWN/Hvucy0/fJqca1F
MBWZBmLpbuww4r06AR+X+6hgksyGS5NFitA4EZZDxS+9H74vhdo5gSDAFCX+tvlh
siCIVyTJm2bHLkkE3t7o9XTMz6KWCnzxDTk9f3ehqSSSYXNq6oKn/k6FwZc2+K1A
XX2HEwcUTz2/fZOSdtW9pc6sEKDIy3gmdLoKz/pofWmJMjHwUrvHqFYT35XuKNma
trQlrd6XHzXZd1OcTjVX77bVJSmtQLwLrqciebObp5ojb/mwO5KbEy1F5BFMZRnR
ICLl6bu8+r5UDVF6ul6K/QJ3yv7zX6LdwSCLTl/SPets+/IvYQPTEgtdmzx16GPr
q4+LaP3t3dv7oip59tBBvhszXJfK1bFFrteJ9dUabOPfirf5cCYP6lnXcL3F63n5
JbnLdsSuazfLaPKv/63BiOLTbsyoiAAkOjYgXRzrg89U8ztxpjGzJrVnqWbqKp4Z
va9rgHmzRfcaxTLBKDS+6eGr3Tcn90t8lozLPr4wSP3MChKHWgTJLjazj9gFEEGM
nH/dGwxMphvBMB+R5Y9V9pwVZkT0hRieBkyo2G/VOHWmhelsAXyUJ+Vui1AD6xN2
L4Jd36HSA+e9h5tm8EGaHofqF4kCY0Xy4XUxbmgb7XXfqrdIZ1yzlWEcl4bpHVkY
GLQmg+yR0DreYAb3lmJs27K6srdSzJAoeQeLIc9nOpK/TxnTJxbtYjjNnYuz31Y7
X8Ku6xRXGMR+GAiYgJPSxYyGIKeDC8ViZruzdzfKD9hdcWPqipIWX0aM6/UI5O1k
ynY7uRAhTIvH7rwPMM0sPjkoJDmJZxMxlDPKBunivoAngVnAyNeedCoP0R2LGjBI
7vl8GjUlrI1gjoYGOKuBcOeQqWa7diXuFKgnlkqEWKRRMS8XDcMmEpmCHu/fhw3i
fL5crRgKMJxI/vXu/RuIs28OS63XPKL/0mxg5FBX9oQUKqgxripLaKshQBgoZnNH
4M0OT3pn2DkxdvpCpcABcVsizVBs97+o86uBLopwgsAqKosIhcmfajJZFm9qwGya
xaktydzV6e03d1BzQCEbZum88/vwFDcNt/4QN7AxgsOzsAOWJrKzidelfJnCTu3S
GW/zRDz8QXjRfQQSL2ILHJy7VAMZrdomU2EOstwXsSBrSR4Ddw9qeYS737sP9Jdw
1ysIV48H3YW5MB0yS35Q2prbxcXO5+Iu776WYsX7A4F+CwpVVXu5PqRC16bkfwr1
v9RzXX/ZywsEZviRYhPfdEgoZQ2UaNH+WIbAdiEh7VPJ3D589hojRM958q6z+QnR
ijTP1vWWtqQAS+ezgKte3u74jjhEKAHq5hjv68wYItkzu4z1+H1Nvvhe9lUmDIBs
kReOv+jd+L4vizE5us0NFjn5PkQogASmpURtFOwbWrrj0LlFhKboMNyKzzPai0CF
Ktc/OIkvcoLy0v9v5HCbasvcXXQWyE1cBmz+G9rb37uppgkSCmB74PZdxZx/4REw
yOBxLOvy5XGSfwzUTtR1589aO2uswkIelcdiK7C4OyemFfN3K3aZuC2WoybmAggC
wKaNeezC7HhJsSxmGYV2U1Ye4MdaJ/4bPuvbgPb8V5F6cUz/+AvlwfJAG6td2tm2
0pC3eylFSczERVI1BxUMZPUMZp61YJHWKd8+1kmGGU9b0qwBu9ChJuMZv587UdZZ
uNshbfHhKFcuOyRd80EWVjtZFyCFbUXwBGunB2QBgVeKr/rkwfYWjcuIfWEr7C4M
XwJNa8B8mzXTLeKr5szJMSll3mA3qZOCzaazyxzcpBXPbkL0v/xp3pJc7tHzJ7pX
3/uh2jp3SSum/AIqqJzTLy3SOo2fyjylSsKOe54yyhznU5YtrO/Rjp2qo+ZfGkdz
AyQbU3KREZzwfW977fKYczEbI+wwiB7E8GMleHQP32GSadEL24YJUfQs7epReV1n
tN7wiPa+u4sDelZnH0cl+9JtNnWoUg0/M4OunBNLW/ke8VDMbCCPtgepWhh3Zfai
F7jeC3PEVpS+OhmKVd0X1fzI7wAcBO6w9E1DNkwdX1XArVh3BuYSeKSC2jJkmlCr
drdm2fhRDzKhUoHionOx5ipwtKyC6L34HUSY1s1EiGMk6FRQdMzuSv8/bDWkHfGF
uot/wwioDETV2HWoWbGbZDI1QUCJjsrcYhq0tOz1jtrCjqMpbsmY/hN+tkti/U5l
bIuo6yVY/ZW6QmnYUJ8iwPzyqBkFiwIUeYMLS2Vzy9VQRf4icFLW6t0GTJMp21J9
YKQvDB4tkn4wX0AM+4ctRc2tkveuT/GzySgbCbh0URDcqdM4Cf2652PXR6nU3vKE
hNIfE/i8/aREvBMA/o8MslZqU8GmhaS59NjqpsMgI5lpE8EjdJiwI3aXUnqoKlAS
rLV6KuLzDCzpiM4PyZjzO/rq8n/goVeyT8/zc/VMvCsd77kUvtg431OC6c5EHTrB
zC6XlRD2PO/F7zJBGVw/jb0MFqNEJnBp2cV7MtzAXX4uH4j2Yo0KZplHmxxLevQK
C7G/VjHY1KwSCa6nNQSjXo6hwTiarMqb4Fr7YgOO3dDx0b8vxJfjl2Z/26EIQFM2
K9x/gB4onZC8GNo5+x1lSiZcjpUZeeczmuTtWGgZR/uaB+Ip+eALdTTgJ+pu71uQ
X7UTMEbOrICN36khi+ECIunQ+zJAzYZBTaGO9UMrspmpwFvHTkcPRhWNKD1kHMQW
CeRsef8yknXEwEfHDN0Pm5+WV8Ow/kBlfDi2bpZhloHlKJF4xwAcUvK9eHHS3ick
/IUDiCKR+xyHrsr007snFFAqgnXnjmGPEGm6aVa7QeYy72ObyRL7hr1FJgHQKb+c
9xeSwj4YabV+ZMCaBV4/xrItnl/LkiibfpKLdLDgjwHLRAubLKb/tHRZ9boLE7qR
jZ/vWOQp+4M0RXE18OhXqjCyweNACdJBvsBDfAEME6z6eJe4u73vsP9AkSpvC+v5
aErmE8OgH9X+ml4SuWAFdwGB9jEjcQxpcw4EUWPw7jnQ8RJo4yxT2dUYHyc7R6WO
JIRpfcebRYlOUQbfkLFiDlbrBV3Oau9qYTSTH20WPF3xaSlQbHlPjF7CmHv1yoGa
NLYHxVRI2/ppCZl3Zbb8qou46NQAaCQIvS9Wjo3YCMpF30h1h73uYXcrgJfx5CwX
yHVJlXBGZI+p9OXey0Vf+w7AQDUDdycRw5gRRI7eNtPaqFE5N4wBpFwDO8BnKC36
HSwXGIGazk359IJnEC5/A7Ly2xqo2mS4x63IO3yo0gY5RyojBLtT2KB3080Jz+sa
yBRRw5KFfUqmoIJnJTwPFHwbmjWiExNJtUKrLn4HHv9DMkYVxAMYXLctNUwiZqwM
4mpQqMbVfe34Ny471wRlvgUeeynMaMcQMSOrEWirV9FKCZwL08ZcYoVdF9ijPk4+
g/YXtYjG27WZqHLfC16qe7l7EWOdKPuF/ijgKdGZsUzCQIMCnkbjNKrqKe6lLzgW
CiVMJvtc32N6yse1s0pVPGwtz7pGgdH1KfP9nmE+ZXxeoHSVCjtBe8vAhOHbFkDL
K+eDuT1GyBYdYeo/wmlG9G32+qIM8jNYrR8YGlT+RCgsIcqaR1ZKd/dkdjxEzLJu
1+moDFB73BwNrjyYVkZGTvHr78CwXkhOSMthBkAn0KqG1YaLH6I+ZJ+q4vsQfBnX
Va5T/wljTqgnYG72mCSngIivY1F2Dkgx4HG1x3pVxIGc/vXUQPSd30GmpC9M4HE1
6f7T8t46wFL4i/q/M1Ffk8Pk5LPJcJaSKp3M9+U58RY48js0BBxbFns8atBkuA/x
XlOZoV14nWxsk0pa4MiZ9+CkwKEblr6ZR5j8m7M0Ak+WSljJNEJfFcCQr1HeMc0x
WKwBPaZb0J0/k0j3dN5NseohA+cdgU61XLPQ2TVoB0a8gw6Vv5OBVWZ6KYHphh/z
j/Ms/VXy5xnLtTHNUtaNfOKvazdzLZrOF6vO19gCI6gsnlIGtreDNeFKNlY3JmqO
gKFbdr9BFgL+pvkahbrD1w1eX84MarOycY8pYHI0yh3OA2l5BNzrpOqC5O6AlayU
9w/AKHrzvnfl2OsK8Di8BBS9Rc1ys+Fg04cAGI1CMgOtzbkfuB5VrAssH7Y310PB
/9qVVH9OKvWbTlWk5YiHdxWIfuFVD5ILYj/7vc6e8Ac7NdmkEMh6aEBZ1Lm824NS
hn7rk/UmR6H6hpn5wZBqnkgyDdVUo5HeDgDnR/28UOm/9b0Ccj4l2J17XCeYbnHU
VR9Ec3ZGFVAeuQHP5k1IEqAe6GecBmRIQX8tIMnDT+nzkIal5gbsSv5I2GUmuC0V
39HMMQj1VteIvxy7ngmWr875PCMAMEL+ksPCM6heBQnCG+PewgvdM9pI/yrIw8Mi
K+qezlOxEfVB97dsfDK8jptK12Da1LU1GlVV74/CPYfIK6a8/IY8g0mGm+zKa70b
hrYmkR8A69FPqsQKO7nT4cv3Igrd64cuDi6exKVx8+olnKC3rJdH0lU/sKD7KXsA
TaLs36UpRwqhFLAs9abOseewuMY7Z071zqCEIi9yoP2pVvM7b6HulnvJJ3qutgBf
jCpNoIUwJ9jp0XNydxuoEaMxfuOkiVEeaULYmW83zjPqEsS47qDdXKy/PMTbDDJT
lU+h7rKi/10u8b+TTlrZHTS3BU4kX/B98GHnxzh2wtr9WmthbodzHgO5n3ioPT81
6eE4gLCzikOAqFI9by/DwFcWbIUnnpzZwcy8bP3SKMjc4oQ1IlWnr1BHkQJP0JDd
KzCW6bCaEvZGh9mvYzZoQwNAUT+vP7UU9jiLqSpabyuvv9JXghuzRw8TyLNe5buY
tjUA+SGSPxgDIpd5wRj4V8T7FWIg57V3GSTTvD+LK6eWPCONUE24ibPdQ735y49T
Stz2qL0a+HCM3W/Bt9dTkHETcd7LgvgghTNRlvvbqXDkLyV2dxIp7iki5a8wTvBK
X63BszklyqwMlTceC6YQsm2idosrU02JAMP3EEg3jPlsH7yjrmdQi63n+8mu1ghh
4MP5y7s9wkq5bC0m5WMU+GPdMaj+Ysgd+V017BDmp9iZMXpBOdfdFBlmKc3hxjJb
xeuKmQMFnPOBxE8Bx6ea3i9IQ3jkJFGrPSFbWKKCpwNTvkH8glMz++zhOMNmoREs
+2EaHUhtnhCVvlbTOaBTe2PwVH6NWudEyoUWe9DPYo7siYEd4G9dVBvqDVIbiEt3
smdnG2IsEm4Lh+ckm8Fcp8txOg/ZgmxgxgTsYFBdjWKat9GBJ40mEmRaEaMUdHfJ
NI4L7OSngmd38+j07I8Y/e+Nw/8UIc1156g2ApCj/l9WbwUALFp9zQB3bom3o/pe
kmcgtQisydQ6tSGcAfOD4MlAGPjkBQmkoJxUxCPPCLt/KjSb6fH04tsIOPHc0/gq
PxVkzOJhFORcTSMWNmhBk9zYv9ylz+vJVxsvJhY97o0XYgkCPGrHBFvLRUJjP7Ng
3f+sED4LwRX3ssDWz37/SCtmOx84FJW5oaRmFbWhNnhuv/yAwle2RZk8bUiTm2sa
tDKsI89HnWXnDwlLx6/wLdHfquWGV6VLYFHtHZjfpnrzWh0xSOIn79U7XBcUDx/P
HgtpAYDvGtNezJglOC7+p/yf9CixJIhrLhDJ2O4UlOQsRIlkpL3d1pDrkFTMmgbJ
WlW9NCxHYTPiT00YbvcFbZpYnsfWD1SlgUHtY689dJ90otO/RlP8YPgN3A/ltMbS
f06Yp7gpkdyo/KMqU2Lb4ngh1SaxH5nbFU4/QmkA5qA4OMrEzM+okVcz1nenKh61
zvkOdeKy7a8spIm0OGfdzY6awVNH3a/bzQN6Bm5FwHINweI8Z2Zjcc09Q5sn7ImX
SFJszvKdR4vpChhtgcbzvEHrh36z2tNvlNIf4YdcDM2Yan2oz7pkPcQrOaWVffPQ
rm1OPXD6VfgKutsr9AO6OtR/pImpSm06LHSnpL1BjaqVDVIMAz3WIhDTwHJ7+clj
FJdglCSpPorJ51BNm1H3Rr3I/VRLZDkODBSg0SFwHVsTuT7Zf75mox/niAeCH7mR
GqOnBq8eReV+BwUrlJ4AlH9hHXyMzRx6vk0g4jZve/Z8b0kgG2HFwexULzzn0xnP
49Ho6N2D/bboXYyjn9WGazDGaZURlo5VYN2v5ecUERUtpgja688wA3/hCE3rE8a8
7r2sQYEKTkQftMSWPLJDljryae8OaXavp6eFNdmFSlmzboRqZu9LqKqtUcY1VG/9
zjc0tORa2xSOquli1QL5fBN26TQGK0ygHrvv6V6ELfUNaj7hQmdSNzBbXaiqNK5F
z4a2IKE+wrE0CJeuQOLSSo5Zirg25pRofFgarasDqbsSuVnKT+z69QrYelYcj74l
rh62V0AlkpagQgCVqVT4qyhp24bTn5p9BJJR3mxfv/eRVKvNckVQzYASCNYhqt5E
ueBfYbg0r4vEAp9ItpoQ6W0FbM0LZknXZsLh+vxldQBYIrTvU5QdBQ+L5m+ooe+Y
Ru+4gpr+rAi3uGLQqyycydCSB5CpIdqYtyN+daJsegRsDKK8MZFUKBjkifwwRG79
pcIpRQWs0kGa7/AnIiMxVRBxGuErRX4VGuVqfMIQAoeRTuOZPH/ZZ+23ESywveeN
oxjIuUwzD/nZ1Q2eOcQY84TS0kER4KdXwrl1hbSsK2M4tUgjI+vPjUBCNS5YuRAd
UYVtXaiAYxRkiWdKxUx2UQLaTmuTmRtIOQg+59GvfDorMaQokLM/2KDkhvsTcS38
qiq/D+/6HPvNyHNUv63Hz2KPHSG0SI9wbv3FhJSvuddLdK65T2Li1cjKIFKkyE48
PA/yuHVpZIvem/0e7KkN3sJvBqzjo6ltNY2cSKsyT565a5o7YEnKd91VZ8IZiL6I
U6UmSypejX6+w3CNIQxIpaU9cNbw0sQ7A1rYXgjzziWwTk9grKV6W5FKItolD8gd
cOECkrcGfKvGYtvzUd8qV18NMR6XiAvOrBVuIBSRsgd9MksmP9H7SkYsizMIx2iq
sNn3DUQL1Bcj9jTTC4rD9EiE7y+RqCINAjdiS6as2kgjR1PrZiTw6xmbMu8hv+ZT
cPN7g6fThll7CV4k3bc+ebyk/dbHPok7EVY7qrI6mszPUaU7XK58XqPpefQl5wxK
30vKbqhLqpmMtNOWF8e4mJYtnbEKmAswsXf64KtZwixvOcz7H2hVkGoM2gJWsc7E
9/17etZSJfLAGxxhn85ZX17MjFjvCBIkckMMp40uJO+00ftaPMifNfO43vKeh7h+
lbtUFoW+Bvcw/V8Vl2QgOltpMZtdbWVkIOz5SLjh9TsnlMygMSLyalHBqfCA3lY6
38BPcCg+enMP46Asn01SVAIa4ysjxp6ODScYevFlNt3D8ObI5t5r52zineDLd5VE
h8L+G2gUAHsdOBlZOgTlcw50cQhLuJcMuzwuGQ/3iATj55mhmjWyJpFjb3NsqXKo
3U8b6FhvAYNBepSw+OlH31pd70V8XaSv4y1c0pgT5fnx2oc5S0P+ZJ1fyl2/2FPL
okG2bDs4SbLVFRWLs6xfuQDeEp1KdQDm1HuZlG+MvKjMwAck4WSPNMjKGZoz/PK8
x69+Is2QopfbfWIwx7xScBFYahKGI5d2ZyR+s7ZIiy337jAAj4cLyMfLV1/XHD3y
DDD++yVlJIZ1zXU9N6kXYGDU5Dvt82DTkBSG/OiATWjtRZp3/AM6vKShFMUzZC15
u7xyPi1x68FLAy4QcVbeuQ96nWh9s+WXTjdX9diYmuDXWRSVZuzqPpfzF8lL19DL
2Pvl/7gAEI5vRzhHd+5CgMuxC0yC7m+fRAb1NJppmMt5mwrx8mhWxgS49hxCLd6b
aEGhUN805tOJvEklOk8Fu4H3UmyTsA0O/sw2muuh5lLR8Y+O0HnvLUWJ5Dzso0ux
JaJ9REYb2PpxuTs/wntsBrF2NTSk22gAHKOGAA2DXYn/0ydJ6PC8tG3hWgxHsAOM
PNaRhPDDUiKg/o2bwk3+mEAG3K61mRcp8vKs+XCsG9apK5eTglYFTLIdv6OLi8rR
kr3Bs9uIwzbyRBRZpAFYsq3nCcmF2CPH1wQPYBgF23VzL9uhEo6SRv/YNNZqZNlN
KAeDHmsdO7UK2wbJtukvByOHmKxurxDmbmGaCbUSANubK2OKgjDpRUjYE8jO/5CX
sVfpq/VGQWpNBXNg8oksZ29c7PMEtNCE/18IEGvNek7Clt8ZB7ehNKiUQxfbAVdZ
oqFZmFC/I7VXqFCuY+MkfYf4c6/ZuQTY4Gajj5LrhffMW0poo+d6SKvSsqcZgAxo
nN2L2S7S97r1LY7Yz/rhGZ+9V7Phrj+k/1RmF1ckuAKUwfIWO+K9VnU/SG/hu9dQ
1LpU+nd6lyg6h+fEZUIvTmSJzZ5MF1fQKKfsTIHZjiHfaxmF8v7iG0zmMifAqD1O
XDmL5vtX1fgVTI3l/WCnDAXpytCHTtKzqjpOOkJe++0t3PF7+tZ9fb1CJXzG5Cce
YHC+vBVUkf5rp4QsruxR7Tp1/8sI4DjgJ8OFrXLucQ6elrp9tLdg/C6LdCBzsyMl
P/9oKTJItDAOObiTyLc83l2WrYzHeJVbqhYGjV8pbId/uNfkBPGRs/gr5sxCA0nW
PUbLpG26qD3yECbaX0yjrLT+buQZpC8Pi79DR8ZjdJuclFTvqeO6zxzHZKPLHU/o
A3fbuG/+TKQhE1n7jMru0TiEk5mNCzeXfACYJQBKih9BkGn0yYQi0rUrx/vgMGcE
KKlu38aN7NJBPajYtsGCL3k12QNfeIdVVP+Dfg26z5Gaw/XyS8pMw3PoKNYpjP7i
yw6R6wUsbJBQlGtDm5pShHd8T4ADCm2+40Q/WjqyKi4CyZyekBpklC+4pbo0XDf2
R2nTbyBfIEBvoDFqJc4AOpUS5Ay2by196nGhVjIlxcSXTNL6TdCe96pXqfmxrZ30
u7vaU3XKuY8RIrsT3gGc6gmuMoUjimdrfAXKTD3v6v71FcbQrhQNyEjc4lAvcj7K
wnU1rgWhNbAXqdNhH/1jPZu+Mz8EvWtlgzCsOZbqjN1ho4h9hBsPBgr6lWc8+MR9
uzY6qhL0Om3mjoiQ5C5fYHurxM3kq53Tj5lpUXbzhrUC8qTh04jpMNRCyR29Gcak
Ssua/IMldAQZtOaIEgcneca3ozOBr3v+2ENeG4GAj+7tQO/z3bsGLa4cFg+tcY8i
GaAd4eRtRB60uHLov1M8zOv81WkY7hwsnKF6sHjJW6BYXwfpBYpcU5ilN+CuxCa1
S7DuoNIOhPdvsvDlSbejn5YsfOLrFtkZWiBShjdHHtB8FPy78qjSir2/LX5XIEqr
iENfomu5ZTcV83QVKEnCkRDmtU0DJQdRfR5fcHxu7A6b7BD+pcKxeSG+mGcN0nij
tGCfy4m5WH6O+31ivroHyWypMLpAX83EDgYg2fPEJzaoWEwru19i0HelhvQKb+y3
ZWkaiExkNrzYEGb5eib8cTDAETDXDZdqHcJqJ0JA/r+wmKICkz9EyXyRtkX1OOC4
jSdOl2eP+e7Ww4quROVLeIaQnHcfkHXkPDISbAQE4632pYQl0wsyyM5qMYgWJfEn
M2TRnIJOcNnbo8CFkGWHDc9RdCklo2ip4JNW/+FYI0t8ZXsYEtYO6wLiC3wzKQnm
HA/aAWQOFc7HBlb1uLtyWVrcYFIMYqQUSe0NKYjadl2cSHJRDaTQgT48g/pzwVqB
PCmjrvKDUvLf553gPjeiUHie5+PioNLm4si/B8X3ZCjYY08q2KuqydEOdTqIKgJJ
CCHRpjM2EPXIjL/TLaK4MDKe+naR0hTePBJoX3xcQ6vm51bggMnUgEcbsApJV1oo
4qChDaDxq7vFqIWtzFpnj5hoi8fNpB+EiQqkfZsrKTVgFX8GLbAOdPuWmw8dOt8O
BMjNe+7FJqmO7Mdbf4Dh1rksUV3xqEQFBkEu47dJhdXT0Rdj8I1tux7RUDbUCHd0
3IDd1TPjji2w0yQNQvjwWNL1GFpusfNip9EE7XS68GtF4RfH/ewSg+VyPsUuueAQ
4bC3tMSNihJspAOmNkG5re7Yp2hddiH/Gz30F7+Hm63kCJcGgPVVDT4g6CTrno2b
e2R9KXuJsY9VWjJ3TvFrgkhhKJX2BMY69a1F7xUhPxut60onh1dJYuQADpJ8TL5h
IWPdW+EP3+tuRaw+hyr1P/5kWkugdgPUIAaaKoBiYUYnXbc25Pp31XwFDk5wklp6
tK74cuf6PK6fkt9sl37qRZWlXiUQdOG2X9t2VSj6xqLaByfL8uzEDg1yQdWVMQP4
8idTYl7H+35FYWdTLUtxaIzY/cmfVvhYRiw3VVrdkzI6yiOkelbxlz7oQwnLiTq5
j+HSPwQy26nBlO/aEK0RvblHAqtJ/qHPGIx18RWG4lAIHcvz2vjnt1Hm7Rj/N32m
3REvyPGzgLhMeRU6LyY5PXeGns5+4bHmZrf2ETnXnNFrVuOtuCBb1l87952wfCi9
bYidXnlu+XGnr5DRNw8rPsCe6qeB1FoyR4kTWIklJuOo6RnWT3K/SxgMB1f6Bshl
hO+DaRvuVM9TKyt8COMJI2F1DRlifgyNu2ln+EWCx2IowiDNCN/sm3Ne3wYmDKg1
767xei7qp3HOJUPFCcJdX5YmGVtTFQdhnVSzTALasBz46XuB8+UcOx83idi8R+Wq
9FqCWM7KnKY+GxSVFVDssKhD1soiwMnNcudEGBjt2+bm1bkyXfegzhaeQtKUCKBK
hQYLhAtkCHzc26LWDLXeAEVc+J2aMqzpKGjTZhb2sYO9cXnRC9EzvinZm2TnBt91
AIUh7/xQ6sq7Hd7teK//oyIn/yCxo+YF19CW4TBgHrAVIBwCKtWX3tyjncDw2mml
lF4CVBxaNYzBp9xT7X3tYrWmOy521Relbvgt6WhaV4eLx3PRx0L1TQTMeJ6DBRyC
VqbzSIuEeEvmTmWoqxc1jpvknD2JGe5KqIs/uFcGABpGP4dXJyMMnFehYT9MZsFY
qrhZ3h10RiWCmqli4Eiiq2i4PcO3IaqLKKKjRBcnidKPvsHwlQ90ElICzTWYM8GB
f6VazrkPOLjcbV4Jjuqq+S/7m+2tXkXBMs97r3RNk2T0+BQmUBJJM0UyfnaYDqhS
/m+41shwkjOBCpyB5Lvkv/b+VUs2yhxvpeHLiMOqGqxGKYhABi3mldOmBzch3wF2
fT9zkU6+6qJ9/SBhKDEPsfLE0kZ+wJFHF/b/3r8SAIcUfIl+V/7zLFZ59midmADN
mYr3wTL7M4NfqXsMHIhyq+LP76aOU4iJ4D9rsm2AnfoJC+ll+5sF6tthDSl91vZC
RLK81/jtn158c72xk+YfX1r8YYyJirOuw9+te8Z7XK/OVrQ3yJbp9qt41zqyr2c5
YqtbJxPmGuLP/axkVhuiDK5AO6s15JY4mnBmi2vdDdTJnwyXeeDhpAPho4XuxnO9
mhWAQlqBY+SK3/DWfF2VSeLhHH77uoODDZ2aZZ+PArjb64hD0EWpVcj0cEHSWYdC
q1sRZG3tGkqEsJHLvWS/FeqM0oKewgyGmWViZ+W/tx4LxxZp8rhTOB5lY7xh+aI9
ZF9wU2h5O2jU5jWMcMB5d3iS+Dt+Jzr01lsGHkZeQJLmyPTAz/wLrUzZrAblbs9V
llBGtRmkJ+uS0dxrX4QvZSiWwsH/s5p0Rw1HmtZGvnhY3iGhGbfT/Z7mzlZlAR34
wIjv8EDc+r6jUxfQhm8LpRkN/sobbHpCfrGeZBXuOuFaeneTHr68uGMihIF/JTXf
dcbIszekpewSQ4Onhp32/mdUS7jwU67z/hkV9rew1cmTHDabSG86qPbD7/RoU1Uv
z8I5n8R7egabXgf/fBXOuEZOv2a15ZkDTWE5ri8U7U+ieWx5rGzb9qqUOiiFfWpn
5wycmvOGGd4if/jQ9jCy/o9wgiLs/N+eTlYjGbQ4xOyGHWhREDKT6FwKNABhzws1
STjl40Gr5qbT4fMTdgTNIKoGUeM9jhiIIO9ukJFtGlA5x/LBKeSI8KajlzkL8mSB
pAHBAf/fgE5rlWG4IHsaORn2DqCTzm+oeePkHReWqFZPVRdhOQKsXIdFIRaNvEo2
iOfQWdgwofdkpflcB0dzLcOKhhbgS/+t2jM9otyx5dh5mGc6gz9p7J8HFV0nSCJm
JThb5Z0tr1GHbVuOyS0rPXml6eTVnttYpdkALiiEFFLdY3i4gzsmoy8bvXa2rgVS
H2utS1zrmTeGopAgJzjseE9JwMMi0vFf5zYE/FBbIit+sDDxbyS3vl5IriWP6oP1
rNPBmJqDjlrvF6aXv/uDEFSad5aLW+A0g5Zw6V9zlIY0EcNpIc3QZFoBgpBqCHBC
9RFkjYFVluhlqIblPAcMfqqVVRFdyFahT/bh0CrK5QetcvA0VNLzqMaRtbaFe/Ee
QBLP/dCER2gXARKmKZsLfFLZ8KnBRuvowwasFEvJC1dtoJqf8IyXLnETEsXXKz5F
T9XJ+m4CX5q0QpWOf4DyarKhQccOCRq+m4N9kk+mdy32ULkRz38P25b/4JSmle7M
uS+Ubh1HsQT+CbIBQYUjYMtaeV63Os6OU+bFBBG65Yw137pW0H4BKJ0nCFwcvRv0
cfG6+zirCYpHcpo3q7q0dLemfBHM1pLchyhm+dZIE0P20KNnDVtsUv5djHvRXvEh
c5g16iVO2CGeRk71qmsGDxG0HPUArxRPsLpnyfI5nqPtMzPnba1LqxmjkEUV9jT/
eYJhnYBfhoR+FUBUO9od2u79pWJdaycJj5dEHRpji6PuwL1tBdCZJ0JOe2ZwpN+/
FI5oBsY88M4XBAxS/Dw8h3m5x2qAuAymDBWHuspn+eWl5lHUdKb+Y6Cd9u16Eq+M
SEWsoNJ5SdM1Zam16pVCJ0WZOWcDwLbD2D0O83KEZSlEeunsHl9SNtOnJK2trjAO
2HisHBkc1YW6tzh9kH+BuuRbm+7b+c9nhkfJV91G7M3lNnOFEQNczDQHs+F3lAlv
GJy1PQy5UEPC5dJ0rM09vvusR8FcKlZh51pOOJu5t92qbvtvP7be1tXg8fuLx7R3
xzLg2X452gmnZ4TCJepHuiCgmB+UxB3neyo/reDBoesuaXi7IjeI/ZgdqD9E7S/V
v8XTayuRT7o88WMnQ1EqY/eYxFo3V/yq/ocvy3EB+MIzVNaD0WQrto/exxePH5Gz
kestKMMu2wSr764yGDIjsAMJk+X9WRQxg4OCgh1APAFG3sTrm0LPIqhoM6dRouQf
0Ju6pH0JqMhFloz3kOdbSK5wuET2RNF+jAWij5Zeu9O+SLzKjy7vYIKEQ8BqwFkW
La8c/CE91YM0xCYgNKBWF1A+vLe32h6xkt8zCaJWo8pSaWA2MoYK9v9dav+NGFV2
BVMZJU6LNWug5wYZkwMGIyB/4r/ei5a45d+Pdn5Vu2Ff6cX52VhQfXU7oYiExzQH
ilHJNft+QtQBtfa27u9/kDazK1FRDogqh/rVbEEmGAoAh41VtDMQ6Rg9rRDqaAEP
uPMvLp7nrR5sZ+8yLP4GtwSvS42YvzBEVhFTpScdl67STB6P2IWw8XJh5pmg2A7C
14iYCBe3i+JbnqoiIyzqxB/SAjQKnHQYAi8VmZOPXa6vNb2PADANZfZZ1NUsFRwu
itVd+qfAfbIAO+aoK2+ZfR70/Yr5CLfosgITLJcf7prH8aBPofC4pGYuKwHzbVmT
K9sr2xmXDjHp85jxTj2IXEIO6cp+oh81ylt571Bm0X538iWZ+O9xtvKJh3pRYUyS
9HAy8bUD0trp4BHFUq3rxgzFdDifX+76LbUI3lbc9i3nfi4+2z5xLIBuQ/ShtdRc
6Zo7A9o5Z3J0CHqjjCfH0RQw8CZGkmWTw+tKKyiysBBzmL56ISEoR0G1hhkdxIy4
ENDiY23jQl+ygRn7FPqy6UHDCQ9x7cwgaOhEbY2FbmMuFa4gnUQJUgGwIfErDIFt
7WbxFEz8+8uQdPiMDtllZSmVhB2/xp60U0fm827I5RQWEo/kx1o+p1f1UZPRXJlX
bKlHZyXN1H/Mp6qtX8ayjPG+FHLYMbTrVQ74g2FejVVbveOMwYbRC+8F7DAMPafw
hU9RXLtFENKYEciSjDkhcI4qc+DGkV3JbK1Rl5m7m60M9yO0vvv4m1QU1yU0s4Ij
wsYUPTqPpvPXiLkQ9Xuu3yUPZid7a9q4ZPzJ2usNvQISxPTJOazM2GwV6ht8kpHv
r4qXt9zC2X/okthwBaZPw2kFt77knMNSi5z5RAdJuzAC9EfazA9TfPdah5TVzrJM
3aFJshtOy7Id6O1pdai13C9ROSG+8HlYfa8CzDPdysF/xxqX/wvj+BjbL8V/vRey
7WxiRkXv2G0adzfdXFwAEbM/VonEQQ5LJupfUkSS/qSmgLpkDdG4QH4ukdoDb8gP
l4MtcqN2tbp6Gp2+9S2WnBYrnskxRWWMcZUufQJOYT56a8QBbQ0TsHNw2BUzJodG
h1fEPRpSpRjqEVOx2TeF1xfU7bXBYYSYE9TW6c/LQiIk5QHVeLFHsKVa0MrdcaMF
eWduIJH5DBsrSMLJD0qoAf+kSFbgek5nBdXWhkt/qnBUy4oFyydDE2pSkcRcsCwe
ZAWW8+gFOD2bqgv2RcqUSALlSEfUPxRvCpDqMuaRCt4uAxZbXIcdnAHp0WCu91LA
sLNlwhzVwW4ccrdEld+NGe5MH+yLpPoV49VXtLAZwx87E6dMneMTbdrAoHAEGhiN
bMWTt4O0PKUycKOEpXkUuCXNICeyOuKq2gEBHL7RMPNkFmckisjI1YyGYeiIynWO
9nJeyasoWce7ff87NlOmTK8ZRuIvEQ3dApw+smZqVzfBxA1m2yWEaourXc1BL66L
zkTi9ZmIBwyOz1JoTOqJ7wolDWS2hWID6emq/8u8KaZj/eUv6ab0VxacXjzw22BB
6DBZhk0KuBlJwcWgJuixMErNtLFHE1kZOFuoj/uPaFfUFn3T7PHGIoJjwoAOP5PV
aZxtOwzZxfyLglXNht0Cb2yqyoHApbEaS4P3OrGcpj6EnGPik3DJEPZN7TlArCKK
k5fmSwHnK989x7C1H9x54q7U2rD4Pbxb7bg+dlFKYu7yyBJH+kUs1EWON18ZglDi
w/0ie78YZFCX50ZbbueidODQavHsUOjdtnNipoLcjxTZ0alqidWa5OSSz/wPIT3z
Oqz2RI2bxJM7XjfxAW5HwqLaeJZQZ6lwofJbBsXU68qFUTz4ZXcNukVq5ZYyEq/c
hNowW7FWNAhqWCEQQJUTUCqTWuJITame4HOGk3WvcY6BUuJ75J3fCM2NkfYB4k7m
9Rd9VpMe5ZQM09OTWhy6Pov8XBerZ7PtqLEf0588cmIO87BG6RC+1H6GOmoKLi9E
EiTevxPOqITA+YCICzCkHhiYItK1Zhz56A8zE/abm2xDXEiNOTmz7ZoxeS9IcJFG
yUmDqHO3XcF4BzIe80VKVXu7PfSILlmN7iUswb+zn9Qpb/ZvJ+8Lf+++O7FltPnu
Sq1SvegV54MwkH0YZo+UchPuMAhCm4WnVQSmSa7EAQUVjm7WoB3CGSbuilpPlo1+
UsIxYmKB0kgY6yKFU9d2rcALq7CSDNQVVh5PwXtz23B+LZp4qn/LBF39j6LMQYqA
hp6zKKvVedhapFjybj7r5xDRw+L1pAXAm62RiHZmtgJPne6YY0yuSt/dkD3zHKGX
W0zhhniTlesXwYrBhN+c5z0a9cCqCFiv6//rgUItC4b3eWTaQNzFr4CaqpSrb9ex
O1rfXGEIoTyfR4ncSIidWMwW6V4B2DkWeo7/VqH3B3pP/4L3N531FalO0EApRgNo
GuomNBv7l6iIUSybkPkKHUTPov9buxl6ttNui6aRaXAwfnfjj4+e3zn9NxyTql/+
DUQuL/qbQ8WYA8KukecKbn4UQY1n88skM9hmwetSxAh3iDCJ1ygJFWTVB13x1w+x
jDizbml9IRMy/NEj+8TIK+Mb4NzHeraixeOjzhLGIyvsAfVIwJb2PTLPX0NN3Ya0
KLveMI9Y7lHMHITGeKd3ZwiK283pZ7O2tsK4PnRzb06A8A2qN6wy/jA23pmDlxgh
SZrKEmGbHx+44yZ8951ymha2IEy7uhlckQ7WA6FfWNOKMBjkW4A5LkaEEIJplXkc
7QpIegi83WgSOAvlEFdE8eu2XAtL6T3YDoxxOQeZ/8UrIE29cDSdzDYoix8QswzA
Ag4LlyQbdFcQl08qmAqh7u69jprISe5Sd4ClpNrRp0uiDWaxLebTb1LykA6tNKrk
CkGC5BPyKhVUvlMeE8+lxKokZ8YzUVmIw0pU8VW+etat7k6zANl2eRgyw3wECJdi
+xjCFjm4s0ZHMS2amZQc29lcsGuIyQyAEtcPWaTqXpeHV51zodqbqOnT9PL8gTjH
62h9GViOUDTBNYKGUTcwguc7Ge0NmeNnhmRuFmB7U9hb+rLUcDySdxKSErJ1eJnh
Ud5lYWOaQN8V0x4S94+SrihJ6Y/vZGuvfQPQTeVdZgePceY0clIZYnxk0vjapu5w
gFIMEsksp5AX3lnjQ1Gd0CwK/lHIZnPbJwmOLXpmsEXVQYLqqLHbMx1UizzLVeiO
AgzQ/hJkMACxLZVPoUc7ucWms8UQQ3fS70FJbvpytseSB96OrseDSIGIIqvuJJVC
RJx8twINRUMCOG/G8TkxoRVKva8KertkWKEI5DVqvSPz2YyJAL4toACIClsYg7bC
NFApWV+TzTUG+r8nHT2QD+FELdD9t4oNmdF1IZFTwDF9gOKtZaK1Wz1zmddYoMRA
qQp3+CHSVzVkEBBPJ/vGLt4qfI2O2MO41BopiUTJ/N0ruOBbQOM/ScZXH4bQjtBM
iMRJlfgTvu0HdG9SC9tx4PnSXf/3krrVodVEAWTbCIkj0D44DOAZyr11b59eD1YA
1vsRph/kR7PCSQvBqU0mc0oU6+/W8xoc/VPzudTfillaklsPMnSm/CIdrBDevPsv
yUoqVoTQrry+4HajcrQYh5iQDL0tQsSH4ZGqnA7JR85/mJvfTpEOmUrqk8u/Jt68
FdvsRCDC6XyUBar5gBp6Bg5fY7IOO8VZ3Ue9ZAYpFQC4G+4DvJ2C0Hbt1/g9CrOR
e/r+PhVIksv3+abwPtwGMRIFK3ZHHf69tyb1Clo1TL+AYgo11nVr6aMD9AIJfd5C
nkGSmjIMZiyVaoh8cgyas6YOIUSgHhqBGt5uEZ5BnO2ZNcS++rjuxA1DxsPZO5gj
x554mwCakhZr+dzAPeEMt47aS3HErPdcFOglfOxmrTLmN//YBxHKPsxDfXzzYure
diEuSD/58KPMEmCrf64g/3NgeusA8qBcN4gKfbjGEv5w68++zB/sGffzCdzK3oYf
3faZt65Xy9npkfjqdusicw0D8+87tkctWX2P7eioIMg2E4LydyZj0Eu3Zd8NfvPE
grexwrjRmSQdb0vg7Go84IkbWuUKWBgoNflnv/xNBMJzr45f+YELQRDmInKqtGJR
lN+C25Z/0im+ofjBsonz4JUpjcMFSQCyqUs+A6ExvwAUMATFPX8GNH9MHNA7QeD8
fpuXJBu++Oc7sHM/jVrv+D+urc5kSfmtr0K5LD3jCQsvAJYINKOmuVtapzPOaLpT
x8MvDT/+NKNq49zVoxLnHNxrwgKTriIRQedVaS76Ib4aQyW77Xlr9uEkr29JtIYl
0YVZduamVQ9Xzgk/7WFP+mgxulcGaTk9l4db5dK/I4NYADH21ZjZiM1Fph+Lh5RR
iEpxpK4Mj6yGfNPf1mzZHN7hwN8+GaLmd+vDB17c1LSz47QdtzC5oU6Gc7L1C17y
+Icgaqznk0nb8XKi+RpMuQDOY6l7aWmhI08LbiYfhcmX1fgHoGl4QqXLOuWBrFSD
AgbU294aDJ9MM2v92HAUAevAk1zKcy4PZZaWNZZZQ7RWczN0iZgcSieO0qxGE07K
vKXnK1wnBsv62mYS/uca33891Ps7NBCr9saJFDiM7BO6kBU8PFczzQG5+39kB7Bs
tdM5GU9jxvDXrUgsmtpc7eeToGE1sOq7Qkj0yF2ZTIAxYMHcAf/vichodbrQo3Z7
tRVP/rUB7EVfnewNrcaMZ4srdv2pC1ppC2RMGJ+V9BUccHJ4/nf778C7XPsxsX1W
dc6WmhaZneAoQqaWOrwlXcIxuaK4bdBFniE/rl1E88U4dCWPNSpq9B9bbEtnqxfq
Fswf/ab8eEQaIzMBBommjYQRT4iP3h6rKfGipdSdZOa4BMaKF3mMbnlR0+kH4dL2
4k5nT9EGnHpan14O9mrp3jwG8DclHDNyQOto5eWWXqAf3MmPLPZf+qAdQZuf48JF
GgfwKFSAjPMFrVdKy5hoLw4PJrqWwLx05ZtmnAg0rMbPUuDv2Vz0fAIjzXSl73ho
oFODFcc7VTlKfKTxebjzu9aEjnd3VnB41N1hr6fu3edjFkOc3rzaYjbwvbZaah2C
PLjOpOoyWFeG1Dz3Qph27L19QjJ0SIxccZWWilA/W3JQAWVl5HpqMY779mPc37cR
rBxHXCTl3HbAhfa0ZvOBuhIm8IRx06IwPzFB3trnrW+ATIAw7lbk9W0nj1myHULz
VtIcdwjUReI/4I12KJ01lEZ/ZZMgnc1fZpRimB1/xSNKi9cxrH95fXa3jX76Ow2I
oRSTNj8aoVZLnVj1BGuKH+oI9aqB4vf6lyXkkNhvuzqFtZdeiF4dmD5SJLX4kuUp
WQXPmCr0DkCZBXHMGQHYU/uorK8NSyTKwJmwJk2Fiku4w07wbOBF9lmcOs/wsaO0
VfgFbTt17L29S1p/Nw6V3Vy4VUNYFl0dB08T9Rlncgi/iZz1epi60FqJY3pqI/rp
TAowUkwn/uC/QMuWHvLVVDauffghDSM10gPaSyGyTJE3AJKGZIq/TAxf3tHQm/sI
wGmDTWSXh4RBxRkhrpKlTMOQiUFNN34/fYfZ0uQwXKB3bLwmgsi3gAwGY3985Gfs
DyXZugD84hTwg2cIJabW5QMkZlUeuijM7lxZkIbRiRY37JNNlSAN+y/UeeATN4aP
JHzrArH7GLej+KUir9T9oqtC1rUClGl5LoYUuoQnxJFFBWkTu59o9bdwAcMfzaBS
ZMWFIDAQ1uuEgn/dskF/VRo21YL/E6bPXlW8FT7YRzS6U3L+RP5zDEQcnWIq4If+
I/Lg3ICgY2VqyX6RTZse6QGHlHYuq5YUvM65DH8V+7V/JQkfBvfiTPeV2zSVwRJ/
JdmE6KGCEPkQAewPVujBaMOnj8SOpb5ACyMLfYHVuIPvcql7W9bN3pghGFQfdvJG
qHo9cOguu3Q1Kn99quBHfiYeWQXj9Y1+AZUS15mM/Pf73nHGRF7DTO38q7CowHuH
F14uhflKTxsrRR+yACw9MYZgR6FXKkOOvEGB65wCrmxBkmZP5JFOQ5fQGHLETKEw
P7Fv5fQHvHFyXkTWq2j41w8q8soN3c7HIXNZDgZVShb7UwgxrWTiFnMAKxjw5jMW
0q2YKAsFHlVoqUs1yD4vZmrKwUlGvFxxg9Gig+vhtNnkjw0znyAi4F3DNLz+QAYl
aqOqE9D6ULY7s9gAQc8XQQ9Jxql7HY47VIisuj+7it1QUtsECK4QfxSS/aF/lN3m
BeN/kblE56zEMOlHyqzE83/LWHeH+19YHVRi2/q6YaIdfEmHoe6uwYkcTqVKw8Nb
mXxEqCVvydn9pi2ET6I+LX7pnmboiPP5p5OS/zdpMX7xSnc/kR4tgG0xf1+LppgW
XooL/PQxFOaWNQwxpsPEWZNCztkxjFERh+beQFK5jR4imUc6zV5dflztE9YksKTG
USS1JMclqsnb4mV4E3VTZtNHm7Hg8q3FjOvl15NPcO8QUu8MJwb7LP+2suMX4Pno
Eghavh/qkEIsk7d4ggS6x7QPTS1spP9R7Bb+ou+t7gJbvLRHuIBI90NZpng3gUC2
99ZWsPHQacIf7NwIPDZmGtAMLnIef6d0E2R4KCfof6PS6vf3lC6RBvixi30xRdu/
tZWaqP0QAHt+jjr5DjWYxpmK6aOiKELenJQtIe/BxB3gDuGD7kH3mWwPtBR8n/pt
g5pRrpzk3XJL5EVyQvBxB3nV6wcCycks8Of2JusPiqcy3/sVFSHWEcgW2FhPx7DM
w/vFaQPNV5ulss/njN+oUc7NiAwYAjRli+gGScNKbUfel8OPLTtDFSaXc/CE2+UQ
8pQ8uw93U4MfEopZYW7/0DsROR6wlUqAqJfJ4Fg6OljRVy6orQrQIGhYG1A8sVG0
LJo2xfPshiIezXrYrw5ohOWi0xb156e9XGfXyE4d0caa1YNwa0AAAIdtjegDaHxI
fR0vvnb1ZmI/cITOmbbVemRGMvkp7f3kGRs68G1Nf41mOjleM1MHE9EPPxERLQ7n
rZX0Ce6k15y0y3oQGx+lHtUoHwnoN1yGEUGIEPfjTthae2TIJZYxnlAgEGr3kp78
AG59l9PJQFWtZtjAtQCHadWeY08u3mI18HvWHQSzQEqNh8mFa18e3LisLXzI2nZV
lW9KJYt/YgESAE3mfLcJmtVOVCvfKEn71Ys1vgkyAcx3FpTjp2S2tFN7NBLadhIq
ZTzAHL+j2OSUeT5ApxX8KwmsoPfAKlw043VLs0H2GPjpH7YK4BDbXnfqEkjKU17w
Aq57qTIaQpVAfuVOGY79+0BKl9P5pPHHC9yFm3DmQBh+aNcTPvHgdLltlsGSdDhR
oBNYBDviPR3SRnRK0DCJKzjHrgeeWc45spXGRF+HFG4hgrfSVKIh2LCpJWHHA/uA
uGxSfT8xRbMtIp3/TKgeL9WKm/8eRxl/k2PLLgD6dNSaY5ayoQAe/WZg/KZ9TI4k
Q68LZeaO15jAVmkVsk49aEmemINUx1I259GZhBxblbG50sRjpjYM11oYy1vytaBp
cO+li4wb3kVCzcp5fh4+wpE5wBMacwRgvHgo7NpS/+GdzYGq/DDWsy1aGvtHXQ0r
3u3/FfO3rLICIBV8q+2eOutJ1mHSv4gHwX/dzZ9nBIZYf7auBFYEPDDvTfbD0pSR
XtfUWF7A6GXVGOyGGrXh+fB0A6wlOcOuhM4RDywD2/22cbFIy/QitgdOZtZBvVjY
Jn2qsy8aiWQcxVLYWe16OWqmB/PcD8Yw+e7+xYPQNcWfP3s7QuQ0FLcfuOeO3T+M
VHv0uVAyxLMmyVtFByt0pfBAbtI9S9W2I2p4M9xqYPOmlb3oTwnS4sRU8oMxO9H8
XITaykqxwVAp4VukVtOlhiOad6DVdv+cDS4GEe3D7r7tm1MFvbd7mzhtX2w2F5q4
G+YA2VCWGO+Q6DOvX+De0iMVw2BwkcZ201FnjTN7o9g50ypBV6kwTPysaKqyF7/s
qpAk90Dwj6XQaTnFSY/hJt9qwFV9gNQFMmQlVFN9pxTEZvfZMN+rIfnFc3v3eOjD
8ymCnFaB/UPFvNznYX11iEm4IHLy1P2MxKKMQymK1mLxujEEpGU7PwCgS/tlncwe
x+gvMGXSBkAG0ec6kvDrjREoOTjEBRogUOIm+d30e99EH2zFMjHzm0nViU3fisYJ
Q/+985HPDr7toOeFomVbseccv0EhmQYMce9YbLiVn/nzmY6UTN4QFNat8PFA6fgn
u4y23KkLPCtQ1c0m4esUHTrYOYYf2bSegLkyFWq95pjV4odJlUqwbbhyDcqUMQ7L
0FWUVcN7t8EtDBQB6sKIzwrwPWTTHpMxaYFSXGjCD02LWtphlz7YDCbTf/Dhy1fI
vDK7TNoLzBRjheLYqYJ08bZsIAtbe9grMTJgpyGbE4HGlRrRzboI4fg8FkddP5To
EjjXuoE0VEhYjVmUp7eBRrTcHhAwVK16bcCMKY1XY42g68+rHGuKS1BRzdPXO6eG
rOIAMTwf557fR+eO0FZkCkLxCUtJVHCGtapCxBvy8H85CJa9NDHzaIU8dckm2C04
hVqffR10O6JTjnlNIbjrTcJlxlXB+ngZmYpKBKDBZqVVJLVUOcUk4Ykj9G92XCCm
N5Tt9njJuh0B10l8rYR3R3UH4WP65PDN5ES+Y4QU4k418aMwBSTPEoOGVDnjfApe
KYkAyMPvlj61WT6TYewyNX9l+AGyPJTXWK2QdBOftRRwpQMHCq58iZKxTaJtlS49
9CL2Q7lEmxa7Vn7Qyw78VYoRtIzifzQGEKetdBcK1zCIIhzTs1Y5gjoQPCnAjN1D
Zzdlw/n83NswWxIwIU47DAm2G4AB4xE4ErfndQpQmS878+PVjfpEYBiblULDljZ0
07OXFzGSkEQd6ZXOw8R2+EW3Pt3d6iSgA6QGFMH9ZF7AyWbwuJr92fHbFEzowAKb
VJfeXrsr8mJdAUSIQr4Lj5gZS1HcEb1hTGLj9zJ7yGZtfdBKhGV0RqYCyTKTu99y
tttL9J5kpC6D1fZ8PUfV4wM0mCLKNCyGZ6Hi8gVKeqKIPZraF3/n+5A8MrYruzh+
HF45L9P+YDkCpPSNEO3NeY0Cytd09qVxgeKorY0AGVRTMjKKbAqMop/GQSBiU6NF
/JwH4EjTxOA/PEN/jSboiQFPN/FYnw4QF41UukPt6vQxS+ASl7UcWdFyVNIcrWzE
MctRy/zuLjOaL32UsN/6w1MgU5agI/bQCyidphjUnptUzI8IwDnPr9TSHUZOQ0jj
Qis+q2EFEge+U3+8v7/jlmcPDYP3lVJrWXZHP7/JH082ABAuegpuIH6c21cyIcOJ
2iW29zXYR3dF49/dK+K1NcZoEhINL8vMAuYCu1l/3PrDNJfcU4O2E3+pQrtJI2DU
OGz/9AuiqcNGfkHnkuF6zkV6Jt6ZO/TK7hf0NyI73kS5Km7pwX88Hd87zA0Su0ro
hNg69DdasLkNesHnE1Qq71VlV2LtjZ0Et+ZKyYeMJxcL4YzmcNwnOOjTD+he8Oi+
QV+o+at2cdGM/5Ywrj5frQSMK8fCae4FAHh1cGeDiw35GwmCeoF0QD/ntSouCm+6
cMFvVaRwSKj+phVz6Fc64ALi1e8Sz11YvxiNsny/L39GP6idrtMqtOQn/H3pADDD
zPc2FweBPbYW+Ok81ySCNAkKaMFJo+n39l00nC2Xv8obqzz83akS1hjb+eS6dRMr
DSnGBxfM01JyDzrOaLqtVyUzpT9GPFfbEmxCQolQDSx/FmUPuUUCiLh3tw9jTlWh
vloXNlZ3OMrAyRehsJJ5lCZ4hEi4X6jSbJ9UEfmCcjpDzaladLk3gu6Vsi2QFtFo
2J0meQv8esSO0WAi7bay/zTCeQ2MbnTA3z+rFTi+OSgfjzAPpfB9WXO22kf/k8VT
u8WFg/5NfmG5od4X210NQgwV0ZoRDnMz6ZQY/gcmkejZzY4U5vME9xPrFbeShIYR
OasBj5zl8ooxRItN//0B5zloZlsluc42COoBXPBvrP0Av8E627g1EvtDX4zpi5mP
zEVNe3Rgp4NXpCWHWpFDrfkqgDapfFA4FpjWHIpIpr7gre5Lotmrv5lyxhFMXaMp
ICesHmXO3xD02SOVbmGQAN4KtiUQswvWvY2qxsIHwl14V5qFF+APdxxhHTKukk7Z
GeW5PqIVHccA6cjjBQOEKqv6APq1wY10ZEazCNjZYk1M5A+Mp2jgJA7qpoRhEYrf
ymt2LTJ8nTcXji2wsd0VoOz4bUkbUCu01IOEFrHlw5jcXyihnbEYauZ6VfDyHTBq
jB6fj2sPRpZMKNcFZRUjziK3ce1VMAsjGS3eqXz7HZngD5o+5erwUZWfX2Vn0bkj
4e5DrDYbpHUCQfStZ7qiPQnMfkZTJJexMy2rQwRvysyqc6fmZ4sE+Wy7k7cYQiW/
+DUTetTUHJmEO/EtsrXkEsyGDRKVib0NECG2j7gEjoozt8oMORUFTi/3iEi0ph8t
/ogrBuVrUyuK3p3k3ivdJ4mZOP6sykiD1DC7Zv2ZzHwqZfGM2gEQX2sqTf52U7cX
HQ603pT/vn0u+z5+vprHyBTMX+TqnOLADVjAyu6sgZH4zUxs3cErqOBZTgTUH5dV
6/H2T0SiQOqVGYosFygrAcBN56jY6EANSLArqHjqmQBjiP9rbaJorexN7OOPAAI1
66VFiMm/7CkVw4w33iCjX5ljPMD3LCaEY7joZN926enyiH5T/PtN17bniXANi81+
0FqopVjgLbw9sXgYSMf+kIbn6Co+7nJJrJh86r00Z0rx7kK+FXXx9EbJ1gmJW803
caOQWLz8rtJK5YowhXEAxh0z9jkCx5EkX0kYEuk3qJHgeKAPqHd621p6goUp4ojP
LNEBl9jzQ5fNdilSoxuuPV7Cl7ceeQKgAXNOwlylehlyZNtUFrqNQIj33Rcf1pWH
8zzgnGSLiv0uv16hfBDmf2sTaMxQRn9eKAAPzBWUKnOBI/IyOoqcj8kIQ8WUO7i9
9+P8I2LWBkwCJzihB/L8g1XfL6jjlu/1DfeVMpS7PCn4qTgLivvBG7hw/G2NU6uf
cb24zqcbumjbMh9EmEFxo71WDDSDTfL//gd1xgostl8QyvfHky3rNi7Ccm9sV/Dz
B70G2NGFJum0WfGtBpZ8rO5YytGNjjEvkQQiVy6QvnoRUjz15SS42J/BCL7E+D9E
skbpt9WcTCi38/2M5cDqODsd3ZMQPLolzwVhHacSN12YKk49zeFBPDqARrl53dCy
/49b4xtwV+pKSLCcY+k8Gdt/rzhRv/PrFvoIy36fQ3GJjYXWJ4bg7+tNP4EgTWEa
HfOXLeZDS3fT7ZClIelasTkqw8TVQ1xNQGZSAXPqPdk+qgghbHxska8IrJk8s8PZ
+seWB07KD3Q/3pRPaPG9tjBcSefFBiF3i+1VLq44hZ3EQlh3W1th+0LNljQJfNBv
iB5vBU18zFs0gpWA9368WckUulkOXNO+rxtDpbOKExx9IhRZRzHBcZ+UBicZUpnc
GV2LoRoGGjqG7TvjVnO9USly5joTsUZuJ83Pkb6hPLqQF1toaLT6/r8MoBpEIH6s
SNcpxZUjiJIT/ZtaCvN0p9IfOnn+/OIurM7xwKsyG46HtEzIswcQdYjLNBQo1cwF
NUYyTzCOvnuE38/nrIFXLsxJW6RcxEjTnWLaz96r6HamxUvz6AA/HSfMOAp6H9y8
nvISQf9k25/UoUD1dnNY3oJukFjeF4TLenihz7huaaGufSy4PKdhAsEhv1xY4+vT
wJRHSb2CkfxZGgyuNw1yEqAqO6JXhzvMuvI8lyOQIx/mIOxkYVNTEhMAjdZYclJf
67LR6XuUCqGOqez5ujE5FUReJvCf8ngPSCypot9IFzOaVosIXqptyhoTQWBzWeh7
z48LEM/ewo/k30MASVcJRbJj9018uu7PpH8+IF/L9xIS9vPsZua800Qo85jpX845
IMz4zaYWoc12IriExf9ZzP/LuVNXU7YPzTKcVZfXfc87WLM0UGLoiQX64GZdBsQw
uk6gXIakrxyJXk5U2vrwRS7Qu+TbSHv1PRRUYOCQPmHuuckIBXS4fzjR8LUj2+Qq
uIFZx/nI7NTPh9YyN09MUx8ybnIirsVQ1O7V4Ipnk7tT2XffMduj1+GR1+toX2pE
aljwaOBQK4x7xVLkiZEvbCTQEKITilMpIToFPsE3iY0trY5kljhkLdt+NhDXVQgQ
lIXTLCvHp1zS5TDd+6qT75BNlVhBJbxRRBlFEGEv/M2ETN9AXAn06pq3CNvTlBEe
oG9qXARp3o/6om6YQFY8Vc+Unwr4gOakjwlDW6N8gpt9oFMDVwwSHr8aXlCmMfLq
t2DLNwbRGD3NKSUCKP7EiAMgyfmRl1nqHr7Tarnyv/ywdeU0KAMFH6iOim54MA0S
qBvG2SZfujTskkOXYPJ23yUtJYRBVswmqisf85k72ZrLLV6raaYy/Q8tp+YZKSk1
kqGOy86jEjzim6/IeUNXGSHRmjrkEYh5D0wu5CRuDy/lX+1b3qfzVfyBrpm+tk/1
pEZ1HSpX6/zosMwRX9gbyUQKBEp4+hfx/4Ybvst28U4aNpX8ZfKmQgEtzbTO7sko
d2O4pIZW6NbLHb0MLecgLodOPh8t6h62PZAHlp1KMK5YH0wZlenWl0l5m27py0NQ
Ka30SfKMjkmFVUks931DwZ/nBYr3UgklCiTMIrP8ip8rHiAneECObzl+sCpKGciM
e22cMOzvd1bzLxCA7rbdNK9kQWob538XjGqJtNEjGwwUap73XtbOcdEXMk5abIjQ
u4nH1VZVAJGvI1C8yGCamE/kh9wkim3JmLBnGqGPB99ywdlETrbnl13r5PJU0HVT
Lu8SRXlQNqaQ8yT+3+1NPrhZsH+6+mwWOll90h/yOCVLtQTgsLVz/yWMzYifsRx5
TuxHYHHvs1Ci4i1gBBBJ21KS+KKvbkJIZ8p/THhgfpKWcXBOILoWah5qf55vJwT/
RjXCMAIlrI/WyPOOraF6en8HcEaaRD0nN9VganH6+DzL59t6y3GhAl9Vx+GCSHwz
2M9jM0SRZr5ZeBRt9wN7h+05N3qNjnDNI3ewY6l+t10B17L1A0hpZ2sqHkYQobmq
m4qPmhb0B8u3fbvcFiBp/gbOP2C4Snm1mj1GyQWN5E/BYwJgk3shYQfwq1WWGgOO
w924EubpEcVWJpwe3AlO9Gy7D0dGvLIp9EfEkNunYiZMOXYcJBMSCE6nDZf/nyr8
yb4zN2RoTY04Hg73PPjMJJzHLUoHefEzWgvifSbuJdF7KVF5XbXNgNeW0hRfNqvZ
j+Ofrs4Pftv7VN9mWTyv/Ql9zW0+TdqR/q51105R3TFVex4Oe/lwvr7eHOOC7JEE
bSjXSV/dirR6QjWmzOxZtH3NtwQiN3LOjGmEKrRLyFQtOpTJ6jl5b5/dY9dRIcd5
9NRZVI/gdlxqiurpqYGz+lMsIAf323vTw/tLNjUQBYGxMcQqWcA1WIoziWtbcDwx
XVi6h/HFnQ/e9p9lTfs7c+To9JhksRO0DfZy7pjt0vkwKtfH3c2RbR8Ltd8cz6lT
ACe3N3Xyff84hqYyajEm4lxro6YDPHNkChzjGTDk1TDOj5uszlQGWMhd6CnV8gRm
BrsV4Q4TIapxWd2ncp3q1gu4bfRF4mvoXQTADrD5y2swkAUotYSiGiLlUzLP6mFj
ibb86KZ3p4K3ptjnwYJhT01Ua6ftHgmPEUOERXmBIZt+8qiERoIh4QsIsoMEu9Ub
d5Eb8iZ3VALe/+VQUOanA8SEx8I0tD5IBptK5oZrk4fqfuUMZRhzT6sdm3npTQop
yDrRsRkiL/PRPZ8n6NoWI2w1Igslb3ilJAtl++VUd5I72vuCKi1eL24818HEpWao
1YpgRxvFe5bZOmMyqvIq+KCjCGBudyefb0paLSYmI49gF3HUkRAneMULS4VI/vLw
kua/2Gtj/hIQDmCGpyHx6FTGVNotFQrlmAsIa88gvFFPhkHaRsusy59AWqYsuGYK
FDuWZX59uiS16sb4gY6ABeeOw39Fm0pPA7AfyngPiSi4NAmd2TxOjDINDqHtHhYW
UxqnQPxRd4gdhgeecuTOOe3kx7rQOdyZybm610bZVKHuOv937I9oppZYtXM62hlV
8+UkONb40VWN/QPonqOZyztQ36Q4tFC72pXY5X/q+IanLDAbeoT2Yj3N9yeUo9qI
SOOkk9Jz6C5y1gPWrKinLGt785ISq1AlBwt4dRHI0R5eYmHQvImPDUVjZRmXfsut
SohP60BFrnklrmHArkbR7DnwQyIo7RohPAVyq5CK0yqbOnMr8qb1hxcije8NG2X/
uI4Axa7HJfkXgIB1DbnJJ9GtCvCtAk9B1vYoSMa+LG744XAJ9+GlQ+YBVV46Vhhi
fJPCWRf3kH2mCMbHtBZ9zZ59VSrskVtRjFzbAqgM92HQlcYi0IU0yeaNTWSTuWfv
MFPRbi/DOJmDJPm8t7d1c7l/1gwx7HAlDWrwUkDPNtROxn9k0f2pvkqz9BbsWGJX
tMeBdp0iXvdX0I9id6Z71sqW1nwtDdH3pB7H77XOZTdjUr6Hpt0wh1We2NBDFpUg
gpBOIY6lU/XuBsOKrEN6R3pNu/fsjhAGKne740TUX7nAVz1u5P1oHE4mmudGoiXT
rSXCFdFxxRayUq/X8wLljYJk5jMdHBUegT1wL69P1qdnSAHyXbXu3sGB1TJ9qAFd
m2mCZyOq7lTYiIx0DE/cfiO0ZFuOuos/whxbhlbY5SZUVykqkizsre5x4xhKb1AX
aROKKB8tCyWaJbmdKzG+KqrVqq+PFbhMyleMslVCA1UA4lgXk1ThWxeybaSgPjBv
LBaBLO8HN6XaRtBTRAyZy9o9WyzzupACbGOCNvJTfDxfYUaPV6mdCg3/boOBer9G
XuaUXfqbcfTYfL538vTU1ifRvWDOl9hu3+WTmnzhrXgOeAr9capgn+z1Em3300gG
vXCFFfW/6/egU1yNt5EsYJ2cHj5qSBLTEOALrAUOWJpb5CR6zvIS9CNcnBluP8Yl
c4o93G7oG3fCyiv8YJdfBzmSUM5KRvELXPz4nz6x6GBpT3RnF0K6pkvi4D2ky3r4
Chnl3kJT/bKg2TjX2nadrJHaz75FUxX+YtQ3kpEuqDmUuJwRN3BhOEKX7DLrTz1j
JrTlK/j7CoCEL2fksyqH/8elvb5tbY8AVTPTPl488B54cPA16NBBPd2Nl5afxtAt
rBD5UOUHaTieHgwf1d9fk+gv2TSmUWd9gpKHHvPf+a745bkS25xASkQHQDrJe299
QSG0JMpnAvLi703GIf8kImr6gdpaqaLiTF9DFfwBkKVcuidccYJQOweDdEm0A5r3
aqOoZOuRWA8CjfOlbHHG41Mv1mmR6ZXRHE3FX2o81xre3q9EuuHO/zXJ5mdGHKWk
fD2bVjf02OLFi337JRJESWHj7k+S/Wuf/HKg3giNi8pWU0P4ClY/QP2BqZ9bKfKL
eZecAGHcvshdixKPSgEcJx7EBqe4Ew9sf2G2c/2wi92FxvG4jPqbGrJJk6b+fRzt
GVhV7yYyrf3evwFPiCaIkjbmIEidDALPdkQGsOkvJLQetm5v8VsNd8/k4/z98a3n
6Ct06driWJ4beW7XJpX2nuk99SvohGSEDgP6H85jcDxuk5ly9RCNOilLbzJolJvZ
4Otu8LwyipIchLSM1RiJt20+fgYaiVG45L4DQtTM7p6lhUQPiSnFlIKlQpkae7oO
WiAxNCh9HDIUmE5xm0BOq/dMuhhzhm0Y2HbUbb2adA7Gx7ApZkGCZ450ItFoIDLP
6VEsqezBdD1fb7phIz2QH8aJScjxD6mP7bNlMxiJTgFz9+9wRIZ9G3/k/hTrK23n
NQevoxcp8kyrkEd56nXYC6ZT9fUxdOFzPZ5w8dtiYEngxb6lsn77BtYWhnBsrrXP
i+gs7geYnmrO0skCfxKjlHjVrb+g7jm6GW9uexoxiNSz55KvRwGeC9ocUmMWQjJO
l2cHCaoqk0HQXMjCLPEHfjPf0Z4QOMoz0LX/11BrbGCA8+vjuhHcHTch3BhNzm6F
xR30mYex6NJoS4lMBwsvqoC2iQdcU6qHFKnJ8pRA4ejnNYMXySUbCd9c4gsep8pq
q+BiTqT9oRAX1oqHhZlSjKMUmmU8VUcgBeczLNhF1yRaGBav31eRj83NC2YuGGxb
/j3hrTwAebOabCdggb7Vkrid4i0s8mowQS08Uqu2IQLrJ9VF1bdDmD7fP3bKcBHq
gS9IHl2qEco02O15xQRygMKnIYzX3mZB8KgOPYY7NFRXvsL9wLIigI0K+BQ833h7
BnvL8WELN1nFLJnaOmGhBo073O89Amz8X7K4mJU7teOs2TGeejqolhCSAJ4JyfvL
SANuoXVTqUxTPIx0TxWU3EehFxsIMlIztm2rzG8q3v/bILP8TiRUJ9gje0pM8rkc
pmoHHDY+6lJpI+Yh2Ah/q94GeDeIw4WEWz4dVTjl4qkFT4mPAdIhwk1I92wJMUHQ
Xx4NA/uAFPNxAaSPWWtsRywjlZaf7aXd3ofgXSxGkypuMhdY3Z3++VV4W3AFAf9S
IPG9pkzfvgSgjzxXAhNxfgXWQmuZY45dstwWOWqdepVROPNb+SnIQCaczvH4xAlw
M9FBaNR5cf4jzTBTlojMMwNf7m2kngm1KjlKZfVqxtSYvC39KAft9Q40wIxdtXuK
+95+tv6mtI0D8eFHdEcRNQq9KgjGxj4HLUuDpHwCxAKMx5ugr4WAmHspQNjpN/wB
DE+OQs4T6Lbfy91YjJTM7LX/68Uqo/R/1HOkIxs2JFGnl4oVtMj+seVn+Pfz2I2x
sv9/ac6cstQDWC5d0AJUEAmrmitbzvkBtd/NY0jjjpjHLZ9p2uRuyfo+FL3E2JkT
41HL3dDpq3C/pad2ASZo5yZ44Xdig7Z+HLN0kRKLlcEWEIL/A1+O87NwHTbvYAty
mEJa/O9D04haALUp3p7o9G0zT9Um1wTEv2y/VhyyQaZsjp3TaEjrFgttPYLyANHJ
olhgcK/TdAEhk66Fwf17cZQ9MBadG9oO3C8HZzxO24yFj6zRcwX1iX296mrZO3dw
jC02JH5kV5YCrRdZkdrUmsmQXwIsmDJPBYMXj08Fe8+Z22k1Qm6cLVM8fFUUV6OU
cA7HL4/mfs2tBi7xfo9qQys1IYB/fqrdlPXlbVtI/YyNvJUwthavNz5pMgtNV4TZ
ZdN/tZsKehxuumtZj0nAfhiU2t4w+b10SNJdi/TxByR/DKXrzwcDUpaJyAwPmBSE
RsfoJHe7ZsMnjJbB0796XY8/sh4sKH8BogUNApjStkyeWOXUB74eBdVpPm9m1eaT
eyEXuT3ArmR9z8U33k2gqIHMmoZe0GHmMzm5fEO7tSvAY7Vuyk2H8Ex2IvDIZaeM
xahcFZr8x4tF9R/m29sf0EVXMQIhWIQNymNLEv65loms7deHizqoBcBS9fuauEHn
mkLApSeKZbPevtiglMv5duyZiBRVzdrGBG1ffHWNDHdKYoIHA1jcGC5gbHsVtjgd
ZAlOeKFvPGA67EhxgNCB+eUQKok/UGWGTYIkxODkva2xlwlZF807ypJepPez/yUC
Vku/qqciexB2qOX0N/G6uvdsLe8Oo3pYq15Uut6qjVg5e8Zd8+sTjgd9A+q9sbiQ
rRVi6hUZkY+IpLKq3dksmEev1DIy7wCtLEY5Pw78gEtXvgov/zKLoP2VeHcVr+tJ
ZHgxBVvvUGRS/3I/p4W9Hp4FK47FtS5fzvAK1TZ3OZD37Po28MsEnW3jbMyP24Yo
RwJ3oUJGbMssUpixC11smhnDdxrI3/M1rdMvUXI0AdoPToUWiX1Oxw8QvwvyGwvO
g4a3v8EIIb8uoXQE9bB7Kczz1VMI0Y4p68Iv+Rz1IAFFxrpQhyV/yXF5MTwl8ReQ
0CK89EfbWdZUlKkqsl/HDYtPpGqymZKjMLl7m98fH92CWK2PR3JwY5kDomfj/Ziw
TK2Zv2R3kyrzUCrrigZ0wnDOPqnvpjJ0OSNKDt5OLqOsaOQg/PyyoqZ6XuJ+/b9X
jnZ0ToOm1YaGIXurngQhPvdggXOYVbfFFm1oR8C7jU1eXGLLrtdj+4LezqYtM66h
5sXG5W37/PBn4zVWr6eweiWlpfpZ8p28KedK1eIsTLLBHz4mwJoE86IHbudhqLHN
aaXlCY52ll0NtD82xGRbzwOYGhxQLlsAOUvKRNb2dmIPp6Hai0aGV+5HGoTVuLdn
aB5vYr5FSSTtG5Annx8XZpk5vY4gDimUMzLomli5ee/ry+TntGgRIUAwGw/plqwm
+QYfThzRxXggcY+DnCUJ1wZjWTZf3itGQx4pVsCbDfdh9l8fWfFBmPGQfLSTP2w0
qxgZLBzVa2vXzXrMZgEK9BhZXGUhtR3f9BbtWzMeI7N0Q3A1qd0YzFRjRD2WhT2u
blxIVPzm7LV+GF3HgkYjEV0cUt1w9pAJSlETMwfDR/Fa0rTsDI97+VHYdTCyXmQe
FKBrptCVvdfyFJzbeGy+uIySusPUYJLXSNBLgqsE8ZzCHeIp4FHsSq7kFByvr3ic
K2uzrNN6HWeAEmxEuZY0M+0BjbUjfhjLkrZeRnmc24q8C330AzQiv5hC0dnUvpYM
Yx+MsU4Xscf1F4X/OT+ABAW549bHS/uDhr2UqIZGetfwRCM49u8NoQ8iPdQvnoLc
Cke9yKz30QnnSUGul80b+yDbxy782AslsnGeoKz5xQpEFm1aMEEKSlcJvGgAwkex
K+Ng/l09u6pFE2o5ZFV168HkBx81C2sqnEfo/8zCCCgtvrXw11b6G90Jq/mKhwby
dOx7Nwbc2Atx7o4HbkFtK7Iu7oYxV6+Ad8CN9cJRcsxEKHZXaMb85L6MC5zc2vb6
ObTG2q7HQ9RI7Ro9yhFVHnSoOV6KlRFWYrF1NDbLLsFTgepXSBbd5QktV1hsuEWp
sK/8Olg4rKc0ojM+VzmaPmPq6KsSM+uthQvjdLFkLGpBErlLzgSB/AwZ9jq6QrYD
999I6e/Sxz652XHSZivfUJIvSQ5k00XiUYRXLop+4yrG6cZozugF20IBJbGhb0Z7
EZuSTIgKnAlqHotw3dw1tFqQzhwbVeO29pVjkjWiHvSqe49LYu0mTJ2fi1jx9vFe
rfQus327oMfZnNbAmkWCS8p9cGqZlnC0oGZLi9i0JaC3vmCro9glAtK2NrpKDTkD
1spLO2bq7p8T6+geKY2JuDWVT7MrzlBVTX1rX7WmDkBH92YzWLPR0JyW5iZ2FXrv
yhYHXnKz8nA8WW7jaEhX1uH8T/H+TbiqTFFg8rL2iMauQ+DjQOp1U1pIJyDxyfPk
gLVa2qcIRvEieYePKk+nVXpDgM/8YMEBxLtsZ3vFMwiaKufcR9XQ25Fo5aq5uKGT
NU+IPPHR0uJg0o0WmUMdUyh+JEk8QKNDDVjXsaIEL9ASE5TJscnXyVUqI6cI3Q7t
Ls6Ix7+ELP855lY2cAOdbELDxEHy035T9PAQ4pPPznPlOgjwPtIKfGA+qUM3YJc7
jZmC8sqRrXyYebFdGaimMk3gMy9G6QVag7rNJwRDgLz7JwFAryKqKfCuOjnUzFXS
O0IkLWVqAxlk/B6Rfef0Q+keXzUQU1MzqRFplTf3Unfg+mUAwefOrBbF0ZWe99gM
W/KwmEJYTl5HiHyk2jF2xqYx4QczuA6DDChl5x4dInBEhz9OKe7W36TZVsW/5186
RW/UnhX8z14Hx3ctmu11de6fdSRfNgn5c4ihZ87L9isuIvNQ9BqgrMvzMhJOuZam
hw0jjKAT56wuardfAwsg2MOKMXmQ8dfy4G7ikh6aRPEeqBGnQr/28r/7uU89c1iH
yAclTc93wAZkg1to6k9qK10AAaPSDzbn33Al+/69vRGD0jfuxmDolnTDh/h/DPzX
sgl6d7QIKOhmK2FSzfp43zavvZkadf14oz+C03ogBVOWV7KH1plTi+j6sXfsOEoc
2HIUp6xY0cFoIMeVWgd6ohbR5a8kaZWRSl4jJG1cJCPaXxfNg6ad2w4o++PGUfZj
RGRNfpVmfe1Hp6d9OQ2NusUxdy+JDQEHscMUYL0VQxBnAF4nqKHnXKhKLYH4Qbj5
WVUyE5yLy7L0HN5Ha/oabeHdclqDD4+pJP+TpS9/fAy4e4TqV/LwOQ8jCB9zn4za
5heS4f2Tmhyn8mvw7VB0ZJqB4BqIbrdBVMI9DPl7khrdw5y83BsXPRmzdGCVhHxw
pylMjEsBrI0xQzXSX0FuuKM8jjObWgew/YqzD5uEGRMqF5o+JWrsz5aNLZyTb4Qk
1VA17Z0fFce7HfesaDFxIoyUS3yM88whA9ioJqCBQ8a2pM4PzXBKHV88ihOin4ms
BW12AkAisuqofjySuAbcyeW9UGI3x1lnFVO9ZM6sw2h0D4FNF3vz1r2Zyf6zVOsP
asO62XHBUWV68mUfqg9tjSQSjuo+JoNZJuvsF6H/P6AI/PfzrloUUpSQIS+ttzG3
nD6scTsy48WcHrhfCOzIuTT+NHXfu/CMpC6qIW1TR5Vwqgp/7OrIpcMH7qHJ0NYl
LRNB8pCB/vufgQx7E2rqYxTnRHrGeTyXqEpDrSvFfUCFepg8XyptrqlSlCbGSO7+
yoLIgC+BJbnjs197KxaiuDv5xtQCjfavO+ozSgSFQKx30kXVbn6MYfYSEUQdu/aB
T9jXDczaT66Yjnc5ZbFRJnumChEIXY24h5TTAGHwybQ2uIO/iPdAMGHfHCkW9+qG
adhZsc+GI74GNO5uZM8JZrKtsJCjCzf1qRsfwquXe75kyAx+l1HdbA/aKDqKz3nr
cAni87B6DADbxwbXa6Dl76/7WaPH14skYoLtF4ZqHSGJ0hPx2f1n8xI406FW7S3L
Ltypx7B1ODOkow82xVzuNbp8+/gfM7uNM8OlT8p/7u2HhQWwm8/8arbqMKR7MzVt
czZg/pwnPZB6Flv4nt81oaLm5729/jtc1aLl8SuZhNNqRL/ZA1FJikZy8P1ZZpXQ
Fq1gwguSAnm2P8wRsLDvw00ca7+ZutGywiH8pZ8h3GJAY7ETcBdWFrMyfAd0NWvX
req0eQTAHNfDbhdEwg5FbFk1X4UczfvqfNXPgA9ZGoMo8kcZeSyFHbIDvTvCDNzP
6tZ1oBmD2+v57uG9jKrq11VscVv90npmFwArRFEkGrmE2ZIdsheNNYJCuCJv2fvG
S2BwMWKmL6sy1d/ecJIaxkq2Vy74XAt8nfa/juFz4NAcAtDTZlU5a1ikT/q4bsPv
0l3URBUNjrkM9quKJXUBxzPdigqWRW+Zik8XO3WqBkx5oobKtY4aORdP1Px/MnAd
tkAHZ0nZaIAjDHTxFEVJy7d/DOaIt6EKp98yp71dqkhxn2JrIAlzTSon3HljnGLt
3jLbkMRUrDjKiWc1iu6RhcmRVW/ou1Nhdk6JdE+3pZYyP1oSxWy0lLgzAZNVaKKT
mC+xI5aWG9TaXrtnNeHQbF+qzxmbNehx6cwgiAUDLqFtNhIsmV5KH3vLk20k34Hf
T4pCr9QuqL6cAxKoLa9t8EdBwv61tXdbGyiJr+jDUWJGbMfknpzybdIZeiyi9Kft
r8Vaq4Pm8bWiIDAtVSQaXJ/LMakqdqIdELztRPGXdfLEUWD6YeoP5n02jTHd7FhL
89PVs3nX9IlZrtjrRnwYMhXaNOIHf9o0pVAhTU4vAKvW0dQgiBd3O2Wsox6xOZMq
MrCtVWbCP4h0ikbzjRuVsSivLO2mbeF/s5CdJPCkz5iWxIjRsCHNK/T0CU2wdbPp
JGl/X1lYRGOphzEms2St7RC+v/4DCLpvtcQtjUYRyJTUGQDfBFatsCfg+jCChWWi
4b12qJhTVP4xLyhnvWdHSf3WLeWMAZEzuaErDU2rCZqZBKJnBiJPASMlfJIGMUcs
ER0qCODiTHzmDotZiKVgQTuSbbWaHzOx4DiwIkeERVHA1GKboMmZ5ACGTnss8Ne7
yHq2pbO1Dqy/w4ABJGQIO/z+b46Y3rna2Ae2LqhMkNrBwpbUtcxrwWXQ8p8Mdgu3
uLZahvi6vv3BvOZ9KHElmtV9RA4MVEJPUrG+TSXf4g2w0vL7H+7uiabAIZT82xNR
1U6kg9OCyYFXYbzaeRoLzBnIrp3KB4r/hVKt8P5GhfWaNytxofTosDofiJoJhdvJ
4xcgJ83AKgF/p0CURTW8AtHLGQfeI/QQ3xiObwrdtaDcxANHjdJ84JAvx+9bNx7J
xBcpi65kgFyj8Iyrm8E7wIothr7Du9T/JTM6tIpnK4QyuIkcnnyoV6n33eemYlJh
i3Bj3FTMQC2cKILiXYwbr4cQhSCaE2Vbs6GE45bRObAcV7+n2KkzapzAcgTwIwYK
fHi50IwMEzjlIJNu5xdTT0YalKkOpfbEWmauc7LegIieqgBepJJKjiXQ62UOwbau
uJWjMts2QOW9VJ9co5+Omrd+qiyIZDqjTN6TrjYfcbSen8hk7sqiPwakppmL2JFQ
PYrFEWV8qQ4TLHXWEEKA29obeZeMG+J480D/vcAHwNZEJ8fR1CvwrN02x3PAXjGX
t7MczRt1DNWczIkeOGmvbwKdU1aqL2gkgBikNhFIpjbuHcscPEoJdfHv/Wn5St6G
kEl15n8GwOxNj9HIUQldsAvkktiqjq5nTmfPG/IkjJRQKZYyn+quHxI91jXrAjgR
qqefKP4nQl4IGufuRclaDOuhM7D/5kF5SzCGywxbu0RsRSFgaI1sGN4cBP1L9KsJ
2PB+SxLZQgoEpSzI2tWdPwSyMxOMOIFLUWxHoErdA+kpDUE6EL3ana025cAZLiGw
cZMTYk8+3hO+9z7r0+oc2ndVSEdEBrVMroMbQQRKuDFzhTndqG5jtGW05EHt7rt5
fvtLvvRxO2BguHHaQFV5cdYAB0QZN/xbFBripMsfCUW98tTlGSgHDlHul0jCY3Ms
HxvJCYc8c/sYIrlh+10v74D2mMBmfZH5GG+wMsAJSzncxwrKDlcPmnCJF2kU5TTH
+hCkNb20bqVrG3G+Hv1jklKKN67GirDTZYxV/pz5xEsC4T/S7WStaA/LxWZKzJVf
YHKmpl3DkqANWbAcPHXz7//ukyH+KcU0zu8oWJI0cC4PNde+yQopekJ610kvRDMj
hMt1bM5hAGRINPRIMoELeTg1aP5DSBbmzaYMkLCncDTY/O1l7jNBmK1NIH7Y5efj
Mb4qMgRyDPLpXdoBtRzWlnHFFBWOuRseI7nbZDEvBN+3oDR9CdjCXXS2hIuIWqKY
yhkgducSJ19XPmFAA6gpjW/c6SEPJPJvrUi/nxL/JKP+gIJPk4v/N+9m13OXHItY
pZxH3KxmPOgL/uofRGyNPWoK3UMXU/8dzP1zwyInm7hg7F9B6q2EhN0eO3hxsbc3
+UDXTqGbbcA2tYppt2u2J2Tl3D/3GI/8V6hQhxCDyCrKsjCA1xiPvAEFKY7PGjJG
NE9i7vIR6gUAQLptuoWMLZxWUDfUC13UWIs9LmipTfMawl8mUsNaf/wWtrCKddKx
p3Hdd1VIh0kqfH6Y1ypV9TEbunuWe6IRFZgtpuqfoSx3Ll3ICSPXbYCeulseOEBU
cYlNAByrerU9JoW6YCnRxPW+vHe4WBd35/mm+3X58vI3KCP64XPP+rOubGxNr0g5
K0VnyVpBeU7s9nLud5vGJrN4KIRXACHvMhABpfW7puyhNnK2Mw5uGR9SaVxn4wHR
lrt4TDdiPptQ8y54FeJy+OGcgrpxZU6Mn+irZHIbMUj7g29/BXiHgfR1zoL/jMMT
svPe2oXjDwY3sW9YeH9fBi+k5PuIWP8JzuP5hkvq2gsYdVoKSIc+a2eVhDjv8+3n
z0A0xnl6ec5ZoXVZA7CPcgIOzM13hfJRCOAELeySeOfE28UZ+SuTtc9b9CE73Rz8
HI5MNpFJJTHFsmg8T4iVvH8+bRWQOpP4qmMdQXbijJpS6+rlCrSElCn/lYWKMG4y
xp1kHC8lTkykd5XsJC/LjrU3sRgX0NnAo0zDhCMXtnaULXnStSBrPkkO97sJw63d
9VIIIzgk63wbER6POtjYZufEEdYKa/HR+q31kXYvCByUp+fY5xZBNoqy1l3hW+Ey
dnBgI6S6hO00hvU9KhQ1mnbLYNdLh0L/hz0pNLYEPu9bBDFvfmjNoWu5bJxZ2eo7
zQ7ogkejc6SLoqmfis6nGKQJjRdctuwLSjFg53kodfU00r7cTmw0dzGVmLutzUJ+
F/bZA+iFoXyPHmZeyX3BH5lZ44nMStRMN+XjHXVaa7y9Sdz265dAexpuTngd+PEI
dzdbGmD0Mm2QcEGJGJSZksIRUMpiTlX32Qg9HGPE57le+XPa7hiUJ+5SrTiNvozr
39EudFEm/D6gI5/zBHD2Cavdy3QKiM9AorIAfiYqwWl5ig8XA6I4Lfp83GK7ulKK
DEFzrJfNxVo3UxjOlnVArGBEb+ROqaco/pX9Y6LNnvIN+DxfNYS9AnydQimD7xgl
lJl6HKXI5EvclXeoFedDemkfnTS4qBOabUuU2kzsF0ymR3vQr36jBFcC502ZJUSg
Ae/jrmhedlOvx4Rfmz1PqPiYeINyh7kmi2Qx6CYHHrxwaXuQLjUpZrkv1Y1GkhWE
bFGes+mW3bhUCLJDClCHMxHkQfy/AM0tQi+GO2EeSkfS3gdALFJfak6JLcNm/OJ7
ZbPxDdfjNXWQusE1UzTvrNMMffLhlhihfcDsGzAuWwrgL+mp7Xtcgs6MRvzsXBXT
1AcBRKOdHstUQiaUXVnTpB0+2izRjW3q2fqPF0kajHLfIAMKrDjzZfV+D/q32h2e
ZMfFyyjManZVsbkgthmmORfMF4egv9x1xnnPlVHdIJrC+HjSzNMtP6VNrAmZycd/
8kKIawUw9DN66T8W/fQjJTLjWQUvO+AMziCDTVe7Qo2TBD6026atbWDPo0bBF/Ir
57/Qh9Y29DZUv01VYB0Ak0I0Cu1N+yPYhDlB99BcQ6G3/VOw7cIV2O1i+X0B4W4N
LUmCESak6CvIVrDheMM1g/p5+vXjhQgzkMLlvewrgaZBd4ew08jo3QZDXZNY4TRN
ZUgF9A/NlfiGkqyfO91XdqYvL+AP3CbBCTYwufVaXiCic54dH/X3ys3ayJxz3F+l
wA9+O/53UVXGbAJJBY4LGqRvWMGL3a7kCb2gNzXWzuSW5YMWuTzHocCY7jw4f9dh
mK0Qsli1YJI2BfFyO6El99PZYxLSADKTqO+ryGkZwH74m0qwq4FXpAVRM3XHloi1
bBbXbm3xuKDmtYxwxz1Rwn5qcMdluEq2vNsQRxEeIFviMOEBJXtllVDnHcwh6r2F
tyk/jLl5L5jhHy3S3gu1fr/vPTYCMpQQe3Koa/XqYhZzCcW0iyvJmCDfEMMgkVI7
VRgCgCnBQAv/FpGpRT1/w1IeM6cY+rK6LiDRb7uUIEssvGceos9rR4dKMAHodiu6
6y3yVM+d9j8GoozPPdjUJpGp8eQnKndKZyAoAXJOmNP5H1HL/0vBvmyGiydVX92R
7AroNDrgxt6Q27K+0/BWICwXuZuMJ8ZaJpYnK13RWkj53CEC3z76fznMhFf7Ehf9
uUX3MfUxQGppMKbjf4NWcdVJ2ywJOdSiDETZBQgmIjkBIi7tOuIkCPj5JvUxYPd9
De+8NEV22f9Nk0pYLkhDG7KAe+XwZOHS0yB6jtp8ESAvKi5khLud3C1izGh48rpr
MNzkTAzbinAJVkkmjyCbr2eU7jSZ/18DRUNAQ65z/5x+MPsD1skKYtsRNIZvv6MY
zOOUGIwmRHtNvQ6pnBTuCP13ZqixS4PbKeDT3HutAX+7VvVe+XSWMiOVzk6T5Kjk
BAr8zvO6MFOHe+HIY1upF4+HRxOLEh7CeYMabGac+52vLv53MSRNhQhiLOph/xtR
LHKIHpTVP23JU1SYBYCnGvyP3hTbgOTqczk8aEfxTeqqd4vvcsNrSaxQwX9KmiBG
s9IaaDZ5vIu0vZMNVv+tVmYIKUB7DCJfXZDJlCA0vVRsWaYsgv5cNmhjVKgeL6yU
HSmqd3PLEAfJEa4dTmlOrA8BJs+dMGRNn41J1uiZV5rF6Cu1O1icmE4+97UV2tKd
7Mx/rt5tOV4Ur2eB4l2uVxyl8fUOGyswc7+6xshcd9hsdEfB5c2rxUE1yPwyaWxq
0weDLQBAyG3nkuZe+1g63b64S/5mfCscsLcLGagrJ96zX9YQp5CH05FXevK60gcH
3Wnx8I2arlD26sQ+JidKUpXlhjhKsMRgLGDes4u5jQ8ZjgWf1KrVLCUkTve8EHve
ApiqPJpVfhIc9q29eDWWnCHRydcgoYsDq2vhbr+jnfiIsnVCEMEA6tEUeIX03dNg
SYvFYW1x/hpeY9OVgaVi7L3LGo4K1oYlxZbuYtdBEAWLs/dpC/1PvJIN9DZZ1zV9
sIUCN/WUhlfR5fnLVYSF3Vhq+p/d7BCr4aOcQOxCop1vEyiRa578/qEAZ3bQVVqV
x8w/xZycRhTPg5oGJ0HfBdE0FPyNP76a0NJCZaQGRBPiaJggpuhDds6DGDZYp5pA
ju0MEHNTBfIVTO/BkLnTBIVxHkIohi+cArFsSW9mDBIwngEVCUe6PnAcrsACHdrE
N0j5iPvpEwdVa4F8rPmbgy/4REp2c3FNZ6DzWylze+SVqgY8EnR8ERlj0Vb7SDtg
rLPigEfqxsb0ePIn71VowXTCM8Zlmh2FOAl0c35IK8V6BQayLShJg9yk8sWladYn
S8wIh7eQ9KfnPCQ5kMieKH8KghWGUSoP+h4xZ1VGx929lzWfYxsSLzUaY3dxcL/V
Z+rs4gq3ovuAalj040jxE2E3Q2yAuFVxbWdA+9DuIJTSsvjyJoaaGzTIC1uDg0cf
9TId4iRVJhAJKY0LoL8u7VnZ0Rxjg1eyuAUSQWpVepdh8iOFSKXIlH/bXEMdq27w
lJTM6YEa5+iaTg1SHkIDDy2o0fsd7BZNuPNoo+fGS+TDfK0s6r6zPadrCz5J4AS7
g1gUID2+Ma9Don9dVAoKNFblWTBFcGG1GSOLAVGja9o6nVXptKcGVbgFLlr0VfB8
gsXb1Dlx3VHL5j5xoIKPNeBuVnT8rdbkTmWIEVccHnMqQjCXNn9MMUGV2TVPedtp
pFjQD/4GnQ5oSUyqzR6HhDvlPMCwHfP0IXvcR/j3E4R5yz+t0h60TUXkKiTiz28P
K4x2vm07V0X2y717ByIVHjqoi8Ziqwx2b8K2DehPJr1Bx4cXIayaYlVynJET+3KD
0Y5eJbiycgHBNzbzM0Sh07jgq6LNvIyuUwKBSmhG9F7WKS2eIjC454quVISrlr/W
chjAwgLFJYS90yvWcd/UZvNtcjvEqOnp5G75t7iHbNnpLmIxMJy2n7x/B3ffZraO
TFQsmBYEQGfAxgpvllG7wjq8oFzxLqgxOybDR1iWnwUUtP7kzuELRrCo9RE3gFSq
2Y9DhMDO5nW3gRxvkopZ/PmRJm2YXRFkIX/519UFihoiEQLbyDSOh7MjEsqufVQm
Pxu4C8k9e/+g1B3giFbK7Nga9QjcBvzRf/26GJS7KbFg9fcPzxDFZG5bK8xvWSB0
RYBqTw0hzyHTb3Ws63jnKXkjbiVbfbgqf/2dxLp6REbzrLhJgWJWkg8s2/6eS40v
UZJNIF0TeaiHDMF7rYzvpKVyNYafxpa+I9kihbK3QHigsAAtPMryod18DRhLQVRd
/yAukVj5ebtWhkgdrQl4E/k0T3EIw9nRGxtrmGwlsb6KPvdz0woA/Dm4JTpO3RI4
1/RNMsGOP0EMaEV3TWnTWOyWbyMF0iTG3+WXkqfhDCq1MWdVId3XpyLhvypNqcHj
BvhLmQf6ZiwxrFcKoNJZ0C/MBAlCRiw7+K/HLdmamianPhFX9vRzPhvLs0cxPIZB
t/Pt/0CUG6zAZeJd0U26fNy9GdaskwT7+OGgrF57RGZegwTD8VG/IEwtv+tOLrnK
j6FeKAKtNvHEreaacnMphKQc4QSwfNi6mOXysxuJhT/5S/RxMA1aJDyvhmhKqcOX
J9nfMNUCPrSpKqT/FhVJjUSfXE/EzFPta0E5wpzpvoQqzY5RaZdtQ/JqiMU15D00
WGtGy4NnBwSri7ZymfWeQueZl3Fzn5Kl8tKnSJrOh2/M8EcFWNZXD9z8c534JgAP
iOaKfa9qBwC/USQN2pguhn9XrRIVQPNptbQiy4STXG45J9zjbbwC+vzPXnuwYe9f
4O8QOAQqxz6j6LAK0QzmnANhgjQEKjt+a4J/8UTKIHfsWQGKZXzHUZZBQCtsqloc
77APL1Od5IzNkYLxYQQGgcsq9s0wdJKsdR1WNqFy+EUOMTYci2UZimnchh1oC+tJ
xNjvg1sYhQkSWmm9sGoNgfJc8TwHDGTFd+qLEyDD2f5WNYgvYWJGmzfsXEe+6COx
bNptWqnFuDQmzv9EkEcwRw5ssIInFFfZlvRFwNngFxU6QjbEsmpijlznJoLqno7A
o9RHASjcAzCqor3XOGCZHjBR46hOozJO9L6INQka8AP34bVh51f04vxUdvjHsyqI
CDSGzucjd8icf0BT80AHTZwgZKF5sTzqU4UalUYtzDykCGacJP4fSAysPIDK3anb
toumfXKhN8nK5EMzgiiBEzK6/tWjVHRlM8kwrfYat26x9cwCOIySSr8tUwlSDIlX
3ZnSHfB2Uk27adr8qyy6Hp4e3gKWRNyk2c/njoo/RdijGqxigdKocJD238VOTgN3
7L5S41TJFTzS1I0Cc7sDlq4c90/ulWg4kLCmIVtdA2Qr3PJyvEY0W5StYSkEVAzv
zuEltxOkWyHhvBp0uxA5++QIAn4gZrwYUbWZiJiXhZhabiytAtKrK/5hRlsiPFLb
Ze8gvaBb26x7dUuHraZ+hEsXqaGPtUF0fnGcVfevFuLZs7J0Cg3h8Mt4BHjez9N6
KlyTck23Z03S4g5zLbEzHyYBARhKAozqychwRCm0oywba7p+q8tqkQDrR36WNrNd
rfuyaTe/opeucX2/kJhF0dMma8rdMCgBR2UQxDml+7iZn6gCxYJvClHXKSLDuZt+
+IM5laX8zNbVYR7KLKjvttDtfJfIuWypm4cHVaW3USiV+ot19XfVbQ/FEGDd/evm
CZ1PzJSTazfHyTJfoR8SxiZjMoTALCuyUn8uNfPX2329UFzPvLP05YX15DDgLTDa
th5zmvCvh+NECVoI3iQu0hPZN1IkPu7pIg/8O6UVSMot/SzC8HnHdbDLBnuyA3bP
Vs7QD0bTl5Mb8fntaQIvzhayx7pAoE437YazZq1wJOv2x4vBwhLcrsWWr8OLM0Qh
bfF+jc/Wh/ANFy9oV84+PjN6YJ9Sdm4Ewf2kRlIW3HvRsNbAMSAjkH8uCAujAOA2
4Da7DvXXUwqx2NCnaTqBCj1D4DopNLWyXylwgffSIVCMvktq98qARyZMEH3mK0nZ
gDapUIhNHGfRM+WFPJBJtLZgVc7HfMHe73spNA6Y/8opQm1LllrIjBvAIaiYf/mq
Xk8Bd+lq73DiM5Wk9AWaUQVcCjgVTVKsz/bx8x3T7/Z/lrM3LSMr73bKH2YSZ7Nn
s2DrDUZOlmrlT13swzuBe0SX4x0Dt1UH1TLmDs7gVhqIchDFLgX86tD7vmrM2dcy
7cAXpMjDTlBYLIubUOrfTek4zoHPqur+FZh21JNq6i56qwHZY9ha9LuB+xXolNfL
7inHfp3pnUgXZ1ITCRZxQcXbnXxNfTcRFLEXYnHsA+OAR4nfQrjNCqLcIrl3e+9a
MAqqRECXGUqhkfexljXAqz73I7l0Lmoa1+2CexRDMUxD3dA6vplOT6ySLEtE8Ox+
kQjPosCWQIQ5k3DLLOJZZbRZA7i81H8gZ3r/rIF/iTolKrOiHocFBsaZATRW9f4D
eaSpoWOd/8faHyPR+4DeSrtf3OTeHeX8Z2MCSHz3HtYML3kuSxkGFg1Gk0h52Ekp
I++VbbIdPQAJ/4caprAcXv+XDlH1p06RYWR3lSS5JmZ1Y794o3y/4RS9ZhAkWUTe
xeoQgFN+OMX53/VSCegBYU9ncnu+4TYFG5aqEOj6lCE7FqT+wNExg/wjYfRlNU+Q
3d0jgB6sMGdZqXsAQ+N/ibAPU7cUhcbmy64EWyhYsyB5Ve8Lc4LKLp2EwbpnWiZj
5nwPfNpOs/+bdtxGIS0f+09aGalKULphwOUVCF+sPR9+1NnfUQvyWDeKw/HsZMzF
nSIKa9iglzvLhU+PmeLv8FhVb9Ah3EQhmKXqm29vZz0ZY02y283rRk8db4tdiaBL
QUmlhKkw9z5dlKjGYFfGXFPrr12N7lSW9YetV0VHAlq0XqFZFQ//J0veqaP3hIQC
uVvwe5BbJWkc6hHRjAx0ugDRAw3XTOsd/rky4wXpzLf6p9e4YT5Whcf3fj5pFFUv
CnbqpHXJKa5OWYHEs/0cIWHh6Fo1t7kWIXfXbN4pIMCWshM74Rrxyjyx7cyYrLe1
Lts3LZI6sU+NnvnDEx69XYgK50m3/EvC/aK3WDrf3GicqAARbyN2is+eYfm+mKbK
YUTwCyW/EdsyYWatsHSbp9wOHbJ/D0XvYV7dC4dNpGw/E+7woaHT+RiDt5AU4qYU
XbJRGLw6V31f1ram2tVOEfQr3kjFUnP1t7PLkEFXATzor9ABXMet0JSx3tmSFbiZ
zvUj771/JsU7JjGtE2qATkNtLLpaH0EK+aWIosfLJwr46ZqKmf6lN87HiPY6SQ71
qVGSfJQBaEwB01uLhVHfIZ79I/8xrqFYtUMEc4cZXt86Sjp4wg05HYzIknCS/U4o
i1lg9rzxF7IFuJqdQ/j/hNtHaEjcSGT2vtpdIliMV3L3hkZbNVYAqRI+4ft+ZLbW
BUtyg3BnRs1NyzY+/MBqCWYtUBUYXf9DPrzqlpLphE/Z197MB7EWWxO4rsQa2CMT
UrXWhnZuAdgtVZQSSfB05h73TCkjGIDGaujvdssyIIP8K2i19ZqDkACbTiTtwF05
SL1CSo/qED5q7DfE9dIstrfOlUejA1g776QAzVB1NEt526jHR62j2GvlIpAwIvCh
7yIwRPjCz2EwpzXR0trumVoEVwKPbHi7hXVgWmmL0neH2q6xWk9vta46euJKIsGn
MNo8VwltUlM+x7cKi5iVt2nRyGM2or4jzGLetvXqca6XcQqeeE7UvycXsDUHBE8G
r5Oqn7oVoCPLKzdKDBwgQMoXEzPbsob1cXYVx3mFx+UiBdWJNrIgFQnqOvsdkL3V
WGOXLIhcg1oTNz/87jXOgG9+C0gPmh2M9csHb+2auK3MCWd/cQPitP88IyEroGKW
nZX3/rvyiDO4dVzaFaq0wy92TCJ/sfBfNj2ku4JD8oYncvDhwXkyWx6s2ADCNrYO
Zx2vmAF7cqjEBF3Y1jd5USNd0pFUblYNpB0xVxT+wIxRW6w4hkCBanYyo+qhcUc9
omFJ9SCWIptcCQdDUP0/vYlNdeNVlKBbrPgR/p8BTflElCfpSLMk4Fc477r21HhH
Xab+9gTJJkBByfNTEAhoFRs4dLJ2XIzJ6UoAvSQRyO8RLGpTKN3NJbdu+zsFEaNo
5TAFZCfKhS23PtFJjaKIL+QL/mCYDiuzKI1RoKqfBRG27Fx83pjxTQBVFzc7QhCz
A+hDhhpKD2+aEMra6KwtGJnRrMjsiMYdw129nioCxAUHwZB6k7p466Ye3q3QK+vh
H38JAImJoaaOZS4vfntAXnGSP8S+5nadUbxOvwMEaUexAhg9ylX8ZluMVAdrjEgJ
0uHRpOoBCsOgbTC+4ILvpYUwJ0QE8nW3kfttUMigYhipJhvE9XK7r+UqbKzudiml
kP+jyfj03GKJJGVhNLQ38j13Ri+z6cjkPr7y4LN4BNAfwzrMEbQ5W+1tNOpQCdBT
vKycdEMEgxRuNobNp9ey6A163MPjv5cmnoN6iEAx5T91pRSR4a7RiCyGhYSH5fV9
15qMsl3w2y5CY3lGfqI4IHMB99OagVhhZeg7Xh/GFpdvqvTqfMT05SP1lk2XjmjF
15oYxzAMqrUCoX5FxWN/fE9Ja4qqI9GUqDnzGQHRWgyGLB6RLSvK9UZOdJ6VuRCQ
TFfDSYNtQzxfuWw/wJGjCByTgGvm2kQOBi1y2yUaYsXnmO/ZRX8h5DMbfUh6FGrq
98ZSnzHCG3w0ri6+KvCsBS3r54m1ZCszxnJ6ArD3bUHBdxGKDmlPwvoncowXeKqr
0mjMYTeGFd3w8k/trdDfGpMi/VLIH/Q2CQwqy/GcDN0C+34ZH/C6pqwzhspYfDaV
1JtkT+8apJeXIHwvH24DjQJ6Q/6Qq0V8gjrANAQwy3vMwkXVeP4kDlKL/YnV/KKd
Em3jEHLMtrRjBAm+Ng2wBfxA8ddQSy6V05oZ87EuBjW+nNONWesmNJtjFQLpHgUq
bgWIQlDI87P8hqzMSUgGsOlvIPvbDUYLaMubatOjl9iYrCv3DC4l1GX7iLDiPsoV
qdTZ7dRksnkQeJNL9P6n/SgxXiiSEGKsWi60osgqPxUTVN1hSNEkxeSManeWOMTv
we8xUbAHcG3vDfAA7VDWRyQPihST960QBmOLKjkz1appllByqUjP3F8P0v0iP3+3
+ugEyM30Npb7iTFa+zYJuFVdkYGfftGxmeEbDNxsah8Wb5vPZtdDLbrMIzqWHjrU
/f58Dy2ZcX3rQpcECfRPr7VSjau39Gnmf/Qv9kwcsz6cgxwV20SCM9G8TtRfPsua
OdbhT/0q6rzVk0Nqyiho+b0Xqt9+S2g8i0/SReTdQv9FOJxkbfEfjjvICeCrqjHm
ZISFEqcMd6jXkM7nKaFtqz2pvZrpnX3L90SnBLWCiYDMk/avE5gsiddVPLLKui2c
GfDUJ9d/iYWcRKqu4qXDpbO2rQXwuArA4oaOrUyAo7jblxjMQCr58xSZpuQ4K21u
h59tlFtEJLR/zVoGBNc/0vBA/bUU77SdsWcNvE709NE9XkrUCBVEIlqA37Hj7mxa
AJR4cfzJkcZgRKdrfzKrnSzsE6caulpg199R9U295rPgxGp4Erx9b53vKcD48JcO
oyb+dBFs8F3Zps10y3kSiGIi5AGCv9pu6WG8hexv/rYqDT9nBAIaEJ9gh8PN/5HF
L+2X6m+4Vecf6LyBFVr8RuFgwy5cQ0VYegMzZXK5joxzzJVyMorQZOSU4BEZwUuV
gCWke/M1m62nKEwvTW4Oyq3sMF7t632acEH5wmjysHqmPeZtHjAEVNtFYXKu3W8i
0HMGvd7vhFRbcKMed2lH15LjQe371zfvtIhY2ySQHxNpLwoaowxsXvFuzVjBjJ1K
n06el681n4+ntSPYtSLys8a22NsPjATPFR8tHW8fyen/LvNYUYnjFijafTvsa1Nd
HmF6ukHgEFkdZ2Js6/bSNDXTCmsaEASiPpNQsRpT/f/G/hqH+z14DE68xKBxDE8m
o0TS6fbVRm05JqESlgTtGiTDQa9QfuS3+iR23cPNfDAtdc3b78OLPBo92PzCL17D
d1XoMoxVdg6QpqC4wcYIGOPw5Aj2Zv6fVbusy76saxQ3g3lk0uvxrQOw50TRYF7s
YpcsBP9wX1N96xsoXetireeT0Ih9MjqtqITsHpqJZUcddVa2ZOtS7Spe4+c0H1g/
cIqEObX/QCqYPBXYOkpf3HxkSeuxuVgLACrX4V0oH8CVWP4zbpsif/9duE4wyHE+
zwt4YV2XurCqaCkH8ehh6FpuxYRrFXsnRIOFykUq1MBjOxpTSIqopMFSIxG/1F60
zfiTf7fCNhHLPzLsOYisuKeYxtnth/mDcEnbDxcgDt9X3eN2Er/0pF3eIFLkgLzX
bUyI/vda/VZlTcpXOtIbIlxL8PjIMDjXEnQa0gl/hCWeqe6U7mZDR613PFkLIteW
JjEoFQDDTmvMCCO6NH9GYleqKeeNjaYeUky6d5Vzi1dzWxIGlVT6w73cid+6MMon
EJ4LW3txANcWMQISALL1CfcMSyKaWF2MV731uHWlYOOmeKdELISNIQ3VBK+mEM5D
2wA1jro5Ycp1uESYN4kbP6RU/u5SW2jG6COwkn38PLQx83KkhvJLtK4SwzSlNg7o
3lCk+mvo7S1xIYn0Jubsy/J7oNARJyLcaxsAuOIrJpDVlBR493HzMGalQIZ7kInj
KcEioqQ0Yx3IpNBnZfkxnkgEqJv8zds0l2Lfpi4I3gzJikJu6pz/KMakQHPGKFYS
wV3K/KMljYzxGHr3e+Ll8KwPaR3lm6o+dP2I2dTrZOHFxYI3xjYyxlmJt3ttiw/C
Gd1TIB2oe6HR0nyu0qQE7DGqxhnCYMqlGr1G9iLBzSmNb8Vmekoo6vjn4Yfnm9lJ
Tg9ix8vZlwq0pAEcNAl15jW4TQBGVliBjxlfpOhyxFkhvPh5+A68B0KGYAeZRasb
EM45qfo/llgYL+G2WLMoHhUagcoGAF8A0vpY/3Ryw/5e/ID7RdmVyuy/I5s5Y1B0
ZJekrynTM1Ggs9RYmnTXOiEow/7yDtxtwTsNX3h9lawXpDei312vJwE7HDcxnIIw
Npaqn0Lj5C1+mUJZ60weyY6Bvc0ZH86KWe9zMIX+BAZTNW2KgaeXIhvWYwONZwvL
i62n0sdVRBPmO+80QX0DsP0NZlWu+nLlunqv+3ODe0Ac8TbZtUENyLdBNtIUvGwb
sGrndICFmO2e6+xlJy3ktjIPBmrpXBivg/R93Vpex8iLpPteUdnexE5/yvtMhNHQ
Dzndiis5y+eNbtD8iBw27JWmJ/Om+mav7vXIEM8v7JeHeeIj+2Gd2roNqCJhNg29
W3LjuNmQKFpSs/Z/OuB3VdqWcjCoXERI7kzPqoE5G7/UGU3YsXQ44ZbxucBpoNlg
1z6wE21la6PkGwflAzJ3HagQ47IVN6A7u0D6AmIojoe/+dgMYSaMKpaYGQmdJ8Uv
MVxPZR2tCPMdSVjNtyZ/MRdGbX7eo5KkgQfs5Y9b1FZrwsXKREucnpTWUMNHsCEG
1Ke3n18w9jPhDl4lnXR4BQXFxllA8GHdNGZrK/TC7nhDGdpWHLH3J+t3Fp+wXgSn
naZGPlUKCCEmvUSUyA77wnTie2W/+PENxiAiKtB3at9qOB+LD37zk249fiVAjANq
nzElFfLC1DAeXu+HXmj4VQ9E66zKYiN2QOIH0O1N5kvpPcNR1tizXTqI+gYLGqh5
314HQvjCoY4N2oFmQbGhEnk1sYMFJiOKcbZywc0jSqe1uoakQ0l1t2o0FBJ9KKAV
l+CcB2nbIDwn7vKwQV0RWgha/sfgJac/Yb67bF8l9uCnZFPASgqjLQgNyr9Pdf2e
2q9cp2CdLfkGtHi0pZZlCHsWx2P7HEUxtw7zHRlKhzbDlnPfxoUZppuY0ikuqiAI
c4MM4z7pjVPlBgypgcFl9nwWoBnYYPLjv9ZhTZA1lQqcDVJI1CwjBTcMPpvUQYMk
0sybk2pD1VB32GnEvndrzrS/o8X3W195TLvpcyT2X3QrSYyhXVRezxa6FctffHDW
bL9fO1wICXXygE84g9+bhTmugfGDimkroFU6A7yKW2UrSLfv39ixFGwLU5yvMaSX
MApJATC4OkqDfGgL+59EPif4SUKaUjn2qR2cKQ4eMD5OEsl0F9yP8eSTCnq7F8sZ
R+4AlbTGaScYbfqEo9PKSR185Rd1a+O5bcvOi0GXM1GARWqXs0J2NmaBfwDmJFLq
6/QX7UQJaA7PYSibjn+endc4EZFwjlrTdqgoaGM+VCF8rzFzu+s48cMVLQU2/Lwn
LL8KKLZAjG/ddqwegWMZlxxkZbX/GqJ0Kry6XXGgB62cm/4HSEQf+9FQnE/001uW
zqlEargn6H0yY1GrUBv8wBndaHtPzcaam8rzyPweSIadRyCKPRr6NK2CqID46QGy
8WjSdNCQyyuqGE+jmquNA+qPXpkQaQ8epbPhySUuN7nYM7TJThCqthFeHERIy+1X
aZqGiRzWxMFZAFBa33aBPCSDwycbr7PCs4gYOHLh6Cn/iWvfsYXTH6ZJ2zORo+Yp
Tw631p9IKXqeMBfw51EKOcX9/hiybJslGOZIP7lficXeyp65tuK5OcOOdZvuhT24
6WZhnroPw4v23DM5KrHfljS1Ps+io1WfL1XerXWLePr/1qwJAN8bLiLGqrQkn5Cm
dVmFTSNBL3GyP9uF9yczqEvMTiwCMKoJSnsomvXei709OMtz7QON24jAaavTMvz+
hFOUBKhG3HPhgpKaDLpH50wWiRY3L3E904xJvetutOX35f7oioMxTc/grWqpSY4q
9B/56vXkxQ98yqzHJcJrhBTro/5ZQRB5BC0S+zrlUMH8D0ujFF8jZugaMlu3OCrc
5abscvafFP2UcZhiYjlZ7WHKml4OMMFqx6fRQhJu6QYcJ7Aixhc0rfAiIBN5ZIwe
Mc5OdjZzmOia+5JTdIM1x3io8lqCz0NPZWtvRUpfYNkVWn2NCXXj2VingT6dSLxC
q6llM+ZGdVT8yTIPsZuAZPvMhDUdvaz0GWC9zPkWvU1vAfQ8nT8Yd/OFl/EwkhLl
em7ncJwoJC9DMfuI1XDd875Fc5uG0wAX1mC0zcj9xyxG+PRgNjfyi4y9tnKbHG4N
ZZzuuy9r4651zEZsS7KQaO3tGIr8Tzs8I/wsbYMd6bnhtPJZNWIMxTQ/Hw5hJ7Ll
Gv2JbXZdrqqSvNMg8qkx/6MC5nloiQKj39IahStLbdBlzwaqc2Vm4CEND8qgeG+u
riE+ocxmqlfR0EwwNOXap1+kvIBc/+gzpTVPZdhs+TA0e72u5NO0pgFNuIe3V6f4
FmZt+RCyZMKzZxzR2i9MrQ/fLQdtf7eW+VQoetZ6FpdAiiMXZda8AaVzkqn1PYVU
riIRKZ89J+XHmn/8JopaPX4n1kctALOmXu0KQDw8V/rtqv3Z7asiNsLckhBZv99G
1581aiS6ORh+AgxeTc5Ydd/08LDZPmfhrCHVaP++TLiW9jiZFf5eZ4iKv1o0WOJI
n1dVzs4C7AMmSmPtYmtjU73FDjZNXFP3YWDxsOPldSMQedIOXboY1KidE6+XfTJm
LHLNKH0E2lZBYWHL5zy7Cz0OES2/R3Ka4yUbQAS3yMwgF1CpXrE24vwce9kY8fNQ
aySAWFoVkvqDCPsPZ5NX/CGHCFgC0BWtzVcT4NYyBQLVK5W3+pTB8DoaaVCjj6hf
amzdocmLm9eqJPtQKawNyS7xCW4Pc/1/Ky8ASFKGG1Rq/RMPmFYKN6ef+vOcplaG
wUurILzVs3eisw1VlRhLn1TpN0ImWojj6I9KQIWOWgf6QKubkvQ0KUhfaw8IqexM
qycHRaKTv101OE/eJiO1GbgduARIuygc6SPwJRoSdoVrY9OoBYs0ecv8ErXgmOFF
WiaaskIwXsGA8K46RssZknMEULJUUNkpGRu91TlmDK8W3uhdooNty5pNLCYSf3w9
LVArVIzbnvoVxayFuZEZoOLEZJ7BIHxMpsid/jvoLXxrR35hrCPkoLYRDhsLDlv8
mBLeYWszSzJNPllczOH6e55xFFTn2Rr5Yym8g/pc8RijJOpJn887CjTKKl0zHVwl
qVj+ct6rxkpW8bXwarwgkA3ua+rjSjdz+40E/r2VlFrU63g5A48ELCuwY8gckr8d
8k3XYfgz1DL89P4V7dIRSEbbnRE8A8Z0PXbJUb5/BNQkGYa2Za9qIH56n09wbe1a
XITgEzLUyC9jFArBC6LJFiUcb/N2Ls1/s3NjiHfeZfPeLLPHyJx+h+fCb7OitIJS
Ii+AegnW3PPVhGAGbpnXydTQVST51jlb23+g6tcwEQObs3r1oX5VJgc90n8oaRP0
pQl2pdhcUrYKs1dIpvMe6aSKaL/+4+AarSSakOGOzXifCU4cbpUbQED5eRfdTNos
Vtz3T5RYpJB8NEa3eB7qmndYOb4nOUlQGEuFz1sssdxhjN0GusVS4ixK06eF+tm7
08q3bN9e9JlULExfmfJqq/X+KCaLkTwdw+xsByjfq8VuV26EFRjGRj9+j7OijWM1
v/jLuiSObztnpSmxhjLp1JsEWiI6ciQMbihBUbb6J+dxRE1RCJqmIE5tt98orO64
e3RCO6CcVTR6bcuv3DvLWF8M9Yn3D5b+M8g0ntkaIwJtY5SRkPzIgERgPEw6VK6X
RKaW1TtACDWNfgL5SLCilp9/vF0b33gqMp6BA8G+DPjy6i0+V71RF0yGbW8ggqRC
0DzGFqSXzhpq9rn4Cp1GrCH1kyWoxOX53AZcDiGtAuYSNNmeyYJBUTV/NPSu3sC9
u10gqFLDEbWYEndfcKn+uKB43RKb+6CF74PsE266xwqr7mycyUWcZF8OIHzZt73n
/GrQOsHrMuwSp4lVExWSeSvOHE+005v3GCKwFTlx1FSQF8qoyDHIOEhIyExsL0fe
16aWy5iYzpjeNtK1/cpFRUPE+e6g+BoycYaaRmUITbObUAhSirws0Ve1Aw9kwAbG
C/GKx0dP41FaVjWAUdwZkUkMBu1DvwOGUNT9gfhJg8XIMRgt0pgt57+3n38ougZ9
8knkt6LPdOJvrev+DwD2tHBhVmKw4fHZusujHValEq53GHyaHaK9mhv2NZM5T1nm
c5NhyVDwG+fmnInEi6mMkd2fRxe615GGoI9hxOssz87h/DYi2COV7F7MvwqzoXBo
nCyXn1ZUzKX95n0mfmKxYZGfFrph3FUOUxZ6gf5xI78aJUxiCkDME+1h6ITx2IMm
R9yd2lzP5MFd0j2LaI40ChuN+XPc2icIouIyck1L5tRVPqY6ASKqBtlIoC4zmRZO
9JdXpiPx6uRyFj32NX3v0XpU/R/WjwwQ0TNND4M8W3F0nPU2Hxf9ApjmklCt5i1m
5AWYQz2XlUADaBLrD0MsrjVkrdlYL3PB30Barh8RO8TR6sLfL24R2BoRo2On1zaT
uSmXNeD2qdFWs2pDSmuaJ+4masDeVagMYrytf6mXDxxqgv+mAOP5pQZw2VnVb4ex
Pa9fD7RmR4ML68oumuqjksJiMbVOatDOiJjvRFJGBexQ5UUmeDRVVzCY3lUNxsfD
ALkHWR4BfNyHu97UD8Wns3ETw9G+294b178qTqX6CzvrnLcEuCdPWNOn8ef6iRZI
6bNoW52yxq9VTIvmrHtFqYFMAzzkAFpp0UzChKmMaFFhxK8SIgGH+iwl+EfzSCrp
LIoIHlP9aOYf4KfEZ0UfPiMSOZ9l/hIsaxySDNSEJLS8kLT7R7kHxUL94QqEu60y
wtgcOg+PYCAOuH+7tdT+hy/tJN+FgFo5/jk62iZoinrLNOXGBaBSgyWi2a6EdRuL
QvGnStSMW+EzeUnbxtl9MW6so+clhXIOW1aHAjLX1A2HUpgWNcLa+D/UZNg9upOS
b7nE8R6jMA4OA+eXqvufVR9fBWZ1LDFXiAtv98yMmc1gVsg5Z6oIJZXuhMiry1Ki
9KZwMHJfR9cXeugmzVIw88mxt0/TYrqNDD/1JGO/gqe2EIg5ijFIcdTQHpqRhX5c
ijteycgR/2QewJ9R1jF4uRglBchDM0oascdoDshY5ntsphQMoC1h6vGETpU8RjWK
Y+gPsq01AGJRHtWhafvnq/U9jQL7iN5WbbbcxHj2Itx96AWOk2zdc1tDz6r6dZcK
EEBGhmlk61l+d2v67fsHpVbo4y6dcCaX3JN+LgcNvZbM9UROv05QV9y/b7Lo9mTD
RbfVxLtjStRgAiFOnsxIR5dWIYeeINokVrPC1Gv+tHZ+2vm/2zzsKFzaax5zXmj3
4zYnm64Qi3+Gjs93FF+tXWr2YSu3UK9N0JOIhVHSdS6nn0er7YFkYZTddR+0O2vG
5VsH10aO6LgaUkqzd73jbvsSpz+Kf0sPIqsDMw2Ev8Sl3PW+K0yF2JYHnH1iB/Fe
EtFQiJH+XfZ6rCH8J3JozqJqamz5nXh2wVvosv64qlAoQ3RUtfAR2LbepMaVeJg3
Xj15oBYt0NEW5dSF3FTTpezOMvgHhKogmPj7WFojMlw/5AghahepP+wH3WNJUfw8
E8lM+geDXVU9GU8zAZ8wHiKRGlGAewR6KeWdkHyBYVraKtIwj1AGixHzFMslGM7m
gAMOiToZIGrUL2MzxxWlaJ8lCebkIkCzTwF83muENYtxqzxyowYJifmjzu0xdSmT
sdlfK790NuOeIjF7+23vmLXbHFwkhu9YeJ49uCPsNYE4YUHfMbeKM2hVAmF4DY5s
LkOhcVnBE3T0uXPZa8rXDSVTDMORqJtRvkWToAJiJfoMAYhM93Ok9kHGd/989h6C
8rRH49nTtlqLGpkvzsV3SMPW/dZ+Vsp9wiJMO0SJ/1n9NEeGJw3h+0HIG7dQGD1s
g+BaNjIAYq0IGJ7ThUcPsDLdP9dKAOS+7Po/HriU7PuHMyhfGM1Y9U8RfcQLx+HC
SOeol27MnoTeGCKQIILb85wmm3uGAx3Tro04/b3y5/5AHXU7q50BT/VKrcDgv6RH
ftM49kYaCF3O5hFu8oFi54PjQfXmsvgUJaMmscssqPKTYFv01QAQu0F4QHYlL68K
6gyK7zmAh4JzJu57bn8QP65dCY9PLv3gul66Ih7iYKss1ag13NKXapr+PHX55Bae
KgV8l3az3eQeqT3crP+oVJp8ZC0axhRU0/ukr+LGR21iciNUNAsNRZ3Ba2vl/XHZ
qJBfFez9lho4ioQAvzKb/Cfmjm5T9StT3ERptcnufTZ/LYYPXTAED73z2qKQWcYw
SZAcRiwsZ5nlN3Ki3eqDhiWkG9n0Ktr3lFcOkq9zPz3QfKq0hWK6+Fq8cQW542Yg
FhLevWx57ZPhohLt6sVzAahl7wV57NPYtqvoTRIUQnAdy8g6dGp+20Q3q+EH4TIe
PndunkvC30v/qQP+qRGX7uezE1KmdVJGWDCPsxHKUM0mQDrrVEgtgL+QOTY7sUlR
yx3cU5dUsWs8FeC7qoymiJtUzS2puOjNGmlQAuchZ4DSxYljn1CpnEEV3oeVa+my
aDbH9NwGqr6vCFLzKuvUJf3YlBwM9tWamng3iheoJD0vrfFgFvj8GQ8VdgoBdCwd
YgG76bAAfoxino1XwNsXz2U9eoxyPKYDV4jHoDliJZ0gnKKfvtDIDbxLWw2InLtZ
TFblAVyy/ORrQKKfpp42+XayREK+LRhEM01ujgLLArb2QhjJ2cPcSUydqiIyvfEe
QJ2HUdMeoAZQ4cE/KZywZZzq5dik5z7AvQE1qGyziNAzTx/OimnEd4GD/uQnq3xM
5RGZwP8JrRbsZOrMAW3ud/eyFIeLn+wF+TwjJOTiYyMBc0gUk3TmYA6cyE7Z8GpX
9eIW5+fUSX0fWrXRB2dG8RSuBsmEGGh92Yq/wpvWIo92TMe5Y9d8rfKu4JuuLi3j
jCKznCAecU44wOZGJLhCwh01wdIbbdIeHojZQwnW7/3ekZOq4T93egwOLxhdLpBy
TjsGSDuG00VihPylH1mJbzdIVv8OsPLaP/B8pYFkLkew5on+ve0JQXgvglpCzdG3
q9XBk6D5l5WxEWJUQG0GowoduZxkRThH7B2zDFmVn5d2trsxPdAQVPTosZgEfGEV
Zb+q8V7WZD4tGe5dF24lTUtB1Njhs4V9aD/zsuKimK8T4W1vBDkFo4qO3GbvREVx
R259bx/I/h/gC/l1VXAhefIUgD7KH+IbaxCjKlwPG4BKDmOZuuD/tIVwZHXyWuXO
TLCQ6ag0fKdEB9KR+Lwcx1PZZsSZsJzn1Yp4tVjk0OhJLV0w4gi0kSgMc7lJzfmJ
+zYnodZ7cJ/s31lREUSBPEIHHfVuQXQkkwEyR1BWd85BSZjIyQwXMK3dzFaXgyj2
Gk4JeotNccRJmXAsc93UXS9+IiwYJ6fVtjdGQltLvpN/4CDIof01hZdoIfmt0k3E
OeJMb7vdCd0hM5d9mLj6mXDt2DBHR7Y9/1neBdMPSuLIXOviPSKexIbRO8abQsDd
GQ+gJmDRFC6Siw5cHN/Ain3jjkck4hJKwMKeCFpBGUnJyxbPpHUWQ7EBWx0yMnha
RwkpCBvbLbM3Hwdad9ozoG6/2q9SAS0cbkx9KNmCgj7OMNobTv8qw+ZXcpu/J92k
rihOdJPemHA9oyjH/Kr7EE904Zd4xXAQhhy4kcQw2mfHbijFj/LN2QV4oDU/YArc
X5R985KIQ9GVTklohmLE0igq0yH0fgtWyKdU+ufwN6UzY5tQr/5kn19QPT12w7iK
dKdOKptL4yi5PPwSg36+2Q9FQjyItmDABrDSStfKdCHicVNFDo+QP/QTeMvSWVuq
9nQNY9l2TexGrnIuTanpJ5aFp7yZe0HLo/o9XFJj7l6MnzwuD+wj+AMEmL+xK+Ws
jOcMRTy8xcPmw99IK22h9WnBApOSvQkWpb9m/uqx7aVMObIO1KfQPxd+OK0M3725
diZmK1UyJRVTb48LNYRFna2mE469g3t4+di9NfszI/ddDTEH8p+GRTNpGUiji/77
saMzUqQieDpw3Dl/2PXLABU0VKBRMSvJuS90fx3ELY/ehWXIqwLqZtKfOa3vYkq2
sjbLetlDKdmMWz5QZ4091rJCcwtGh0pX+swNCDfPFBZDhtbhY4m/TQf5c+w0T/b4
2ayOKyKh3slVlSUz9uOxaCemafPI+0I7Uglxg2DuENfvqYRmwAhyx6FPPsskV30p
0PZyVzqWpEwhxZnDzLK7v3U3OQsHzG2/1jIdAZq8phBWiCwGkrw3IuAhWYFArXQi
72CPhGe2cWg7KHptCdHXvzmyK8Ulx+TLPg9WSkPY7lOGoXGODG/VmG5S1EkDBlGA
3Zcw62/1myH/FNADGLuavoB71dMbRe8HLMxdqGIixvOvBeShKRiMMMDFefrJ7+OW
K7aBnio8qzA2YKG5/P276MI1/IjF5HVTmcH13ieqH7gqO5iGz9jhEiwuOEvptSOf
cJz81k+OuTNw8E5cANXyVy7d+0fWvAyA5rNhBp2JIePSh4Wlgv7o2bZaZij6jhrf
ncYB3N3XuzEmCgDfD94T0InMm6yJxVowVMVhRXVPEUTFhjecVqBgUfrnY1WqCSOe
QJ9M/tuN3hdQsE9ytj41rfn/5yZvRtAvV45icATm692BMWe/8YulgYQ9nocPCSXe
1s6boQ1LTMWKwBzkzlisIvYeeYeNXpFw/SJiQcklxFXCxNj6gEUFcBJmwd9YDUlQ
nerQbnMmb+iJcLMlShzqWEzIC/fs2vVV8z1HUWBsBBs9QEkPPakqCarBokIeeAaz
R5cW5/ffj4UrbyIgQiV1/4S2DcbynKEWH1gE/ycr3XktOmEm4rBz51oFk3V5fbkN
wGEfhEUvFvUHUHHkUY79W4w3y7BjL0NcbviUcGdmTyiWVRAFpKUpoSRk29cAQZjw
50BXj/L9S+mwZNuw0697hD8NJleYCGhnQY5Odu6qRM/FitDU6YB5PdEhD6UqLawD
lrLZNzWCOqP1wJJskBmS76Jdt+anXkvj4cyLiJMJgwThnCYA3QdJm+LQC5BDR9vr
6OgeHUeomE1sOqFLZE6W5e9fMy8qedygJ3sfLqawG2TQojNDJbLH4KuEQEQRVo7L
XkoY/8m01/e/3bk6J4sngWxVOQJIfT7wC66r7SshC/7bhJVzDwnpMBqN5WbIwqt/
MHoB1bHIz/P2lCvJ2kehFvCyMzsSnbZzPTjzG1XovpX/i5Qq77GgCH7I1FYCTVdM
XR8fePc8bk34cfWmG5dobIK6gAdhinMGJehLZxK6MN45NAYl+SdT1ut6dAVk/yaa
HMhgz8WxTxXJhHQ6bP3LpW3cDrS5lNGcDf9hJYoq0RnHZcLVuf6KDuY8WDgMJ+B1
AunAMOl2bRJk4WK3GDlykecmqRwA+YIVdxnoYCY9qDwkwv1zCjFmZ61uOcEqfJo7
OSbgWHDQrIXQtC3cgO99yp2Bl5mU9g3FB6/91hXUBWXT05y/de93fRKpGz8lTlnb
5Rn1GlhTwhdQXpHw8BEoTB7gDtBQ3PEQEx0CRC9NNbeC2PyJY+gC2avpBSwPGoGZ
LmebKC3ecYr7DzFzWdm4/Q7EVTdiZs5Ofq76MC5a3kRjOQ7G61y80KfPN18LhXaQ
rzbS6AUsfNanQRj386H85wag6Mozy/pp5hQKLUmlVGhoS8OPDeqAeOQjyOW7lnDD
s2a1ltNqeV73bEB9TPtCNt1oN781+anmvJs0bE5W1WrLcom/kiTQXOr04uvbpO7d
15lGX5znq2yQPHrX13DOq+wvN37JXOsge0skksmc2uE4jLUbOsovdouqDbhbWmo8
zmizlJbPaO1UqqF+zHGBoKMNdAscBnfT9y/Jfct4pyDkIj21WQkLy++HIuta+qX5
1hECt6Bayfk2nC0UqvXbT0LP5YHewBC4TPHVcyStHgHEm4lB1LitX2WJP0QERbY7
zkL3eTktDHz9maTks1NGpPOQhKZpvOz20CjfRce+0FaohuODBc8YtVBk9+E57IGt
MPqfBPU6zunam+Cc/buvmSvtQ/l4SZdikqv105u2OuOMglKLKZfnyZNOKJ76FAn3
pGPiHc4g5B4AC5DIVVYoPaBKe8hDoAT1OiVy3V+1GElomRb3TUI9hkk2CcLiKEF+
wpMeaAE3mYnvJ/+KTbNc8hSU++ayVwhxOSGfhQ+spq20w5CZsvnvzAgpF7E8pJe4
f8p83OqTs4Y63WX6VYYXjI4Ndyw6EWrwgEy92hoEa+zDA+iyxX8Jrz/1YATJo2Ip
rH75+af1ENsJAUlcGGvA7G+PsW707gMI/9c4qWbFr5gyEC9zZnWljhYsMrHjpGpd
yYUAhJte12ptjpypLJAJkAaPRE7HUMA4jbF3w2v3mpGq89M/2W9hkCJ49ik5WhnG
Ja3OKEYedjvGokzF4BHpeGmLSTtYrq14BuKjAAiyk7vI2r0UJfY3gnvQPh4Za77a
71yVlmkNfFiV+hBo/82NUMtXtmUo9Ll5CKYS0v4+Ro0XfzbPki2A7zze0/UNXI3B
LGCmRv61FBwGOVvtBH+iJ4o3kPbB6KY69L5XF3Oo5Xe4eblq/C56eMYxNyUo5Pmo
WSpaWRDp8BiaFXiNSjOF6vylFABbidVhWDHVAmF2YieZr6ssvltTbuzaqzz7+h9f
KRinUL5u84d3q0zXNwsQxUoqhnuA8EfwtxJEiZAvTV14hzdI4k2dPWazrbHsxTOa
V+MybbyDESdI6cw6pFoXFV/5TK+rDXCRpgLrnb7Bc9Ax+0HevnhCG4lxzrzNdJnT
D3eRW7ZSOUO1pbFczg0M8m/LbjCpWwHmzQElugvAk4mqOSB5Z9+GkANx0PBHfSMn
ES5c1mlObGT9+FjpHulUUqMLwxpLaauPU8WVLQpIIIt8tDe30PXZlBFEW19ZXkZ7
aXJ882d6Py6PzWyjYZ4uY1bkHOf+Okd5njHoaF1o05+tH12255qS7cJfMqnrFn5k
pHsuuvyRhcnMTANSHYHsni953/Q0X5soam2xj6NSiclnqteco05cdgMWsU5VJREN
9DvfSgHEpNJ9MzyD6YYMHwxwt+vreqMeUvgDocOG7G2JCkzUj9VjY1r+rK0aNAUS
w+DsjyLVQtRjWnR4k2TPions0b8mxQNbgrkkvR+u1B9/PDRIsjZ381mpRMZlz6/y
z0LOGoK2v7NZkDemEl1XaV9V1yq08z+xFHh6so3PdZL+R30ILAfJzT608lG5vfvf
m6xIqTJ7evmvwNXkH2RJX+Z/MwooEAfA0E3bLiks2ARc4iUZ8dY1D1FXxZ68ejMd
dK2L9drpZGintRXlCMGSvYAc65bLgMTcEadjENokZ5PG0urmW67kZBSyv8PwmQR3
vDgVK3ZJaaJLYKDXHQSk7AROWCkiFxk+Ghieu1o7eqlUrqfLcLhl1dH73fK30D0Q
0t3gp+FR8Z2eHJ8ibSeFPPcdRPqHyzaPbpKEm7ZIlpr3kipbgep8eizuytZyHohK
yacrSUHqldSoA9alK5HrdEtb3ExzHugGn8LJxTBfgbvEDebLf/j35KQE+4jeJBP5
O+CYZsbF/IqE6wnRJ8AQaC00sf54YDGj0YjAB1Fr8Q3C5WSsnmXsGQoKL7FrKIZa
43kQiO9OTDFjUJVEa2xr/eJPru0B80sBbGEMWR26hB4JedFDkSmVNUOXkfIgMLIi
EJKdk7jo5UATG2IVeuXREPLdq1I8hVL7YeqKC7cnWL4y2pMo2q5Eif4RzSeC5alI
FBffKY3y9V673+SaJ1hvqzGjlCPaAKYyknNhzhwCjsIfLPpe+t1xRi1WmVLp99Nh
O//lQN7BrT5N44sz07n6KvjrEiBGKNLJ2ILrDdxGkAy/2tPi91Wxt2LKq3dpsom4
LYuQ7D4/FljZXocFIDVFgMQzLGZe1vs0CmO/gxm/WE2wIunzCwrOKQ2h0e72J0gx
pXwUGEyLERTL3K2qbAK/crNZ5V7A+o71upWuFBpMXf1bhI6/cZLd3VrpP81EZkoU
UIM6fYTRFmsj+THKWX08knDicmTSywHcL4uTSCnYVNyLkEmBYOdDDH0AqghGXlGB
ZTdoenAOtnVQOUKC0BPI3HmSaBwbN0LrNBiJXNpj1BhcJ0tLQlBa2MoeLPtwpby7
xFHd6kiBvhfTK9g659ixjwgXptyGzn5xChqpO2TW1oTlOWlN81ZQnqn11hRqNlBA
4Hq/Zv81oUZIgfU8qzBcpxuLPvdBD/EhTc3ihBPevJv5LbIqLTPnK1+iv8HQfgIn
8xbYiN1bHTCiHckj0rlKEpYqS6TWmGR0+33khvPW4OP3wIueLln2TqBI6l4n/j47
6E7aXr199LYNbT0cLt/hGSIW05BYAODS36Fw/mNKD9fvdIuNMtWdVngGfvoF0385
TXdbRPG+7ndwa3n39CB6rni10lpZ9Mxj5fzcDi5icu3CpgdBP9XR2FHjUyJftBrj
+ErySaKgdoJj2+vrZ+MtU+tpjdEaNz/u2tJXJIi+RFRu+XTY+wiT5rqfe/6JJwJJ
Z7rD1v2wE5GawbDGF7+N4DVPHNkMopF6/aguqQGQu3RtcNXLP+VwzzwlXWZJvlhi
Pjrowhjj7ZZiiooCZurPabU4I8TIajzERunvqT/P9jI/zVjHwxGLmJ1gJ912vULF
3vKh6SXPP647guvKo7aeHa2Ee9kopb3zA6PbyL9l9Hs+mUb9iGvx0FxvwUERxwV4
0TyulJSfFFcdNsIip4kX1pzBF77SjJY8npf7tkJWPy1CiJiOlU7rpVGnbKlSad9e
dhzA5EbIlz7D+UqSKFkpqgadIHq8SUo4zuOp/WeTUaO6SKGpaGxHRP+F95sXUTao
BIb5AjJP5VjMNfmpYawAMavKwPJhRgY798wsvDhyYgC/tFTD7DSFFqdI3raC8wdl
I3xbNIxJNaFXLGXSW59d4URMeAKeVu7HgxF/Z+roQkZJhYb9Gw4Kux53XXT+Zwao
KuoGXFkZqQ/czrmDQhRLHJRAAB3ohnwtAqvgwQeJWDaQwKz3lRkbMm7BZcqp6GH0
6BRanXIKMU/Kn/k+Pxk/zR6n2K1TJVuJ9GsYvjjpQTniSij8sSsZFRfBnOTzo0zZ
c8lO+GwEHatjHIahez+4rfOxky5hkSM3agF6r+HqbOIBLd2tnY0YeYxmJcTtb6PD
C0DUNs4HFH+EJS9ntE5D89g0liPh1jcJN6MvROcdWnlBfbpv5ONGT4pKKrFTAF7i
oxnZ6ooyEs+PmWXpe+/pdGtbr/Q1TUxTraSijjkmpRT5HHGFoPEJMQfSM6Vyqnii
URuanEKrK/zcwTCrQhkccz/wAZUH/u0IxTZGIShRsQsWuXYUtESYTFuDhI8jOxyr
PYYNY+9OwVg8foEi1J4NuBde+SBSeDlmQRqILEG7NeyBpO91dcbuqxaCjs3kPkTu
iCViwLJeJ9Zrk4tzhhKerTjbg5mSv+bS2BvfgUzy81YociM1rvXSFgjo3vPMfMsr
uChkXzOJguf2FjIesQnNNxAyC8r2TrSWCEMsNcHT3WgJcZCLaYAjwoV/lrY+i2mb
YBpxS3e2iW5KjQ3zLdFpGE6BNnNTrBfeJQd9nozj2XEujyBkxGCyh6+QD70yprco
Cr0/kmcZaGqmGUAqVKBi+ujahQ3X2H2nkAuJC5xrRr728Km/MSo6lsltvnISi/VG
M/YkGl44Z3PmiTYuTusq0AWuJCoRK7HKX1w6nhZ1DolvL0anPAcd5vpSKBTKyxSC
PgbVtWvv7JLGUuE9K6nvrS0x6/qEn/JQGfBx+jwu8yLbd8A4EGHqNJU6D0TSJ0+I
YgQQqX1E5fhyVg8Ijichz5sgHzYfXTw7FQpzE6BrxUWhO8AuDEiw1vE66vrW0H6R
uCiy068OMiJISjzyhWi2yphxeyfMh/rOWZMp4aUakSoVNAHucZK9g/4nDVPZ5RV6
zvb4LFnvMw3bPmHL1OGsS6/7HQArv6QX1ZGsZ2dG3EBDwngJAJmbBTBxS0f6mPjt
daEoIH2nKuKFX9EZsP18u3m5LY1hq5qgvB44I3gDfA46sbFdzCc60fdG8Yfw0Ah5
g+YTDw/FkOQRgf9x3kddYZQ3rIcSdQbNniJYPeGR297L11Sip+OU6M7S1HonJIRn
n5WQZTK8UomRleCiPtn1vFOuXGUVk8xbdpfBk366foIZeJOVDykq/SJHIKXoqitl
so0FvqUJ5o7W/OEo+63mHV4+TbUsZPjzshdcMbEa0aRFcQjbFIHm9wt0VZsFA7U5
J7NN/ErbwXtTWrDyo4JSTHXrM+k3EPvSocj9EyZp3/mytrLI9SE3V3LPQzHWSQVz
dTP8ELbKw+Es3+xT2xyzTN/rcHA9NNP2zCkBnUyvdGFlWC7KDfSkZCRRaR3kmiIK
ZnHo3oDSD9tCx/u5xO04mQ0sEHp71RaI8RKpOqoH71m0SNVUwtmnu4mLmRBl0NDu
dvauyiX7AlRB98BEVmZRarqYCtdHvypLiNU0j1J66xLFoQBORDh55WnPZNVqpETW
ZTjx7C0VcACNrf0Z1rX4RQvh2X6pRgY5s5QJSwtj4LAk9DnlqBmLvQmGGnxP3Z1r
I5mPRJaTw0EYdcftqOXkgCdW6BYrq/+XeduaXK+WUKhozUDwpjgoTyqtKeJcR33+
HrZeVwjLBSl9vAZ0LH3+raek8XEH5RIyc8RdBqGvROzdd/jpq498vvb6CCFuDMcR
MwgI5q0FjlUeVIxKF/n3sBWTbtPV0YnVSom5i9e7TveuFP37bzbtVc8/ao3cCkPJ
aj+DNwU0kYx0sLevvIFE2q6IsYFeGC7LzLdgKFq2bv3gq5xRNUwB8ohK68yQhVZH
nlkDlSc0NGilDIqSJ0HyBU05ORfhmpwF34qcxHyzsA2d8kSn6McSFE4ddbkFbjSp
UK5Ok5IovcDtstRh0Ut4oqyJJSZElS8BvEg4riN1I8nulYWpkmFZTaKdimy0y0qK
edo7gM7D4KOTGY2bTQXqBJEHrBRdob29Y8nO0V06/X859lSVEa7gE4rnC01dnA3v
x/+K741nT6DCiwBtWe3daHXph9WdxRNNZC8PmHS1GkGWGpp90x1+9W9HMk95dtX4
ZaXozET4Af1N5xRC8/tv5VVH0LzNaadFO20ISkwszRbqfOtEodm5D85IV31yLz1l
T7bOVFE2AbOkzzFYe5IjhGh3alfKaYisvSuOoDza2EbUE0OYbnSJTbckYFoHTLqN
1cDsKgwoP0wiYLdX/NeB+NsNOJAxYW8O1Fh0gIyWSq/XU6YYpgIb/pRYZZEk3kRf
957tPDjQY9xTK7ZLii4sZjKJSPtx/2bFnXszl7EuMTWyGD0k08tLxO9p7IVLTmxT
KzlmLzkE5G291UTE+vaj5EOgW9mHHTkT6Hd9B+uWzmw3k7I3QKk3je26r/13BKGz
Qp4HQjtDt93xqBnAG7UVTWLq4JQO9NsQejOfqRz2YoFzl8ittqUZ8Xdjy217hEYH
AcqMEEodGF3t/9W+J4ncTYB2TaovbKq2MU0RxWuBxe1PtlIOBoWGf0vIvskhdU/A
jsRDKXWxn8+n0uEG4RaaThgrpHPKBZgBiPwZUj3EQEvLPBSqssElnlDJTzwBGnVB
YKcPE5qELqM9r4VX0wxzCsx+dkT4hnRSrwb6JH0uCena5+XKXGpn5mMYSQR1VdbN
dDwqMg4fdlh0tSK1JClFfqSPMJPq/NCKRm60oH/6JB9Fm66fSYVINRU+V4H/oJgn
sydFDVP6y10DqSAr+0o/uJVkMSCilQ09j3/PnrpyWkpGCIenMMZ4DrxletPEn2P8
SY0Iw9j+rNREqZg7jsiDgtNjztvSs2uPkkJy53kH6ye2mUUtzrjIxK5bdjxRu41L
Vi2wYZ0OTe1Jm9iWoUyvgXUISUcVfXNyqjqne40A6hNxIukqDf+spPD/TNzVXGFo
aqQvZON/X9HQgbdm6o+tuRe6DiJrWrExbSfyOUDS8IXcHDK3aags3s69dfiqyFH0
rTXAtWnxiazkp+A36sMNXQyiOjWApZjZFD4EadQRIRFPiNthEQ45N++Y28vxUsNL
6BxyXfjCEGWNt+IH9proiSXdOPx3xbVn3EEumfQDryWNWbdSSwHlPvqnkblS9lMP
VwyDtRONu5Z0iY0nVgbAMWQKjwKYmMuFi0YE+KguMFz+ZGmphi/+zxB+PregXvy+
/c8Lg0HUsxb9ubGm1NclMsizSkH+p0IZYYieFtqr4BH0hVdDmlzTcjo5xnHsVW6W
0zZIebvQDnl+QwT2Dja6L8u9ZbVTii/cxykbZRiKau8aEXAuLFrnB7Gcj/YQbJHu
FA/JrZ0KX/bJsY4hmr87EwMPkfylt63mr55M/weXcx/3RC5RuEQi1gjSO98VEo9A
1wFeU03oM2/79/hUnH1MJzF3N9lLWj8xwWOW3j+RgHvVAoOM1a/x2uH8AbZtEnRq
TylCcQL5WSnySzIBjLJ9xNt3hd69xzkFLTFqX0WriAxjF1Uk4DpNANrPWJoMgrK0
qHzFMBidMz4ZU7WWzQNstpQ4tHPUkQy6U6LY443cftwdX1QGk08mvhulDsQZFMNy
511UsWJnssP7c8ZV5SAbsEogHJw80MMkmCHaMaXSIqW/j6UUHOyVDX0ayv33OqJq
g5XNiGLfNKMS3MpsScOT9BGVNxVqSB4gpCdjVt8PdlJ0kpLYyHcX2dcvrdfj7pY6
GPC/ayjvWrNcbCmzzqjvkZb908y2ZCXQ2pYlXUjW0qmCpfS9YJaBBbhaOYcbqN50
KU/tbnFJbDRq+HSv8iZgyUuIanUJJEoKYyQmB6/VuBqg9G/aBwVndPNSXW3jII99
gikvC7mO0l7iJGWbBok31jQnzmQAeuqGlJsz654QZSJeaxf7125NzYW9D7SMolD6
GIqaU6g2TFSRoAbqX+C40lD/2M7Yb2uKbQw3MqRki6K83k9CybrpNN/4jqD7szCw
LWaVqG1//kubERA0lUwsCEy/8CH7fsg15MCSxA9qg99YKNMjm0381TeclzkNIofN
UhX6TNuIPVCa8hBvy2p9C+/b3uELgMwpWejujKeUDBoiZMYw5N7hO3PcIuJnkZo5
qeO9+m4n9NV9iAZWczmtC5fLtazL52UaAubdDn88wFmcIpXf93NSo8RcG9i/pMiB
LaeeQHGBDpTYOV9ccbZDov09oh1eyV7S+znCPTEPmsN1Px7VU4+f17KoUdvkZxpb
5CNfP5qKiPYYRmuC/2O3vSYpUgdwVQFr+b+iozZWiHmsAcIv9q07+z8xuITuKjGU
UyP74sjdtICvV/0XA1fnUViJcr6bW+JXpSHFN4RxlMO72BSobYZAj01KKlTM2BCp
QEkubq7ljyZE2J4Jvp0T9vejktLmsfoTVC5o8Yx23GQKqv7zQqnqErJzOTs7Ydse
A5UZLtwPYm/ROGsISucnggFryejF666IymMaUMuefKCyfVHrCU0xitdM1arfkzl1
fc5V//91iWhGfoRz8X7SZpuu5oFCX+4JQEtpQ/VvuK3oiDoVGdBhahlkNSCvJyKV
HJIiYRK+Ei2wJ4dnlbsn15IYyjWYnoiNqnylxcWBv8t1QSgwGIsa1MySBy2akwlL
4MQpl8pjH/G/5/bO8Aa8lC4i2XHfUMwBdmOJvXbKAXBcjOze8vfbojX4VMUM2oYw
JFX3DZ0bikHbje6CAZgAyZsTfl5Q8HaxiAlVDgW9nTpd3VytfQeMIySEsH+euVIs
U6Nwa+Mw6dKzIrfSu5MwZNbM9vkw0Y1gxYeNd3BJgogCO62spXgUZ2HL8UqnK3U2
cpOteISDjBSavgCCM8Zk1JAo3m08Bxmu3/4ycgxX6UVOVZV+HF6xPlY1iS9soXaD
KmtCWcLt+Bmur4uxYcy613pPItpKh5LjVkpNMW4fwzuYBirCHGqsDlO4ZogM5cb1
Azv2Hrqeh1MqLojaloF1yOq33t3iES2InpMyQ4GBiXAWEwhdEXc9+UqqEG6yrMkF
lZaxEq2q1qnxpUsHA+L2U7dekzHqtPKJ6+qEH0iFWjfLqU4GKvYpTlGaTfD7E5Is
l0XulYFvIgwcqqfMmIiweIw339yexLoG0fzBVJ7Eo/0eDrQwVlQGCW9TYWet2kk/
8EQ4SEqaqsF+JcOeHIm4lyemQoViWnC2mSSpLH5CxI3+afAYVstuKK/jmjJPu7AK
fDPq2RPYOzLG2PGJlu43EeINfqUsg0svJ13E8lL5XfFC4RJWGrSgQTroF8h3K2+M
SzYfzAmtqSPd8QRvUwZOvN+uhgbtRrNIZK7SyPPmBvn+eb41y4iHa153X5Lr7sok
2zOjVxbhe9fIMEsz6NJssut3Q4W+dTXGjaa7ouWhdfVyzSoM27a6OcS+m9XxSxJs
I6s9xKq2eJp+0EADONBmlyQXWGg0H0iWbsL020hGG1amgYP8tFMgu25+WMkKqVbz
WxtLM6v10g30/cTpQn/eDdXauYP7clgMrrJZeeywf3btlaEDRGQDhVaMq/bCpQz4
O0usu5SEUAcLZBOSKBO3oz0aiRT/DHtP6l0wPtnjgrpI+Frsz0IH9JUsyibcDPZn
/F4UXUuF4snAj9+b4GOJOVZdyOPOJLx2YtSIlKKuDd3ER32IB47oIOqBM+EmRnad
LAcXyLgZu16UVguUHqV8hqEog7lVcLs6Ck3KKFhvckQBWFB16Q0kqTQ3LBpQWJhK
IdestP8ue+9CcMRsCYpYeYaz8jeF8STv0FMhFUkDc7urN7UorCobrhCysGlRo5n/
DR/zBMKvnVTCzLt7gBhFp5oBksBjkUS/jOUeYoto24VnZZBaw9ZS79KXcRlVZgMe
+DIYjBV0wDB/iaZGxkd0A9RSkue5jvcg24pB5T3tCY86PrE1jH40uAd9tkJH/tfG
z2JIi3SmrGZSM93RRF6ZfhScSURjNFw0g4uvOkQyli4JEt0PH4f7kFFoOJGcEN4I
6A5nW/wt5esZjHYOAeGAmLsqxqHsnHU+l1TsJF1oCQBiEhNvER86oi+liEQUNFoj
kBujIc/tnF77SoAj2JxExHoYPFUQhWVTmi7IVCscMbsSyJs9Z/KrlCwZoq+M1GZr
0u5cKpP8xaR6ZUpctKnhhcttY3wDGwxsFeAZVph71SBe+WXY1r7PgHa56PSMosE5
wnWL/28cMP8EZaJ4bMgsUA/q6I/Z5615P7mLmye6p5gAIgWVAs5J6NTPecTULHU3
L6qHYaCKrePrEF9yBbLf0AE9DQ+p9pzQeskWvcyF6SF/blcOmYEf9Z0QihlhMjgA
oWcqyKyt6qAxd1+7RCVJ3Z56ZsTT7A4a7MTLOG1e1WshPAihh5p4VtfZVLsO+jxK
pWtGMeSauRXjRIGU9oD2GYmx8Io2ew3t73VGJumMKNxSNKiSBDhXY4dPqmVV1VzV
5aTzItexG3Uwqa7vGKnCJtqEQ1pJy3R97LUGY1GUG8OBGHLbMLKdoBWNvmprBoDS
7cyz58HnGUEFohgIzhFr7IU5JOeV+DiKy6m4ZNeUjAq13/R2Ourqb7zaFOA/QYwR
oK8kxqa/9C2hnjYuBIuInzeeK37xJ7W9zEQlmJjbYA5kY7zQY4QG2fMainXts8Iz
sNmF31uO9tEMBa0GCOtHc4wYHAxvmfepRRXTNlw8HK/snI1DF6zzKy7CVBOiJuQy
a3rZrIkGxj7rlAvMIP5VPOGqWY0wBGCmVXQKr0xp06Q4XDZ2laUGabeu0OTLUwiW
RDE07C72cVy5R83prVQRLvXHRdq1XVkh3XaSB3N5dKF/YQj6prlugsMUQXzYnlv3
f4f96MbHMJkZm7sGQhn01M4DeI9z9oO/qNXKs3ZQwLvt87lEB7Ka5HHG2ssIu6Js
BNfLS2eAc/TCM+/c9twEd5LHmLGEcejgTDLZA5fM9ooOhz2QaXla1hCwXOgeqFCm
F9R/pvAoqFNnWPppd6R+eF9WGHmr1ywl7EYgnAlCmY4nmfV4JHAWM0sWPAb94uek
zR8hkhPdjKAT7meg3g0ZAeGXZxftTBHBPVqFNBpTdgkiCWxhXZWi6e3wZ/x+F3TH
t0IzNLIgepSJprh2hQEHRv/siz96jBuNwoEDCLMrQvGOLaoCI9xN/6whBIzgQRZ3
PNWcHKqIiFlT6u54Dzhggu4cBOUDf5Ijnqa874cgKhQAyiXYRAud+VeRQ/tJqeau
y3hgEo1DeY//0x4HSOXota/qxJzyUwBdMuH4YGH1H4P4m5X+kSf5HmC3i4zKEc45
RRr1Lugrk++8sgh3+Gc7VBd/aPkl8SaaWjGK8SMw+dMfLfdlngPRMkk1FU/KjidV
x/2cCbhf+1Y+25N66V+IIV3D+1P+y9JHipnHmJibsj7CF4rNjYKHp6gADNhCQvFJ
uIK+B/tkqG11au0r0SxbLmCKJ3b/4Ex2AFQkRezfz9AphVB0OS+jdQRWqDkja0E7
yYF8zWChEJaCMQPsdDAobpMDXOb8Nf2nJbDiuWJhVmA5uJPGk0mO7eT6Eo9cXrL4
nRGlJLCNKxHvybriuJLcIMvw542DpHOj4JuyJO7+8tVa6Zv3eSw1ZSLTz8S+1tab
T+Z4pcC/FHXRoMpYKl4sk68gVq2fUrgPY6s7xqweb3BE3Fn4OOeorNlhIE2mrO9S
AHoGyRIwbxWGqz+xuN5F5VGXD8oy1MLg7d7+Rxv1J7NTCge00kscz3SGUy0Z9II5
tqno1n8jBB7KFWKYCnLqt8eyY3kG3HVy5gTQjWDM5IxPmghrnr4FAzJHeIzEJxp8
t2tcpQgl3jVCJ5lHw6GJ/1PwywPxn+EPf5iyE2ft/OXFYcCfAXtPGBDnGtc95HK7
7jqoPsavYarjR+18oS270YEwAIZbvqGrc3taYb27MW9XoyjaYkQiFufprACHHztp
AWt3XFb+sMt85gACwDgjKQn9benNAXdlry/QB2IrW5K6F8c2ol32vpZapkLCt8TT
EqJXFwt95r7qEeyciuoVLnJtxNl8Rb8lQ+VgHqTc5tAWXomLwetL1+IxOBgRfzGh
Xvq+guDAQ39KIhKDdmWV5xCATsiOKTVoDevwdRaKTXvHWejxDqBFGbbYuwLLQeHA
49B+dRBtxDvhE6q7WJnIhtHB23jmuSVi5gW+s2qrHLyaUT04/xAqzx09EVsNDyqK
Nn+Ayv+/TFi5RaJZm9XzUxTbI4YMOsy6KCx3Mt4ZS6ZeSK24pu7tLRubWtKsBV5R
V3+WT8hkrZWO4kFzefCUlkGJRlvf5wnmWyS7nrqzo1xL0Iz2m6t6LqBZ8V4VeZ/m
OEBMX8U2U9wJv0+kv8AujS+Blk8UK4f3bV+sEIZ9oTisvVZlBVBgQlb0FWyJ2Udz
EF3g0og/lUJ4fi2NMEmSmGI+5+suo2G6n+bW/kH56rrTJEyh00+92MZoesClZH/J
vVSEXcAKLN6/KuhORUwXdjedgrQ+d9fPflFwGhyXbRcLezwoz6X23E+5FDYyjPM4
5qJPIP+8nxseuCYbmOXgd9qvMmfFQ0aHBYSAqGMM5LTL1LRiUiXKEHvy1D8L96M/
GTOvgSAyrx7lJ9lkUaqKtMu8A6bl9E9FfhJEY00Vvz0YVYZcgaYmI8KyDYHVAJqh
WdrX4CFm0ydRPDtJnsk5nCFBruoA3qux5Uc4SBsnAKnIvvEsWECKKFS5NKXaraS6
Pq6iktoGGHG3r5EyJk19ut0nl6QtzQKGRPZHxsniVgYcIx/GFHxaRRWnwKMEaeYv
7FI7kvwRG2E/B4MXmPjuPSrPO4v2elFRrJKLKrU2vZTQFDv7orXfuNP4dxlzODZz
VenUx0oieQdHfliXKVrWetpwnwcSE7SK5erB37V/KrmuGP1C0cfglblsby7en4rb
uAFJfnmL5DGQkn0zi+RUjzEycW1Ze5Tlekv+1PRzGAP9qhSvSxR1L3JBv9x0JUlE
niTCQetvbqk2zkOIZupZOxaWFx6iACQHphR/CLiukNOxYwd0TveC4J+Sw+cv+Yce
xn2ArnelOZw293fGSitInoMkLjh5gXzqHUIKRLLtLXhwqneyQwTvBI8Y1BWYpI/V
wHEwHnbexkjM7FfbdrAq0GVHWicHyuWJWhl77mXsNMhhJldCIzUnZvMjtJ7BTtV/
Y3C4TenUGl3fCdaa/wrC/bhDBkC9ml/dJY7q5QHG7FY2P65Ro+k7vGRde4CStiZh
3uPmCikkfc3LGhDTjNKYBWeaxxXiRUPuYuI8JVsHN97ZOP35nnWtXsfitDNipCQJ
GHbUZvbZIKbMJrTZ2Cr0Bz61rHMBYSpnL2WyisqJrO6fZdu9Ssz//MOfUiSSOqJM
hmqiC29HSlFRR/sYh/aBvPfH5dDsI1AJwGUfafCTuqSUcAQVP42S4fK9XdLfW4D5
/yTqIEOoNFF9NgFACK6L3TCpqoTZ062GvstWljI8+GNbwVjuMQN/sSfJMd8dsiy8
k/upzI1EgwJBf+erfyAHVhaNSBpSkiPKiy+XCOuMQ3DwOxBBqVD/vN4cQCqZSkwF
Do2CTO5bpHm9ZlaJFFG2n20x5t4COkZ2gONW5iGbDEExaAnckCO2Fw1l9shcGJUZ
FJrkgMvGtYWqw2sqDk9fGZPzG9xnBoZ/3QJAiTkgQD9pID1mYUsCwjk4YUBXeA6h
J9QU+UbZpuEGv5YuAMF6VyHCAey817sKI6xlUvE23TTaaYLEB0UoTg2aBAvnWh0M
rGt7GamTBfW+IAkozJoulzzomhA6JDKs7dnygYFYhJ3/Kgu/IRa2V+4kuH9v+7Es
KYG1uConpBEIFDR+Fx8s/fXf8mNUceMbh95fEYNIZI8qOeNV0sw42O7/amncsAO+
1CJtfyFDadgFkEwzjM1otE03tMGXRMiyOR9fGn9N5YTKrroHc8unHtmwrActGY95
hBVqRdI1wywseQrskMhgOVG7l/GeWvHPFwzFstgyLra7oO18mSmnBDZ3dbf/Rjt/
+T5LAboZ0d19fR113CdxCi4pSS0jFMMGCuReEVTA8aWKNDApQpqsFVArzYxcN8qw
32IKhybLg3/Tc5BR70AZ2fI+9fIENpL/4qI0uSS1SJunraCZiE2iI6gIZ+ZMbdKU
wyr0cWoaepZhryXOf1xMBjiM+4U7FlG/hCOcOEPVt/MfUzha9kZVwYxz577kZRNr
HXq0hXqn/8usKxwkGjOAue8+oFT2T3kokQ2FZs5cH4BmHVl2y/+tm/QyR4hd9m32
APljyezjZmBz6yQa7eeSnwVXsy8MCSbKXc63iFZhuxPoxhoykWcmEBePwEJEGpCy
thIoxZ4upj6mfboiA2pnmdrwxkDXDi02mKaSYqYa6JlBh1Lc/CKwccwqHVZ2U+0L
1W8XU/K5hPuTmEzbvuniRwfHSXPzFdWohVdVLkAasbmucRhPNdBfUzsqOqjnme7X
PQihQNjx5Cp4nfCwZv1YPTWMm7Q+w3Fq4d9yXlJD09Fig5W0XbyrRQVNXbwBupGA
IDHyPRvm+OsP4UywNccR2QPyhsKQtaUkyCbHZiP/3tSuFEMHqoBUL2HGVkyfR7FK
J/+aVFyr9lKN2ovCHamgCrhh1ZJL5JPR8x1DHf5Z1/zvkabBSRoLMfeFvyF9Ze0Y
eYS6li4QMxXJzJcMBgdmVLpar7Pl+wjtyvJpp27KmAY3A7210sWqdN97vop/+OxC
nQPTDfcF8Fy4Kb7vYpThserswDzdtS91Gxman1Bf01G5S7AxX2iu9h6nO9pzUvh1
2bB1rJ50/AP8rx1AH2SrnXlvDRCxIe95EOomdfPw2eyt9ghmje0tUtCD4u2HJwKL
xndjkVm1FJTEpRbmlFeNml4GGakk85HSBUY2xwU1FYa88zPpEfyIzMZLl29Z5YW7
Bbk80YVF7SSNrQF5xEG0nhLDLK66BDJ05RBtQInmcAr/JRvp8kBFmNWDi3Z1WLaL
XT8Yx7NQC73UlH2bxkxqgb1yBgRKhVTxIv5rwUjsGSe8nhtotdPexKBa+WBzsP2O
xCxh/Q6ICFMxKlyLzaRKAX9kvS6PJv48qkzYCpjmrhFxYEDUerzkq8YIF1LHAk8k
YQ95qhrrIqSLLeViydzfw+wFyYutyPS8fxbdLd61lIOl1RRECmdP5YsxsD5MJXZM
GIx56JKk/COLci7TeQfzYEDsKXKq6IDtdxNSgFAhlLBy2pXUHVb9ChTP17OgUiEe
+oMh+kTo2zo62GtD6ebBqv4clTtNQu14PHEB+jg8IqUep6KqpAmx93pg7PPZZ3bH
Uhd6CVSFetxKUjtE7VcN69C2R4th2KcNcdU+jG1ogfJ42oq2fOXFESYBZbtLUtDX
EQlmNmhNKG8NBWyfQyR8hrVlTfb0gw8KVkeV2LOALXgLLYXZB7wePrXA3bKblT7C
Qhn81F8AlvMpLmt+MUQ9IixeDvCs06KPdsncGqh9K2hy7xjyDToiwgLe7ha07zWa
TtAxDkGGGtvRXAmyK5yHl5+th1TscvdfFwaN+oZXXStEkEQsaFXKmCPi9icKjCjo
B/fI6kh09JBzLf95aSfykI2sKJXTREcFDNgfcvtV2R17QdHTXp5EsD9pYSsglqwl
0QPzDF8FD8qrf6ly2aL9nvGOJKSsG1MW1xcGzbKC+v6L/na8s1DzlRidzoe4GHwX
gWWO0ch5u63DXJTRFnUVe2v5qJDAYXu2phTOgd/3x9FUnQH+SKkjw93StNd80Bt4
tCZQpMoUG/w9kyfn0FSw6GzfjKTctgrEeRa+tNpf+PalpcASJMaSDwXWkhsRHxX3
RjTPx3iTlgqD4+MMKpq2yMZLdFL+GQobyzDKDrYkc/jArrtJ6Eq2JsLyVsjjbcVT
XfnO0mMk3WcMijiKtvvtmlfv26+p1SRcEhYfuOncj0urZa+Dc9CQ1RswJSIMhHov
7heL3GS0A0GWe5LXDjGnqSjjXr/j/q/2605HN4SB8lFuTx6Hv1rSp3UQUKF6Zk3C
MtxxzUDniktOe1hwytMqumifF89Gz1A3FA8G30N0jtZVe8mhRIoKvuACW2b7XPng
qP65eWpy76Zj7FaTj+hwg0c2qhXq+i1CUkuebkvoWUOHHVaCeX4y+ru1XIWihVYE
ab8cimcPesW5+OAamuSY/8YkpRq4IvUGgU6tD95jrFTiryg2LwLLz/0rnTAUp0Ra
uSqAV25FhRC9ExJbMBsKIiSRhxq+urVUop1z4DW97gExRwfpp854w86p8bI8+sSW
ywxf2z6QGF1RLp9L/WZMZgYuHbeU6uHs2nIHnhagsNMHGZHM1soiBB5ZBi2g+KD6
z2SnPgVTwua52M9l9YvvRgK9dxGuazt7HqJbUFiZ3NDTx4RIkR78DstvFB5Yycaw
WydrSnKI6iqfpcy/AwyKYBpEuGtcjfn3Z06+uqdk2AkI7teppzcEH8QLiGWU/W19
ZVw84i5w2IW5uDzAuuSXp5+QE78trgfH0cjr/moRZbNlvIzaXL1Oq/inwgkuYS8c
jLiiIHq7Tyh6mwAlyBOsQVdQRCmADbG1tibJigvxxfmDZRrvUgMNrP4AUpwt9P7t
g/MZEyg3Uq5Ukb1UgLoaTVufakoaDH5IeteVBfEqm8eoqcuaFChsyiynROU/wvrs
QopiYluqC7gn6MtfeaMHKlxMNU104DdNtmD3QT8A91cXlijWUSFI8R9DyjtHHW/f
4tI3/dK5NeWshIJsXYXHR/h6wskg2cLeEAAKU2MsX7qfcRUacYVoRoAeb7g3jm00
oCZ+2In+DJwYYi/5q39+BCAKLNlXrytKxAPc7l4A7UnzkVqzsKsTLZHYOKx8OvLG
PP/Jy55jsFWZknhGxND7zscRPnkdbqp4I2MGBM+fImQi4a9nllU356zbzYgqu6uE
ktsk98aVQBp3Rk3junGTJE+ilHsP6gC6xJ9iT+di6QT4/inAL8Iqi02WFVKQSAhE
ooU4hUiUO0owyy/igaCBlN0e1Q6grWN703SMXH6PYpd8cwj9moikEY2+oGUxuq0g
TE9dsjbBu+EEp+2BlIZPUVG/sz7/Qe3fBQGIsLujmzZf2rXNzl190/GIm+VYDzfn
sG2+O3PNYJSrYmYNTaXgzpfDKjJjd6pHHGvYD1Xpjvmb/jSU9l7X6Y0Hfe2YHwr3
XivGn+VyUGm2j0dyaJu84W4L3sIUTNz58s6LL2nL/7OgIVm7kemVwoTcTMjtv3wQ
Ajhe0MIcGn+3pkHP/OStj1+R0rDi58FiIF7jz5wLByk9sC6Xu0sPTfkChbJse3oi
frHfEj4f1LvTY0sIxAKfNq0t9CG3TcNerqetynXA5RYX2wJNwOLazFqovOT4RZwY
AhlNNks8sAbt5znB715y61FIE+YZDCApcfUu4eNws0RqEvnHTKLl3eebHuUJySNc
bD9yxA80zjxk6Z++Bp9+rSXXPGxk/tgFH6HaJqtl63qen6/ypPt8MDuQMnNFLVLZ
CLIYIHZV1YOeIe0e6Nu4MaBfu+MECEzhPbRwhJTMv1BqgbcAAmKzAgyMH+h+WzUS
ealB3CQCHQH8+1/AB+hT6O4lv9Bh7Yp2fEwuMzd4gp42KBu8awA+GM78YckYtnap
dD98EzPSZvphHkDd6tOUiULJa39EpchuwnGvk/xAoFCZX6nmswBwSdVDcHZP/5GI
95JSfI96gAonw2pU1zv9TMVHb2rU3PJppfxxexm1yFl2UNFG3dfI7E84JmZR97GA
Hs7FOBHT5GlXe+1H/5nctbak4TWSntPLVPKod/T29B+kQSCB446p8l9x60UFrEK8
6gytHqdwex5hCQaO3cgBXKOWWIWOEREbQWv/hsSR/HnnGmwjObeh+mkI9tj1I1SF
ZwbUhO55eg0U+HhTUhn2CDDvMu/GzALMISP1fJP7SofFC2al/O6cWLr6kQiaKtOu
uc8ehN9/wrywyD4Y9H3O5Kvppt27+gPGGhg3uaNkId8dGRk6WLGMiKFQQXQp8zVs
kCI4nFawwxpRx+wmPWvB+AmM7uH2jA3bXRlamW9egYehTiK0mIAx5AiZyua78S2Y
usDgWI6qbiMEVD/xvciYQ/KJHv9jFK+iVlS+iKS56kEKx5x6wsxaxKQG01Ycqtdy
rkJOUOV/TZAITRuOu9WyD4r6klV+4DO6joC+XTLR/1oMrJ/tWwkfMxGYKGOgUevQ
ch9GqIvS+U30YivOXuMvd8MXUUxkAh1WXqaGa6eDI8FEI90iv2bZdJF+2Xk1IAxr
HUSjvvNJkorXtUT8UdnOBcoMUJ0UX2xAV0fz5cUxUquwMl8fEst7ZNqD6yFJehvU
KAb+NBHcq1iIBfVUlZzSREv0skplZJ+m4LUk8lBTPExIimSUxYImNc/QBFKbe/po
uYDVuRbIMkrlCgTPzqk6vc0VGQzPXpGfRTzEA0veukfF/z+S3ncCXC/6lGfT6vcb
LymOmkCdTYqSYlC4SJQDJ+sEjFGIk3ofZu3dzDRwGOOsNayQHxcWqP42JHSl/65P
l12qYBQZOHl1e5ugsFeM3Cq44xD9VvBlwdUTGeFK9dv2JafATdtDsK2WUuKMPQ0G
ouxGQOhradedR+trlXz+vD3bmnHQRtdZrBx2vKbFUYXKWDOf5jycChuH7HNJ1USV
CwtObPS0dmrEIxXlbKDO0XXHA8qAOD3rKi8EZL8iFjgWfiXz0S6MpSjU6mmw3HvX
MLR9b2+yqMzaUG3vp3UeHxi8BZp68L06cOU9e0YACRoex+vCs1+RZJgialQSbIo6
Blph2L4Mh0kL7vHFosE9ocwFCaWG1pjtdV6rRd9hrudMX2nEBXQM67iQwUxSwC6o
8l9QS7KUEPjiK3rCe4Pk6k9CcBeLtAvrH9ZrNECZae6/C0waTusQusPlosOTYls3
fzHTTII8ozHTDx88RtMmcvKD9oVpb6sQCkxo4pq4pTYmURAujesD5Y+2plGfU20k
t0h21qQcoBCzp2VJGyn7VaztmF5Wu6g/ER9yk8tgR42yX418bTGgZovvHbu3nlui
FLXBzHxzqYppmwtO+foplkd6I6L/p54mOzXxImlZeW/Tjt/miN+9MTU6N7pmJm7E
L6jNOA7Y9h06/9RBMDGTRFr71KJ7mkBhEaygNeYWjFA5xbIMO/ZjGV3OJJXOIrZy
QNvB/Ao8BHM1vx1L56mM2zkRRP7aajXhdcXOe9Rld1eXIfwUb/Evd79yd9bs2ySN
icob9j6N3srUJFmac5IE1qzWCvHDM+8JhipGhQWDVIlQqN3YzyZDNYBn2LYJlyT/
8olS8A1wdl2nEF5QbMHTUCpfPhWvZmWNJmfO6DXERod1g+8Mb9efhSTwwgLlQOpb
M9BqSQPDTiT+XfJwrM27NyLRCDAQXvD0TvsbTO3dF147+/VQ3d4GheJ3kMW/k1xE
3sO/GW01jCSVXFKbwy7Ct4pJsEbbrysQiueZlT7+sjKbbK5ulyYihdQArem25qf+
uUjuoLf4+tP/iqqIFiFsS4OvK2EWMOZFL67uoGhUohcfyEyd8nEBy/IxuHZDQPhz
R7NklHmQrTbrb+ecTktGYapcDZbYrSwxLCNWDnm3riSprgEOXmcm9fLfkzuCn/oK
AzeEz5PCnZVdqI7WtaoHLssV7CPyRVrYdGQfbXJbpX5ZfKBHD9pOqW0ezkJdrn1k
+cJNmi/H9+4K8Ku4JHlU0CA6lc7+8+scwVUkqnwGvfqg8by8j//cgJP2ckemIHdO
pJYL59My6hMcbwAtKbV7Gvx8pP5VL9eg+J4wPLkDOegCGyXXNb6eFoIKxiOUYPWh
9z19a8MyiNxZEdSRZ8cugFcmhxQqbBlNn3wLdaVCIXVTxsTowxo0UjcM5fxKfPy7
yWttN5IShT/KlAojb+1bNMsV/Uhd+T6vzr+Mn2YjhIGe/gn4R5O2o2pFpUVx0VZx
Bv2IbjZ0VX9MCYkuMAg8awF5+eIHDWuHFYSc0iNFNNFuvH112wKRwOLc6ivHb41b
Yx0j2H2I+lGNB0OS0GRYNmhKRmvMuqJvYt35Qr1wqr3wnpgJna0ozpwooN8CgAXK
j1FrKwbKG0WHieYl/TfP3M7kxBYD1g2tr7fux8ZNCntu8MNddVpBHLOhn4QFyMbT
yUdhA9Mo2bRXrdI+qI5ZyOhcZTKPjED2tFu5UrIcrzLJ06pqqTbjU3/QO05MXXr/
GMrSxQsaT9C4Aw5RILGSB1ZHdFW4UWXUrx9pynuMzg9FMO5eMolYmezJ5Z4+8ee2
S8bqF/V5pC4FgUkoSJegbF3QD4v8Ht3TS7aUpIZ3gUudMKY3jH6cTwXl+566XkfI
0WxM340+PrN1uuH05ldGeerXeK8pdTa1hPlKdoakZfscbxVhahPIw2uZbASTXzom
tB+BIm+itRr6skeSRa7rooIq6YpCp07WFllTlAyK6Zfzt81i6XLZxp0zRP2Q4QXf
aVm6a7LQ/z9ROsiW7kEpTsufQhEKDtK8mMBhArR+sUjdVOOHnZsvWfU72bhGHUfp
nDX0Wd+90IwqjNmQpk3MVBf6F8fGMCzEXJTmHI0QpmtSZJ5piUyACwwsCYdT0zhb
ny2KiHQlvwxcZ/T4UrB7P8Do9An6TS24QTIdQaaMUfxiBE1P4TxlgzNM0dA2o0Tt
QqYlYHlDvPbpsq8bP8SnYQUjlQPoI7UKGe9/pgVMhcnnoGjCMBwmb3VeTw/nVqRC
5l1qS6x2/6F9y6XnndfiJIHjjTL/bmMLVmT6Q4sgLCWaCylVcG1SbM31B6V4OUCj
u3pq4JcQyrEVT1aIypq+98B6I5syr5SRg74Y7To2soEwLaP97g2F6TdECJmtgfpF
fbI3Oa0DhVXpWbCVCb4njfS0j3Uk9VEpDNkK3vKrvqFM1SMCf8JGb5OxVMTFEvwL
QbV3sL9JVQ5AHzCn2pVxHXTP7FY5nvc89iThecndgt0Sn8biDVa9jspSB571mLDw
eqAi10OroIESoK81QecV08yj5M54NCoz5s5p1OpotLMkSkSqnOFcjMcfutS5Gadb
lzVeh9nvnYEFLalArWUwWLoqWOJ5GuM2KLtwbBQvik35tkp7/hCpuu8IkCnJVneb
lPFfkDauvF1+C4yS8PRR26fbi7IxvvfPQi0sprsFt9HmQreBW82GWYPIx/LgjYxN
C1c6n+rzXTYscmwHZsvQdCZ/rN6CYLo6BcmBw2594f0ytTkFWNoQJtgwHnMsqNu3
iOwXHuvNANW+WAgxbOdwHdNDsW9PnXqOEayavEIoxQJzxtyNDgXX9V4vpp6jft+z
rCGZORgqJbDSSmuP4cDaqtv3fIFbDBsFommCHTt4LrtBQDIT7rZsZP24BtQXCYIZ
9Sxk2263+Lp1ISnWotwlT3KG8qYhMLoZbOtW+I1VMP7F7uH/WVQmfzoGP5Ely/X8
3Yk6i1eTJwKpdWU5Dd4MF/FXFXb8R3yWtreNvo+k34wSR0igptqeS8/3SHSieVcQ
Pfsx04yNuBfwZd6+0ot3pxv6lDFkQgrBOzdgRI6/42LRA1iwWh7gdLW/Uymt9Zqj
CxRn8y27Xl+nEEeg+K/W27STH7bPg5GgkeAg4X5P+S9Kfy1xbska04nC0Q74Bb2F
17p+8vSAhbSj49/kOEDI1Tzb4C+LR9Cq959+SzqaztfHlwhYejZNvtljw0OjdEUh
uC62itXlz4yNaV8cPTCi4gin94CI7Ka64kOCOmjYCwGYAlWrHBqKJM5IDdAx3gOP
GInpgMNkk2Bisi6yV5PPGT+555WcYDUYf6KFLR+AAxXYoNsvff3GocFiLWRth0CM
E49fhBgit3SPpXXb8+89oCwShGeJGj3lH5fzPs1TcJeM/Xu5HRu6vD7e9tEC/9bw
nFZq2v7BBbAhWticj7trxxzcNJYn4qZX/o1kurBKQyBCRRop/U7QcGjU/OoBRIPi
sWQLaQKYzxQySimcqdud6pPdyZ6W9tjG4fVwbRomJvjXAjOUrnoxd/bNuM3b0DAL
fg1tBnCYhYDTlK7zJYAqCLPF4+FHb9udThyp0tIfAzkgaKAMv7BeyGdE+KSLBMC8
AhdRfKyhuiaLwVEpH2ZE9vxYNHqOnxt4DPHlp8lSz2SQdS96N8snuLY/R1Ey7HtP
/N+K5EmjhKsp7muS8Z75Cqj//lXLWdXGUJT7k+SkfQuv+77HIVPoOMjcbF6/OTR1
Y4qRW5uMWWiAco9+Q4Dl2Y73ROFwVR+zjLSpaHuMlFqT+7OqJFNYLSFx9zGUYYZn
lne6C2TSmYK6GhflaNE1n3eUw90PEqczepckuGYunK9c0hbzfxW4313EO2axcDVi
O4rXvIk5teRoJKetpSJuVJUo0Nm8dGCwE4NWjIx2J1DItTLK2GQ8bhekyiCByz6V
VqDEdfWZYznPqJ4vnc2sxq5HLN4VMvkpBgN/R4XregheveJwwrsnltNn9AcW60Sb
7YmlUqmccTp14Gw1oONyUeK1aDj0xhMS5xrW2QRFlvHC806xEk93pR3KWiHXrxKp
5OQCb5nXm80O1s6W6jcAU2ekp184NMUClomH0FMcVLUeIyQng8FrY0j63e6Xq0oA
a5noaBkly89fCd0WdO40qt81a4wK8rauy8r1FDTOU6DHBtkz7E4wj9SRuFXvu0/l
wZ1o7opn5JkIVYvkd+9vnUHNRujcEBe+JykWrVM9JBJ26yyU6GAbjRd8J6bN10hV
mZmuaQH9YI3ahMTAUYx9DJTiejeFhFCs4zO8KgZZi9Ul3b9NNFIpG/OOfVtK4enU
grfHU/a9wVGoVOM7ey8zBycTnynS5RgwTlVqMlzt1K2/0H9xBis8mBppNg5oacg5
6dKTU7fEbaGCOY/Z9mY84j4FV1r4oDLyGzuvRDtiayLRC9bNK/LCQ0y2wys/6ofq
6DQaJunk2RIfTAlLpjsDgrlcO8WZDRjMUwbKFtEJaB72+hkCyhE5kP80qcxo163G
dX/rcGDf+jAPEzYqvMQNrnB39D1FYHhGtoS+z05GhoTD9QpP38rb+acg85s2Qk/N
onWczV9pvbLrX507/zyoeSm2MRmD221GEn1hlGbeUk/PKHNdQCBunsuheF61llyO
RnbwVux0RWgjOZ+GH9CkGWpgwX22waoht13RjoCNb5UTgWY9s9+tkFujpZCNVCGs
svbZQix8z6EZHcMLPdmHSPLuAEXxLwbG+zL8TEpphe8jNzaPw+GPECtqY0I0Fbfi
KXjknbpmtKRVKGonmxYOIu8JI9JjxA0Gvo7kkcHmA/6Cex3leuOeCwB4+fN9XNHY
EbUMzbgKzejWVVvqs6zXxFj2vuRGwZWrQGQ984/aSEIiO9PKXxPVkT7iz9247JIM
/37OQpgjGtw17XyrMp8kQEFAZb3r5KHL9YVD/OJwZGRy4aqA3O6rzKnOZXyLOQH4
6tsA/GRvdNkn7d0FlOH+92INVh461wqoXJlrX4c1OHHezUaAWBvy3GpY4r7T5ORt
F8Rsvvvl9sQnoCqoSqfPP6U+aYTZuSYU1lnYZ9WtV2H8J4HSoxOfAWaOB/f/JZNa
TNCcZcSpE1f7BFznNQRqgp9dPrVdlIrHAIo+Hi/diFqRQJArFDV8dZE457nYLETB
4hWiqZKj4BjldFSJUjecSaKkRJPXNXbmU6pa+EjzGDYWRLkKRVF4G8VKMThK+C2A
HzRygYJxUl1PncURPVFRT7ONmTxDm9nWcDvQy53xd47mgULIM+WMBxdHFz/BuMSe
B4JlFxleouOe/3RjhzrF5RKxEJz6BPYnvzNt/gKkljAQ0oXsVWIxUHQiYtO6riKu
swcicNUkewoBr5mx9ojjpWsECXSUsx7FswMxVOuOGc0NsoBsrsmKX4FTBVuBKkb1
HsCe96hyBfHmSTT+TRTd0njurtNA/0bI+V5hdmKNISDJ8CAX0nQO0xhxrhPg74+4
zuRT1ebFPaXvIFC1/+XGWNjYktXa+SznBbHyOwkJUdPZM4RaqS2eRak5eSc23UMl
ddUcz0G9zx2PX11M7uN4GCqXx8Ixi7Orfehp8RYs1RW6lMNrrarozdcxkRa3i7+d
IvcaV3KtbUi/TIKVIOHsiONT/banT3GR30qzMnb0qu0hPRuqWv8ky5IyDWuOvCHf
qTVcSXPeG2B5J7N4R6sG/vO+ogmbXcSeqXc3N5JWLfQEm0u6Ycy89JCMPqqxmyUa
8xdTNH63FV+A3QIAVgHzCdb5qtVi4vQ5LL33bpHeoxE4EPtpVTMPgEBlzooestc0
8ep3mzh4aL92M9S9dTCrpeN0hVR126bKYtIBujpuhHBYEwkVGDYwb9VHtCNoKpgC
lqLhM6ccFBXqKwUA55Zknh0RbkRYP1tdJ8upjhtqDPQ4oVdU835sQQ/q4lt27z0V
/n8/N27G3rmWI6pWmJQfbCijKhdwrbulrUY6AmMtZJEx+k3bfLFrSbzzkmwOZcIF
xtE+mc+dYUykAePBMaVl8DdWXBcdqC/Jmysp6nnSN9NaEohfdg3x5LJgy4F9oDzt
iTnAoFKl/jSoEEceFDb/cIyFu1/4GD2Ye9zWqMpNeFxa5JOKxcXJRqwbAO+rYAGA
83r+Us77MW9IkmN3wIAEWYU6Esw0kJ2Hisrcs99gLpTYOI2Tcnr7B0d0GfVRGjXN
i9z6/0YGAPorwEXjTUqhXHhK4tuP0Z3jr/wUG/SSCmNOvrxXIIf/7G/R61H6TAMs
eu55buIgTaor9+V8i+0CJeY1WPhu8BuvkF8FUNEW8K+zVe+bQWAvK42JqQO1d43U
UbEJXyWVhYY7fleQfRBKuQ8QkNoBeUXLmPdZrOCT5byJezgspj7WLHLRJ5vuwiOB
AK9Y/wo79qPu7mPeeFEXjgWW0Sy6aNaXp2Xqal/2p8OktbyIrwNb+U27NdFhagCL
/KSL42OX7l3Uy3tFxYCUtrfwkCW2sCbfT/jQthtHZaV7jhsXsOX1MNJsrwtB2JoY
b/phWy6U+Hl8W8MH/xieOu+4sI0+NnnnS0LnTrMnj0jH6IceyC6iqfZh3f568PkI
WLHcGqV8QmYnvmcHhjk2AG4wpl2HtuGV1VI86piuj6KgFTl6aUIRmbfjZdfJZTBD
Mnz/l05L/MWE2U0ZvVx1Igl6mwUe436wkOp+NqBJdpNpJg3m6TcyhT3sYI7KDdor
u0nF+IYQWvte/FTzeBT+uVUiozwSOvlOwk7chweBXiNE3uDYYUwwHF5V3JQKEL9C
Mx9hccdLrdZl2ZhiKVG+ahHqtPIZI5NSZ0MzTnrYO919kY/xxJnMXQMZrzV3MO++
Y7nvG8C/gxxNYC2Qqd2Wk47uZij6+hvJAsTZ4j8+DqiOnBETK+Z6PlaHs3SC55M2
MG0Ya6gexas1FLgDkFsD2VGvc/6Z/YNf2sa1bCq1WYPBQhf8qY3wRqZRsjGdcW1F
p1s2CRAelk/15xI/fR1TtbDvMxI+vP6cFX/v0tc5c+Wgc9KLGYJyVV0fxnXArTSR
ChcVJjttnU6kZFtBjqm4NoDYbNJAmxerfu70/zCPfXymruWWftLda2zeppm2BL9q
HFohGbjHxU9NszVBCjVVVaUXWdrU6lWiPjBYCV/uaYGjf4IkW0+E5R3ebKW0kBig
SbkaesWJxluJzpRLP8CtBJ2WAFThzUuXQ8BeS/A+TYjfL2l5t2VvuNKGT2q1EoWf
t69cLb9pLJoHnMEEWTesfT+4rTZKiw1ScymGdAulnbsoayYu/xvX6gvKiO4+8KTO
3Fs/axl3czNqdtzQfOmCzginEZ1tYU07b1PzVYeUk7wvlzuf1AWDDC+TwYNK+V5h
h27RdTrZmcYDiQw9lCYOjDTS4RJMxdsmY+neAxsN/xYvazq6QOLX+MXZA5mIf/rm
6N6fNAS9H5QcozADhbIa7uRENQglp2HXJxHaysxld9iSUiHwXX6JoLJNMFxZA7Kf
ST0+6/rkbXUjF2oAClgJ25xqmN5ijIMOfPAQqYp7q6Hnu6Vgiqz3jyq1Z8bavIX9
YGMim61YL0VyAT47A7eymeE3pj6H8GBJleLqtZ3V2olrLL0vdRESa8p6UDy38oJP
s8EAXXHXXVtMdnW0CoRzOflf3JqVQajTQwxDEEzVmbSjY1CD44Ehwn/VjxK7C2Lb
OVSvmv/Fl2QbMdArVExxYD6SqLEiHV5vY/POC2g5xGukby+wJxMaHHfmqsUa24hk
w15h/QAJD6OMtzeTG2A63Fk8RKpHOR/TIlaYRLRf1tc6extNwnc1nZ6GCGgMbKgZ
qmslNPqW9CVyj6U2+TZ6zzhwMmZSTo10IZYyKpk9v5cMmKACtzCW7VdHbu1VtucJ
Ss1/nM00/MHrP6msmZK0Up6iVpVowtVg0ZpErgCYGNQlA+RtVy1F0CcFqozOSItO
j9xLVI/9NvqjGbWA7godcwwefG0JiDB3Os2WKau4UyQ4KlvE5dGQztYRzg53Tv2w
ZSzgTLhtKdZISyUEXYptGSH+Qm/sPzuwRaqewchX9wcxAzvmjifLfPd6Re/M/dJe
FmAXszDaxK1iwbAs6S8cAdYc7QlHWE90m2B2MjLtF6ZE05fsCzF9HtE6/1DpD/TW
mZJs8BrRGF6/oXAWUmC+Ib7ZykaOofsYhdw4ROjuJrj2nWAZy+d/JYTc3pMBLZC6
NtLpKsofkiUwPgtzjy4CGwpnjYORCO/O0TpOJ/21K/zQ9XOR96k3vHL2jEIoGY5A
a73/euGNsxqW0hm1M5wLxVRn1dqmZeJcvnKhrfiWYZodkzgjFR/n5z2A0uw9DD8C
Ps83C9DNGdaahhuHNNGooAh0YqAYcUY35+oc3yUO3hP0dpujZt9DZm0GksnMr3Pz
Xkw0moialbBhVSyOSlLka6iUnfakGqVp1QHRl2Nr0BJUSHFNkadFHdaGjZTWTA7K
wHS76GDj2G4ksH61DxiLCpr/rY1c8Tot03mVrKkgfGcgCTEA9CL2lvOJbJ9voLxz
pHkAj+5pjV/Jr/9UARH1KRFJl4y/v7Y2nTV82DlRNpF5E8NrfamaBE3lGAh+PklS
Tp+JcwTR4vsTwKb4xUeZyEnT+6J+Ij0Ht2AXMiTEwJsIWxzf86s6qGEgnpt/PNqg
VwdfgMYcVMYa0Un+OTe8tUvt3hiSVo6MwetyEW3cepeqOWE0tY6FGlIB/80zph4s
F89zb2IYTCbRwmYmpff+mlIwbJXdwNeK3NmVbthnRz8khz1tqS0LUYu/W0SH+jZN
/QhVTnVcbscOGCbo6TWPNIlroFhhM+RsFKdvDvcAqJndPaeJYcHCZlPI7t/MU2Oa
Wn1cAONs0lthn6rS40ZN5o8a4/lgMeZ/D13vBo0BWaxAwNSg6nzhhDhLODfxRepj
ONZpTviFjrBQ/VLbYdHms4IV0zUE6ri7qH+nntgKAS3zFfoVXGmOFgrdu4dTA7vg
8J/3T3HEsyEFtqq0bk9WQma/Tf1uOOskpOvLUyOJUybcYYltKY3ZA0WwZAnQjabf
baxKYpABiOI1rm1EfqYYhuqTXSW88wtB5JmL/OrwSsLyXlbLjJNpwhBLwBN3eztL
wUuJIvyYg8WSqn7e7Kv9KJslFfnm/u2hCYUFSaQzeOMiFJV8R6rzjYihNIVW3ZE5
DxAchvcXwN2dD1YoF2juHdakIIkl7qX1PUKvroip48SiVwVYOfd/XjAihbdTReSy
3Uc63VNRjR6ZDQ8z8VuO2zEycNjJT2DcyDHqAZCZD6Nm5wRO2usjtwEH1uadJG5i
ujvHr/NoSyzQZpUX6ZZrOKEgy7r4OiO/hO9UDqb32RVqdt0ceaP/NaQkaj6VvW7G
YwR46YKunKrU6wo4EJPhRr6FHOucZjiy9pnjxYvCWgVXrhqZVNAbYrVnB9lNatpb
fWV5RLMveOGK9wNlVgVsJM3yycWIw9pIvWhjRZsZqC71WkT4RvJsXh/g/h3rPhn8
r5RUVMzBaUU4G+x1tPWTiTBiw52F97q2dtTRpwfFWYYYlcj3rwsFo4DGGZPSVpTr
V35UpYFVuxjgABBuZeXAIJOIIzf9IAuNLjO90g+Q5dwZD9GMFpa2rYLrFBphexCn
0bEztkxsvJ8njLr2nw4d/QNnw6Cz37k/5wjIPKdOGgqavoukQjaK0bAt/+Y0G5PE
nX/SjSddSJVieJVhgmeJy64juE+8cDK8z9JQzc66VpMn5qiv6gPdH9579vLkZ7K3
vWYtGBVCCtchrp/4K5/k/+iTozMy6+ArNTtioQ1Ysfgjg+TBmDmN7Sn8koJLGDzK
nsWiNyXtMgs36ov3gzDGnpF6jlqYmS0cIZM3Zaqxxzw8UcnqFn454grp/C22374K
Yk/G+CHMpmWSiEN66p5qm2nJs5+nBJ7ArZljouV0rgAcg4A0JIb0eYH/VUsDpASd
2ghIbYvsGlr2jbT9RfxoQUjfdHrlU+fB69mdDvwGBhhBT7HCUjr+l75xYE7IQMtq
aivK+xv060umrAUr+aAn2PDQpJbXHuk9pWZb2J6+lM2pPt0wJxZ6ZNTZU6PXrXVS
y1yIUk/gOV8YkabkJmJTePXzvJMSK4m4vBGjjvHOMkA1EvnRjJO3Tf9/gA2TMHJT
h8ixI9vAdBFv1lVccuUs/qIPrUdQfbPQahOCWKz9PkUgft0h20FAOkiY8zv38J/6
fw+K7utR9znD7IlnZGXqKlrp36nBCcxgwRFf0ShGMErDsm2DE9x3jmWHGG002LTl
+K7SxQFCCUZCc/VPeG3Vdw2c7CA+CqJQ7Xn1J0nFhIDV1KmJsIg5ynBCBc/6oc8y
jkGkwUrjHnoTAfnkkz/21OZXO4AN0x+/XjTpvuJDCB5K+emHbr4SzSFH/ouPV0uO
fOHgqs3XlwvkFdFRqlyYwX3ixuPsG/UNZcZ2O7Pnc4YhcEcjEGQMBn69I2nt314g
n4yEWsMVHoriY+a4SA1LFd1bJbK3ZcncImiC/fEpQ8P7jnSJfqe15aDy2AOk2+Yj
O/uxSxcrA1BiXe5oS8Z1XgO27oI5VO9NE9kJ649RdRkQKkH9aUudD2amHFd3jogJ
OkajqbL9qns/whh4/4SKGz+vi4KuVocKn5ZVcCzqt8nTO6ewqGcR60926cWLBct5
iGWoSjBcEjyox1fkut9N/f3w5fACvy8bdm3xBoX83ZX9pgvhn3SDgxlTo3wzk8yh
3yK7vP8AyxxYaxaFMc34UPurMXTmFlB6Ol/X8TG8C4A/jyrytZU/tpM4d0nACUtr
yKVbIPb8y14bDY+iri06pCb0Rdz71HKmg8YUhe9n3Bm1PC0QRUZcfgVXyWl0yrFt
+cjl678O99AtLF2GqTT8FcnJgx1XydDi4vZVnw8J24j6T8W1tSyC3oZVXQHl1/Aa
Ld+pDCoVncesuKpkcZEGv/F6j26EJ8HHE7fMehNaQKAIZpwQ6FP1sGKA9iOqGHRL
jMmb0Z5wccWon2KpcqjWTBZSYexEHix8sbtH7JAJ84dsjY2GehuVvfK9aMB7POui
QM2gd8CQX4jGK53sf9OZ4Tryd15U89E73FEMTDmZkRoXczL0vptqrl1GmLwWzxOs
eJl5/X7oFhXcPMRvwZdil14vqA795l1B5IVI9yXYI/JQMBc654LEmbfINv+EXgD2
3HAW83g5p91ebZHuXoM1pTGgT+6t/wpUqk6NZBrDV9L8KSn2vtJYKAiaUzZyVrk8
valVnMoo5g5GB/vfqn65QUCIyWZbMYK0hqUhMGaarVR0gff0fDmSGptplQteB8DD
oNsl9JM3pz/z8qAtH7OIIk8nPwBj4BEfm+jJvP4d1ghcyC78P1W3l5PoHDiuIC9p
OMQXzfB99+F3hSD5kCmWvSCTGoclRj1AH0ofBYxLyBgvq4FAcH7y93+5qK+/5jFn
C+wrl0LoXAO41XBoM66AYeNpdeImf00EsVqoCOyxphoABZy6Be6qM9yfBsftTLl3
QwAOiuSaQyUwdxlZOBDdlM/ju2p80+Lv/qeQ+fj2XfR8IfEUJrHzxsNp2KjkAPaP
wzy30PZJNqpHlizD1iA4xDrfUbeTI2/x/5ZdSSSwyFyG/Qv/vuP9PM0YiQgPgQTE
ExGOZuBVm5iWDGL5/hY4++ZYejHTzyB+7IVI1xVSySQ6j5Tu1ofN+LKkaITF1w1B
O3RrvCJ6PryOuVMtU+bVskD1NcrhonkxgutFwO8Qy+XAngxZtFg/7I6R1y3iArNu
bRz9T6+aoox7Dhk7bZtzJv30joKsF7pe2tgbnqk+I+mJhDkpbz+eOicT03ITsEmC
WNF/SfnBZAJdJZLoGMTRE8Pjp+lyBeN6CAtyzjMgZWzDoo03HNo4/Dle4ZM8Vj04
q/RxkvgRCM6cAYVc3lxVZOzrkevdkd3vXqYPPX5P4fGpI/MqX/vWiuysmsKiF8wf
8nOG7ZHX2if88Av/Z1F/N0aLIFSmmuu18wCDqbIkWor/AMuuoAdU3HkdeGqN6hse
PqTfKaVQeCIgfAjdsWRwjokAkUgnUSIbswWKgPEnNkTZCXVNhLXg9TdhWIEky9ms
x0YcN1KJOQlR5LNGSdiDLFvctp3nOXHozCRLcf6HhQIBYIb3vnk3Lw+X3zW2p/2b
xOj/FSH+BPtY9KjymoJ1AMUVrrsPAXkR05R3RZYkMFIKfTuqBPK5OmW4R7Rx1Egg
T9P+mLmKjzj4jrmA4P5mRAKGt7+q2EKadd283ZRTnJm0qlnl0260UABK4h3VpV10
Mxb7HNCo8n6WBFS9jCRDI2m8n66iUZyLvAbPstAC9oT4u6cG5W+elWeidXuS39x0
0n5hWh6r/UZrb+y6GSZJS1Xy0cwGyqs00Lwj+TQgE/Y75/zfye6mmOOf3yItUn83
Cv1/wMOe5Wq4Iwjbd7rWqHTFyRXBWWHtE9zhyOTu2SplDFRqZJy0/l7t3FsntRxm
SJRw+c7lATZ93AOS10kEqY7rOyLOE1evxTElJlkAG03yS126bXv0XtWR1lkE7Kmg
aLdYqstEjP/2KJV3QcRMC9VfK070iWOi3NKaFilztn42kgP+ygU7eVzGf5/OLyGy
bEY8O5K/andcbKjzPNaENCyQWklCWAjtiwfeFki13mt6HEvd8mBcIzP1q+4+iFYH
k8EJ0gW0LPsAQumXJMIODpq9BkA9dliX1QqSYw4Pk82la2/Ss1zcnxBJP5AF+dyA
xpXycCRO9qzLA2QnhjbsmPQD0sWnVX43Aqrab2OW1x5FVpQlTCRQV5iqEFK4oqnD
+s21xVAYOAtvDIthNwdchSucC3Dloi8uWhxZbuaZksJbUjlHxJuj0f05l0xFZ618
zSDVNTx+ctHhqwRsPR0Wzw3kQw1J6lzmzjzuBOC5Gd3fxCpJubKTVBaSugw9bAKy
D9WeATpbsk4W/kxELPapSbnLqZEd2oGKU+by82tgTI7BgNxFCjrPifDgTshoKupT
/FZHipXCjaoSUG8QBK/zsVXWLuhcIZXx+1ktMjp09E/Abw4eJ2h5p/BvL4IvQtoh
MjJzcZhCiMpd5TQT4FxqyVOQSr2U/KCYZZ/NW7F6ecS04tYvHwqVCVsBTly/XxD2
HxQjAvmA/K8SxPIm3JeKUssasN28YvG95wvYHCeago+pcMFGg6ADZReqbuB2VarF
SaXfUWb7gFlfGPj2lYHJf2SJxvhE/a/RE1+hkA9azDtUrYPW6fsWh/A6/RMZZXRx
73HEe5Z//npxUl4HyPCedgSxOdHipkNVPEqMTKSWGbq8fc33DGa6OD6YtONnChbc
aPjtL0uEL3GVszsT55z/Ae9m5yHT2DxkZ7p77lXfuH/hvmX0eKIK8CFknWMRtyKT
o2ozA154ulKlwzs/a7lWSaxunZqNJRub+OPCzT/cqzg7L1ysJW9amEZIAgJ9zx/y
4KbG/KYsGRADuNjTHOfm/I9wQ9G2W8TlaGLyCsw4c3TBOFAKFe0LK/hWthUKPTWa
+NZME5Xf0hFv3qH2DNG80j/cNGQXSwHjQZFoPp0JuzrfjqWfCnSHXr0lDZW7Gg+5
9ngCSPZmsVGH1dpB6xoHSHmUoCnMdxv79NC2/0T8L090dfsye83XQDjzutv7i/Zb
irc49/0hkr33Xe0XcYCcqkyDW213FERlH9CWpVZ40Oe7ICxoLwwjtrt5fNNI5e4X
gjv6aIZpBM8MNAWJcetyqNchI2a53qKWil4qW1VBXsg1qMN/ZxwL9vgGQQww2IUV
OsyOXDBLGsIOcRxm9YqcxahozD/2rHyq2eCMNPpIbgDRGJhpR+JCgTwS8i6eAMds
inZNWAzDCROS3MPk7Y8946HXGQ9rgmf1n1cUsXTl3w1UqeKLY6vFoQMukCXUAKYc
4zWKqPNP1/+oyJRfrBrNbsic7DMb957jpiap7q5LZanHkV+y+EKQ1yCxRq1thR5a
wtwaZFuWAEKDjKE+d/1+crsRi0i6oRb86R1DXTlabXhqyE9pdSZMz3ZNDfkRKube
Rg0Etur9eCmlbl1uBWpmbfTzRbIPhzsrzn3rXmVKeXV0vOew96j3mus7Flh880O2
zP7MGcoC2llwAJNqVRW/R8g3EciGUPcT0g1LPwrMo1hbjiJ53ZWCvV+TVsOjsPVO
ZYYiDA0neIxt/W1bNEbcqbgz4FTbIKXZApUtI1QiEmGmN/kWTu2yE+ZCZpESIzz5
3xTmWKvJWf1Qg4U8pMFigGPnB4G2T5szou7B8Z13guXbVx5mon7NpxpWGtGXCDh8
e5OcT2RAnG+I6gssBsPRrv17fVFIO64IOlNyE2TikhRDeWIWqZ0kCVAa0Dmj+3Yk
Klx2tU1bxpNsWZ+7JWrw4OvV3PbX8S2SputfUQ5LL5bAfDOKarZ1uS7pIWh0oA+G
Bm9+/PwOfxoaH0/+SFXNz9wwHXqkp+i/iJSndj95rHh1CHfBp9+JcQmDZvxJKNZR
eTv2WGNWlWI1Ulw7Afkvm1OZuljtUnABZdj4O+YJFqZUk6tNOySynZMOGVqCC86n
dAwfHaWvwpBiV+N6OYEkiAQYNS//MI/WKnMg10EYVRIXTX1F4f9DqSCnLcKoP8TH
lZ3txHjZjaIHzF/ZjhZ7zrlh2WznbKE7j1pmajkiWfheZhG5I6HNbCWTAMUF5gNQ
BrtNJdRDwwqahJIxX4cCm4nhsziNzrcYwnx7tE7uRtndrFZ3X3ExCnbYR8Ruf5yY
YWM9zXfMsXgaGcexPI/3vJOU7YVRFf9uaDOLlxBrgGI+CY6MKWGS/CBt8lrYjTW0
m/4au5U3pfeubDrQ2GbKFD7vDmmtrxjUvv3uC6iw/rpXA67qn++LoPVE+M4z8s6L
QT145Sb3YOhWpZSlVJj++9XvFv+DLExfYPkfHmFNe8S4zqVfx5l2rRXoayFCcB7a
6s/Gxk64c7tmK7jeMnymD8EG22DzeVcT5qUHE69owG5VA3wSOWthR3nWtd5c4mdt
Gn07lGjFdGAwEfDE1t7JlMOMQNCNl89+eTQCU0Fa0oYq6YxQ+wkV39niBe0hkCFO
shDJpe/b5IkDngH56TFjzNHMyqhStI3xdWggSxfPe/bMPylpg3aHiUlsTeX+ee11
ssJUkn2hfgGdXBRKzadoADVY4CqSgZhTkNupBgoXpmnPKxML9Jl70sLQ3vCppinU
De8R8C59U+IOgqjS7K/smrQz2AhJyBq2YWeem3No8gXJOPdF+krXCoBsxmoJvqCt
tI0+46DHed/uRZYcKOAlKxptOealkTlJJnzoHFyvsA2B8UUEn3ksjQGSdWzJTo0U
ODbMWbMdbNcc9K3nFedpvB2Pk4AW3V1HfTJPP5yyQmvjNtl72K0dMJiZt0H+s/zl
ol5wf6qCuIVqvTq3RtSAKhoEsvqRdnb9n2OYO7A3qynwI3oUbOa4coWZRZapZ52L
N3wF1B8Cka0aAjf1b9RJ6P5Q4HKeyjiUEEA1v+WQ5L7n7zREjV4FyzW0us14Ns4P
BDKtPjxnsXAHE+QyHWMdMyLjVD740NNwlRMloZ7ijE5v4efNaI6wrd9LPd/8xbBB
1EgCjlh8YJ5lilJyThHFt+bbzYCA4kWkHR5bmkeTVjHFAVX0ZbHIjcFvPivEYwW9
EHnqqhCjEdg2t50PT+KdQs2IGewDKlq3vSiDimZE3sSzZp3U1gV3F5xzSpKR78iQ
yqIIJfGPCPXnPTj2ug7Ns6/oEx/4qUw7Z5daBwWjkzPpAI7yHdMxOMVkVvA3uymt
/xwbxv9tcElVUgkCP3f44IkVGwq4JtBpf8h9TaS92sIMsXo6oEmnwwyNIi0MZA5I
fMmRF/VlCKJ+UCfF8J1ouIjsT1/cAWPrHAHfZabbjeDZlgPbmZNH4zZB/xnriefp
Bn7qD1XMxlFKDYh+Cvgw2SxQVL8uSBqiRYrl5Rq5KWx4rvHgCxoJZR+UzbreNY9M
UEmRS1CrKzY771HuHDx0u95oq95KO1C3KuPthTpLbD4aDEt2tUiGWQ0Pt/wia3Kq
VCLUo/n9jPS8VgVOA3kjxe/sC7tXx2SJdU/bPhFJXd8FCwyVTzcUGy2IeK3beXje
NpQUJUlavpkh6Y+GB8JNlcfMcO0C8pDD15XnNCnRUmuuTPsGHlSb2aAeMOJ+vKHX
DGQApz9UU/qjFZt61MVQzEMw5f5EKN6EPjFS0MhZ2Fv2duphuxuibfi+I9nQi3Gh
uQp/CtHHoChiwVvS8D49BOU8AH+gZKCdnLh8MLJTZTka7t9IP7pxodrfagkhmQD7
zX9nF9W7qWxlF6sGgjuaByv7p4UVf6m5QVwN2fS0kKl50xV0mWn8r7pygSCzu7vr
vBWxxTIruFtVjQSUgPaN6KdhtGtZezLAIdpjGD9SAFNNW3GlaAWkxQCH2hcgA0/3
oWJT7HK7q6jOvzIs46d+gYmIN+W35XZfv+CD9M8fwk2VWVm7BIysaGp1ry/D4oXp
GFDXDxsKJ5mPR6csjvo0sg/shNs4HPVSOy1u8lBKuWla0Pab0U6yMqF9jXM5XPN0
CakZQTSqMe1omViM6v5zqUlk6pOdMQq7l5T26gyb8XGEo3GuvozMF2HPwOp7tPbq
EvdsVlI5LOTivsgQ5LkYzeDMkG9E7Jmecy5hEFQa3MLqWmR++DPrH3gLJ8FmtA++
PL4ZgTC6jk6hf7iy+VyB1SEVJxU/6PXLB5zoxkaXOlEpE+Mi6Ja9a5zN/SgDgSQs
L0UgQWzBBPCP/DGy6xM/vpoETHuiaFtgD2GUYONDT616ZTvU/5/ZiNLUXPcX5lDU
Xux96FEov5tCLrwkSkFOWQdWhSPayqi/12mrTtnGpAGm4mbmsfaZE3PLFWnXQpIU
qi1uLuTFFKp5eLZtyHA7XrH3Ogy1acl83TeHH39wOpz5j2tthmRzYdSntp9nRQr1
H1HrADF+OxRoN0OWqV3VpDAQJldkBqmYo6coF4qRsmb2l1D/b+3057jOVhoKjdJ7
TtelsXpRIGTrZUEO0NoRWX6dZheypwFV53KMPsaJgtkeY2XE8apwTcLwQWPmIo7J
dao1DesPx1BoONmVuPhG871opWUx2RbSLR3nYHXH0sCLa4+nzQEI+ixbTSAnfw+w
Ow3IWxXb+yNJY7LVD0n4c2t9F024GNBzGp+a5906irki/DvJZGNEE9EAxOLnheHM
cGECSuOfoP2m4yDiL+OSkY+qdoCY33grLtvQdUX/S7mGTvVzhPkSeMcQpQPCI1QY
HRGBwqTEkoSBkEqPkqJbdEU+RAPh9wlicndZ6GZqQQF/L2uKS8tQSAyGpx+VEl2G
2kW1MZbIN0D0yslcs3MXm89d/Oy1RVNCGapT9eFL3mlVN1Dp0lGopO+ghw1WrY+H
zGMOyxWSwXmyjs/4DGFoZqGwSTqogN9BhO+NVrNITXmte18GcGrYst+A5ezdTuqw
xWd06WXJAEfv8FH1uMm2xAjumaxRqJNqHcEnzZRkMsJVwIFfSU82h1yLfyRB4pRS
nf2CpSv5QDnq0jg1eOw5xRg8gpD+oB1Nr2+7Lkx96+Oa/w81IGtgKstyVDTNxIQg
53FPLP8oYVZbC2xb7uFKeMMkW2U86RB/w0JVA3ZdONlpoBwQEfcxvqk06VSmsOHz
kZgMarPt2s2oR41inoqs8dwUGuNhrbCCLP4c3dimeLuL/1+kwfmJ3Prb5lRUw6kh
XkfhOVSOoz6s9HHUiEEQ5Kqov5DbY1B0UDiAUIvHgV4wmeIDG8pV65D4qyHEeoeX
Rzs+gfSERo8AhNSvgQxK6PBzuQTu6blj8fyFulAhNbxgCaCOppJGkhCjiqpY0T8G
Nf/zD+E5WdoDbR/AoyAO5FKrc2SPKlBHfQqtFB1JYLEcvSy7ugA+q3P5I6gijOEn
BoyT1NHbREVue7WvmNMeVlVhGK+OjLw+sc78kFCWGGULWbsFxzTG8uLtt/c/jANG
3g+7zRqrw0blSSgZ3SLWoraPcagP5eiLZWmRR3aHkQjAHKYc8AstoD5DoLszhkfd
dxZiFP1lTTAC9K/vjzXLvnLaiSkIOAcnTuIIggc+8t2z5HhNRv8/PxZZQsSpdsVB
eHlMR3M/icL63m2kHC0zaSpU9/aK5zLDbDE24DP4RCP/JpBqHCLLSDmmhN1O5xpV
QFrV//6d1rf8285XxJeuSD4/rx4Ks4VNJNk69s1MfydgOuj35orfH2H4wcAW/R1M
/3Olxt+ScVdpgJj6GBOjtXMg2qa7z3NgDKmHP/LhMbEwgmtU5fW78lMiTbKBF9HQ
4UqzW4OB5QEdIl96+cZfRCtob94JtQdp6mPQwiL4zvvRbLSV0WBotFjOe4XvhAYy
6H9lp5QOSTQVstcwKRXFqkY4oMQFNsSiUxTgqYV3xZK2qPQM8aKC4tJU07ilk1QC
8ZqbapcRZ0TqIHygBxeNPgpw34DttFri+lMLixBlHM0nSaIGymreFkkfz4YZVxcm
QBDQCz/CXh2vfrtBDeSWECrL7Z6M7LsFAWQTSGEU/733ByZe32Q21WD+ZoqRbbyq
HyU5IKHZ3axy0CGueHDO4m+2dlQAue3ot3Pu3AjQpVW3FbNtBcS7BwxULjyxFdDF
8HUI3Cf4HeP9Al6z6YubGfagkQqI3eR3Hejo+lzHwHVNm6B5WeBI/Lth8/1WafqX
rG6WD+kxHEqXPKgUReADmLHQJe51O++E2BusGgpnsAnjsSutmex7bjKCJeO2A6Gf
kLinMMy2EvldKgNJ+C6M1q0XZV/AgRJ9S4r3c/nmcrVYG5csEDGjFlZ+X4N2Y2YO
NjUw6M1TIcnxAEhosUQj+uEF2yHBHpxRMhdUHo6sDyuXE4kTLTS7Ne67Iu8/tb49
YR0t0Lgv9BQtw6MIeMNse9oYtG1f/lyy9d/ExK69jUvlZqqdC+llN+oWU2eEIlAt
xJn6DG/u4z1zqFxkhLDrf2BuBI42EbTzOBBnABjAwwKzB09tJlp7eTOmR2TdNwA2
NsdiPiJGXduWheADrSOBJ/PZZOVxh2MiB+aIoA0Xyy6E3m/WSEi4qfl2MsymWfJV
U35y35oPoM4TghQQ+HYACh0q5woSYUJUv8f+ROCrbF+TCXlr3w3Brq/B26dE4IMM
KLA0/rF3+MPc6HSBbeAOt5HG1nSAMR8FZ9l/rj6SpJx7FoWZYZSj9nhKcrrt4bIP
spzSBXAGWjW4lFy2eq+aTGhF8wJ6JI5+dn0Ea5Zbeov4wzsic88Qb1WMJSW9uQz+
oWKlZDdrtPfJOpgWaPzTSC9ZEkCuxxws82njG2UNVxhFLOQE6A1YH6BOHwwT2VfU
9gVVX6wn6b04X2wq+YkYcVgk2R8tPDlwNs9ywgT0VKVUXqeWMZ0EuRdFQ65vKR3t
95G/+nbufMr8UaIjzUq8eq/EvP0VbuwzkMI448fAuI57btqCcUKWS5kSl5tkp8KM
aiHFQFlVKvdb8AqkeWw/w/5capvlCU30nXzjTGUxi21aGlcw/jjkFN3V5joOswXi
eDdeUD5XwALC5G9u3c6glYRh3j+O0v3cHB7cYOvWywzCmNfcVwxfPEBk62ylYDuZ
bRgUidgi/WYzL7c3vzNh+Id9NmYZ79PBKRS07kLu2PBIP47r22gg9CxXLgYTgLpr
jABvHRCDqVqhzDzg1T/Ru/ivCQCeTBscNoCqBfUYwO4CMju3BO5QxpECeXLD380/
Ch49R381x6RqAKpk4nnsUjtSNeSoXhkfLDZRI4CxBh67ZBvNCIEC8KH0J333VBOx
UuuJuh7JTMe7XQpCOYmgL12l7dojSxYj4zZRJFH1cqpFto1hT3wRFcFwTHD1xl/8
KYcrXcFbcK/zj13rGjeNGmeST/GywzgX+BbKhvrIbg8LxqCnTf1zmlnC17mP43Af
0CC9b9mhGHINcuOS5Flcs1ISlurwF+d84RB8R7rrRsEEtRdbRmrEMfVnCY8nz/J7
PeDHkFdpXF3L8LkK4zxjJeR2VAdzgNYzjNUl+o7ZrlTSyQ3B9t959R7EA8+WxZHE
GrITjJ1ZSyX1lpafw/6SQn45Px8Qx8IA2eT9Eb8ZVfUFq7ujekzXW2EB7h5kh/nG
mDKYucSng6+Vf2GVTy1puV4wa2a8QoBVaBy3+LCXf1DR3CwNDd9hdHo0e2lzVpPP
Te2vr0iFbFw1dUfYEngC34NYtlyDd+9+M3Gd2x5WKzPz9etKY/aJG3hXXFx8THZv
/qKqRGiHq7FltY6ON5n8vBCBfu7/1N19ajZTcpaBCuqXM7qbsYMbRK7kuaQTCOcB
XiWt4fnJkGGNf10NjiyJc3Z3InjiFht7HduOk9RisJBzBcLfkzE+vLl0iG1QmDVk
3UbSGPj+pR18RkFKdU5M6rY16nreBiGcsWFEghtT6DLAvb2qs5um3F7SuTYStAeA
pGm8poYRRMJFGcEd+Wd8mXr6tJ4oK/mIcuGUEqM29jaO2QWB/LaaJUEeoRx9LeFO
giGj9jmiwbIbDjyg4dFp4Or1HUfXRdvrLLZhf8YuqN2I1KJBO2s8hNsUe7IO2Ynl
n+nnTPw7saE4lijXLX78OGJTdry4P458Y/EMr7iInfmGPtDi0XrxWSKcPTibm10a
nGuBNAT/w9bnvnSEQTjOU0FgkzSXxdMwmNvhVx6PShyZOKZp6m7FaohoUjfCBK1Z
2XkRIfaedQKt3qf7qqv3yRlChKLaqISQpRwIIlS8CRzbwiG7z9m+0YV816DGOStd
Map9fjGLzSiPtneaDBtsoF/5R0tL+UJu4DcP2iV8UnasTWxIgdUyMS7Uy+GUONi1
MZdfpt1CDFjahbNZSlnhV6aV1bJd5e/aT49B57h0srl70VLZKSDHgI1IIxhOk3BD
e9i6mBih0Z/mLbFhD3q9ehwGDGU3VgXHTeoJMvhYBhXYKAd90qbnrurR6MFnvxb9
EqOXV2JMQzLbMujozPESuQHHrsfbZVoaIVf+dCMTzftQALMnVuCxAZMNMPqThLbM
NYSNJD4EmetjZ68Wvy/DF1uGxrDBVsyxiaw9ovs7CgzQimU10UkPWULYQ5suZjiQ
qJ871AhjJyoHDJV62Xv+vwTOtmV+hbw4Od9t0ieqtlqd8z0pncAXi+7t9xfZSqVV
0dvtKm4f2ricf/vn1TZCrhCHGqWj+8lN6EfUWnkZ7nfI1X3mh9NgZv1EqkDrAdqR
Jvs2LaxCpCkk/xvyw+O9U70hFvWxNqsac/02BrFhKSj6dlfa1116uUhf1RSqIXbc
Bi8eJEqQrcOi1irLhhZ8JZtuFclWV26c+S3kjD37FCTHSghw9GbfcUfPFzHwzlMS
nKXRs4x7EDchGn8mSuLHoRlB+MnhqYq0k/CY6a93PdWvSmMB8RXTlBZknEyryTvE
Xj8RV1KNIeSWiH6u0LjxevMCAW98tl++yGp59fNid/JrJkzqcidSfmP64aON1r7d
c/ejdgrRGdhXdGyvS/doRxeQlXJM2BNUYDymlh4P+wnVxNQhONQl4NOVI7foJJCd
HghJzvlFpvDRQY09bh+7lGaYmsJoDiVv5s2LmSkE7NOD8GUl/k+/tMMqrarxFv6j
znBZNojsfjSn3Nwuu3L4omfegERMQgQN8EiMUbGhDm1Ho3EWsY0DPXte57V6rziv
9Bp7d2oAENhDEIYivEgIB6g68MdSryOGgcTLmQX/JhzD8L8cpq8brFb2/Y4NzRW5
Oz7Sgr0UoA1rovC0pAMMXzhnL/e2IpEOllD6VjzVlKyqgpqvzWp7YduIbCo8tvy9
uselZXmuVRAuCt+xAHUJatguVpwRGEFIJXCxVVqS1DTYNp4N2LPKnviW2eGEg+c0
zP3ov2UWvrL0tJA0SkhDp0IFLA+xLev7sQkcrMKH1M2165wMwrFn7KhDZrac59bk
iuxTgtBfksHcNzbnjMaHjeFyFzJLqRfw68SSHJps3MQaxJCrD29/4AMiNntu4JXB
mkpAcOcgCUTm5JVHPwpV7G7XsWMrTurrx6/Ik3Sw7+FjdB0/MaHCJS1kyjbjVouJ
jY6XnBECmVvIov3LWpe2WmRKViF3ykTuBFNZCQioxehH40k1gNZ2spOpKrnaLiZU
qz1EoDQY92Et3Z+EDZX3kOS6IY+XfzO+5xrxtSYtw6uQI7TVMsFgfm88WVcIJR5z
50GG2FkMO5dIStQj1c77F9LnaByZInJX2Lf+s8WgdVhw4nPHR/B5TRahbxO9PAbj
2IxKGRf4GIvNwg+fz9uMH9y1zah2Z2epQvCZzEBx2okPg5Y1OQKBgtqCPUMHSeSr
WxoxNSq9qdh3ssJUcxxzMlUwma2taYOgWnKhFceTChxdFKM0PxNAcKGmmPVUVebQ
g5AmJixUyL8bz2ob/FaENiGkI8U7yFKzmNNRBBMSdIfxSXpP9JsyHbdz13le9ra3
WUJq1silujKY00kApkiJn6jqXnm6XnsEKOOJupXNtW/nb1Yo0m4tBKaxyF5okyhQ
XHgvehcNXQCt/3bBDoqfTnHoeXLVFfMaQcRZ4dpK+ctyZgMgOTrDZS5dVhGtAwy2
Saw06QsBWzbAsE1j235afg3stj0xx8nqF1+PSHqiYtY/qxbMlyMINNGjQHAh4mGv
ZK06is8Qjw0O1LHJC4iBcPasNmLAvTaabky0yUDAe/e95IYsxWXzNnqExcB1scPJ
mmBbhM9DlXlnM+XJujRpBVXYyCkXQkN149ooese+G3opzy2AdJaJ8++RhErevapj
1sjI1wUUbQ2AksO1D2GHghW+A09h3tTRZne36zJmoKCOCKiPLUfSV0f//Juem3fs
BahkVSeSXKgdfUQPuJCGUwOQgtThFY3q/lmSB9xfqbkT0MHECS74gId8unbuzy9G
jIPVuyeIooPThKWGUZfhzANhPC/9haQjc/M6Tzy4x/QwjnLNJh7jbhpTqttCElH7
ZML51F5l+zOF8tFNZTziMLRkgWpxYxOeb7BNx0c+pKWQEbomrt//L+Z1yQGOH8Bq
L/zkrcXllRD7bcEb69J2LecC306KwY+Mi9RWtUMi8r7zs6rMGC/PWCHjeGM2Z9n1
qxuiw3p+WsYlV5xLiGHYOj9aKIYvNOSKUfG8mEvbM1JK0bfUCkQxePoj/fRpGaLp
wnr9o3K0NKSx2RV/sy5NGg2yfkjffQtW7oXUIxpgjU7hq8xA2CIAP1kzjEl/Qcr6
pI0XesZxFD3dfzmsz1ONLcun3lD6ianSAAcNIas7B++9To3hqzyBRYbVIWahC7nL
kKLJD6UK/FfJAJH3n/I5Nh7lBYG3Vel/MSoA95eH6UfvwiujHtQnsh2UWdXKyLNq
OjXLZggn4mbM/5MH9GgTyQ71EMhnk+3VgdxjRZlYMYGaLQbjCMoP0FDMf/8nLopO
v3MWg6R+KVcbUJsKtvdCfBjRnmE7Y+rYCaaZYkVxkePr6kG69NCbMU7atLxv0OhC
bAa8J/8NJ4WvfY8T9pgx/WgRGJeUSFP1yAIP4MUkeDFbLXuCKyibbmdVuxIyb7Rl
wu2Js+Rw74XHlrsnYJYmuj3UtbKsiUrY+IdYAUsCaCJM++maPX1LJk7EU1yUjStA
Za/Ov2O5grDRYOBXbot+dDdhezaSdjhzJlpvG3f27YiyKpIxCReYHPIBxZWC5bnH
excSZA81+2iTeRYs8Z+GmUI8+T5HxuPUvn6Khz+DKFt+UVCP9LSAroIak8BAa+eS
MVSOIzYqvz3jSXc2NLVUSZsCBWalgr3ngTuyYK+lhy/f/QPX8/vC/HJqAWk7noVL
L+3BbprE7VDt4o0XcXoQbMKXHtiA92RKZvJFgOGk/yhGt/3RcmKE6FnxU0Qv3Si+
nHxNFBtqcq/nh17D8iX35EQ4ocPA7AOl+p0Y3esV1OsdJl6Mh74BC6GcjO7Ce7bB
DcwCTuAodZM0UXHcjQyiSguLErCyIw1cBhTLFbO3O9UVXuW5a9PIKoSy2+2esghS
9o18FL+RbiRaCu8HfQAF5CoWkEi1Q0fzT+CknK1IJozRW2mdZXhZYz7YdU3C7BrY
zNetU2+q3+pO6Je8tTNRD8/X5i05ZJA6+L9KufL19mAbBJ/3MSNkWE2LcsNqjJQd
XzS0FNkDx4mjzHm/Dm+QBqVZOtTtB7EGTQZUJfo3wtJ24MbmVJYPxRdaK3eVaBGR
IX/1slje5gQF3QyvvcuGdo/IxzNejZGTsFoLqXwktqHrdjR6nbLVLTc5Q0E3JOju
r+Z/GaI2XzaBTTp8HeRgyKv1vhw4pN0C4AUrUZAUe1O7rO7bcRVd0Or2ARAVJNiN
jUWKtSwJaQhqegX2CIDLbU/5HMoE3Xxv4N1KbGE7qV/LOIVaQNYmzCUMeJ2lx1oc
2H8LpzZcNYPS6gMl2z63A0VVnOKcroHI8VXzWgClbS9LdY78x6YK616L9XF3+NBN
eiIUD6N9IewH9Oo+fUtMJcakf2b8KdWtAZL5OzynVo3X35NQ56twCQs1ekYqi4ig
6CrMQY7vCgbfn404LgV2sBdTFwzx3pw0zMhrVwefPdwnRNuSCeqscKqT9GRUS66L
Lk05rXXLz58NbPxUmkrQvf1m1/lgEl6TDFCsVX5trOV3/DT42NMw6wASgk9WGvI0
/BeOjpgcWM4CdD5qkfR3h5BbbrtzKjRuX3b7gMdZdruqx5Tk8YL2RP74jPBb0Ngx
/x0V0n1bl5M6+o7aV39yBdcnN+QsJqj0HFF0TW365HL1aOz+Uo4/k+tE94qsNsxh
LyYLTvAAyBYW/jqwT13IT0iybqlNxXGlY1f7vT8FpB94Y3Mzd7wZ9XYJSr4tYhXd
26NGh0tIQHFmT7gTbjStyL51PrmgTDGfhiQyrUOIUoPudZd2t3s3wSWbZq6x055k
1T+WjHUm0S8lgTMfzj5wJ2e9rA1zmrHyayNiHkK6w1KLsqCda8r/ntUMVHOJr2b3
4pccwH+jH1rTGLRTDIrxyfoT7EXVCbjVd4iVOJ6BeTbqJ5TYtMwawMOsoXv9599W
dzFr8oZN12eJSSpo7/2Jyyjz6sHssKagwnKkscJuus2ZBeurReCAcWdEZwsCW0wR
GejyFGe9wBJyoYsq0Thzjt1PvY+fZsQn5TBJxTCdkqnoUg/HlDtuQZBzEJNBXmr1
rxI8Prw3H9N6N6fTTdcBlGifZMrCSf6V8Fn5on1IIskO+6s7kgUxl5Sda22Bx23m
ZbQRgi8FLMDrtpzlZ5+AT+FtfcX73c7urOjIihyNWEOrELslHH3WQigP5vCmJs6Z
+uSlvigzJCoMO/oK86TRVRVj3XYEGtKS3R5s5L0CxRCjZQvhdU0oIYWti4as58b0
V3DfkwigB4/MgCJ2wXrXAVJVMii5pJpn/vHdd6we/o0XFII2xOLjTyHelDxCA9QR
9sWT40hpw3qqWNHidy2VC75jKkLyWJWlr7I290NcknJ4V0OzPlXuK8pvyiSmhswY
OJJWK+qWa3EU3WsZey+bLWK1Y64R2+ukNdxdigOnfQB2/Jk8gmS4o8mBMlkbgKBB
bfKgnAve9rLA6z+zYp2Fy9b90GY+uEZKWvgDvys/nlb2A6P9yeetTjpV1DIywgXa
GWvb53E7h4vbBGtZ73/EI/mMG6K06pqdMK7NKAN0OLOGAOEbv1cDfp5s91obpFbw
QmqTJhmtCUlLeurOrOQ9RncF1dAGbrfAK2aHDuYfJos8pVTw8UpwF2CNYunpEm1h
yEV+5rSggc7New5h2Fw0Mz30M6SazqUsavxsiEujUQty44bkMUE91AC7ooE2EXRq
9FXzddXa67M7RdbCszBpWLlm5Ys+A97LgJ0MyQBSQS2p2tww397/HoT4dMSUE4X5
zkJ6D4Cy6nd4fCgpI2JqmsJPVsqV7Quswoh6R2EctEDE24m8PZwy11scwGIm+ikt
g8s6BiMzgue7OkGtuDibd7QjOVoD1HJZNkjXVABoumRBtydbh35ytKy65wdZomiK
OH/OIQUj434mnwwXiEbzdKnDdcKrEoQSAokih20gJKjyZgNPEPnM8/rA2Miqf8o6
fEP8u/TfhXh9Rf6L+06XuDMovXvaoR55XfYq/6IqHWZbf5loINUYoCt4ps5OIXg1
68X4xRPAzqWkLU2mMcaqzhAgupw7TO+eV2rROmHLnU5+q/Arz3tWiUcywiTcbkmk
UJO4RVDm5S6oAUHXyGMGpCw4FwW6PS928dztUH/kSdGmO1TKnx9fpuEEXaPztr/B
TN2ZjH7I9NG0BPzm5MzCUXE/wlR9mPVIRNH0mjiztm0vX+ycfbr6TYf2mEbGLdbn
XJ9RVLe6vYnat8HF7hkE0b5NWWSKOnzpzsFysLyi255Vq4Nf1Kn2LzQkB5ns1EVO
Gons1cVKw9dYc3QtiL6enXGElf2WXH4Vz2qRaSs6Bb6WFmpJJcSIlVb292tXUlgZ
rzclfWmb+MW5gn0AKsIFHj040xDaW4YayT48RQZWEZon/+XMUua7dR/U9Ve6Bx+6
tZcHcTqR5Tn7L6Dbku3WLEecl5KdVCKvGop6m4unpQnow3r71mH4KxF9aVnbOZCw
vRtGEUi3W6+B9lQNqA7GgDmVqI/4uIeuLaLM19U1U/bFPj9kOFNh8gAPtOR7q7Xy
h4/aPJN2wa+qodxfTsIBgc+I8kBw5jQQku06clemNlTXOSz2bMWj7mzOA3tFD3Fc
drkq76j3Qiio8s2mqzI7wEPV4saJmHiYSh018YDXq1rXPews224QIhWwueWpdVyY
cAZA9+/Sr0RvmtuVQEcNHgue08cJVgrms3fJUV29VcmwF26FKyJqVMxXptLvJ34x
9iZSsbCybNjK+hKxWmTrd4Twe/RBeHqgCrX0J4C5LafWISbjn7uSpXn8WRrwZn/s
aaHWNnVv2bYCigpEVAoVzi/geICUYNIlC9L95gxIKE+zcB83AR7nqE4f/0IZYuD8
LzHVixUMn3xGaCpyDs87S9RCaX+rmYFI1AwbA3Gv0etMZah+7o48LOYgZPomrvAs
U00XywDoWAa0RIQX7EonAUzcD3x1LekmYRG0RqGqJCkQyJuPXUBlmw8COH6nZETW
M9c+41+tvOJWwB+UXEi6OR0xAhz7qp3GaLGhm7p0Lj+d7Le2FKd4kueBsehEx8Lg
STdl1zbhNiUK8LvR89/wZR1h0Gfj/s3UrVnrg9bE4Ul1T5xfgHcmQGpYuV2NT4/w
sY6We8Hm+dCW1nsH9lEENzgx5E8zX1uWshnXlRcJPjbAufJCsP6YiU8OtkqC6eLO
KOCJP5rNYBy269pja5pyAOE56H0snmdcLEBnYUUSoXt6OmD77ffAIvmHrBPVGSU8
88lV+aZDr/ZxX3lroUNW6ryIoxMXo250mZoDbHAfPbpBySk2/aFss6PxylJ5j84m
ikgqJVvSm0PojMhTKGXUr6AmopEyrUijJnDAZSlcu53KEVxUp61ATsnsOyzlK1bR
5NFFUbB3fn7fgCNMSsIum0KtCUYyExhyY8p8a0bJWs+FW/zY28WU6aD/oPzgPHcU
TZ1U/zlukBRblPhICrRLmDDz0FAbYsj/GmnF8MZyuObu6M3l4NPtuXA6vfLMvhrX
A5JaiL3aIk3/Y2GbyRTlyERY3mdytrfc2KVQhrC42F/+YsZ8KkUo3hsmKqMn66MI
1mnIYxq8I5jd7tfitL5Cm2aQFCnS/Xi5imaU6xUQZT00e4VJOTBhxIIAWXp0gO1G
UZ+ogSAJG+zcqWfB5LG6X3QspXGwsDJA4QlxGvhV+xze+1vLGqp5LSygMstdHxKg
2htNenmqEjiLb/+9fhMxOQqgc5n8EFf+0PPzLqg8AGFe04g6JMXKcj/3c6zJfIR4
zfV4QzyFtoyuHLt5WQyapWW/vHW98t1q+WB/Paa7lAOlvlGvzRt+wgtIbM9kOuJ7
mjrOoKCunIdbEwNCsa+QyU5PQNDiGbA1CgulNTb552eHtEH2Jaq4sKt+zIcsYkpr
NalQUkQOsp9wsZC89rIk8F4pd/M1gXxz/mH+mcicdmxRh9ICYF10q3a2WO/fA/4i
fRyHEp1/cIJ7ug2e90qH32qQeo6pDgIv7YDQoHZGblblaUIyAU7S25ZB1HX5Dibi
WcIoY45sQ/+rrqV7KPEixH8Q5jqwDiC2gcVCq71PWnRsOxD4zPoVY5AORkIwK0Vk
9+8Y/22tmSWy7aGHcldZmJecrPUI0eh9XWyh/yrWEeUhDnuFjH/u5qWinL1G8fpD
XJjdHBfgZ8Qej8OTT8YTSQPJMmz/5TRMCxvl+eo0vSE/3FvD+0Qa9E2xtNb5KDvx
q/EECMLGlIheh0qTaQdAVoHQ9IuPMlnd2Ptp6ZS6FgNombsK141sgfCqipZMms0M
XH6XRn0wUW5Ss+j7mWfqpmk1R7P/yyz1L63IO7oHHjgaeFOWUzw63iey3zaWpvOt
pG8RGG62sFER2Ze/AOVMHWKE1a3PX3rmpKn46j0bXmY77pQmtNH+jvPPy2fM3lFS
f7lPo6YIDd3U2EMa/ZCpIKcpoYxKuEo7vl9FY/j9Q5/OWPpOBOeEF9jMWj6ZHZUb
QLohJKffsrowIQQRJk7Xz66kkZp1BFzt+WfOeE2jXbHwxicqmnRB5Y+E5L0b24kT
suMD5g7ePP1tLTy/j0xiYnEmBdQb3bswBTeLc+4yGnaV0S4PfhZ3aP2wK6k01jKQ
iZiCEEQfsrBUdlmXYy5QdhP1HvGvXNq2ihn4P8CO36u3nTVSRroZpH5oGf7xdCiV
Mq23RyY5vFw+zSnWIZpnI7YNEZp5sTKaBnZ8dj80yhGx6obIzHdH5b3s+19ua30K
vB1Ewg3WKriMqdGTF/Y3xUkxI91R4Zew69ISMbCfYi87A1RlJVamNIqpkMMQuI+4
axaruwpC05vcSCYEnbiw4MSV8KNFJ0Rm7iswBTQHiO2Z15YGCicCdhYeFHUlg1lo
tAeLsHgS7QGHgVLoJOCRk2clv2sMmkFjwEkTLWWBqvyyq9B/Ua4nIAZPrgv9inIQ
aXB8LM78G6YPD5s/5vVxx/P7T0E4eOvHZCO+bnrK4g0JvQccpe+knkdWwrKGtfYI
nx7YaLL0oHWVLqld7S2/MwA1j2D473iWvjfO+26ReMKa2y5YKGMtNurgke7tt8s4
5fqlIzlhdPsNuF615YJU7OShzYregyEASJR+Kq3NhXTx46WmAYVT8Ya9oLiNRp/c
r5aR4gL1oqMvk4y5YLb79rHqgonO5GbUQGiXOkpaOS9MJF7MD9NwK8qD+yYucljb
7/h6WHOctEsvuqhOmEHlg+Dpw5kq6kKWIxyoFKSebWZOYFyFjLuyQR2hF1TAM0sj
rxjviz+xRyUnbkk7F9/9NljC8AwmacstAsQVVgAeAzXKk/iyHdKQRd55kdaXPhc7
tOH+JzLSWhlIuB+lxw6MMVAkI/SUzEZyb3B3I6U33xxlNfAokUye44aLoLaoHtJh
cPIju/CUOkB+c31Q5LlxhRMrEQum2kMXSeVH0Zw6JGRtVtmoD7YlFxzRR6Q+t4hM
McfhEI7A6akMXO84mPgmCkbdVvPQQexac0Eb083pnY4LohLi1chBqjyDWQjOX2am
2o4lADgc6w8aZPrYCJa1OAdm5JxzfzI8QyU+zdOHPpn2mwEzEBNcaOrbYTVthCpz
fY5SSxHDrLY1rQpGvLFaM2AjyU4+TZdQ3bCwIfnPw/JdL5MXmBY4/hFQfhD7kS2U
iADDs7XB3b+Ux/rI2qfGCE1413wROGF2I5v0PAppBfk0Y620d/Y5vAJVztL1ZIG3
Ym0wct42cRAarzS6Zh44SX0IebGnIyREdkIGcQiyCMsq6DRVA1WYsh+ecfEiPs3V
Hw9kwZ6LlVtn2CRVDLJaSp8vLQ8ZLYWmi053mHQoXIAdAUkr2Ltq/SzfIUQn/ATi
ckdbFkJPJtmoWpwdHD+eWkumovIZrZaPnGIzprOZyyG6vDfFfBm+tri6Lawd03jS
gDzns1Eo7lDJfaQ20BM9TmzH46T9yXZhL9M7cP+Sa2JhOup1mFjWi2yNzgJ3NRkD
XqYNar6ID9PJW/3nVvuwKL0QEe2kYhgKf7qhurtVPfhAW7Z1JK9kyOBZX9f3XbKW
NAdQToJTsUpDEMBqxqgvxoMfE3tFHUUBuxyFqy6FuCDW0BJVlPG4NKz617QpQdUY
km2KeFBf5KgirjfpHjN5wcnfYfUDnK9QDOZfdvWYMLRyV5XGYYBVIhTGJehyP1m2
WGc5K3J+GCX+sq0soXAAOfzGtzIW37OqdIlZwSSb8bSdhqNVf2X2ZNXo/g7R4mer
gi+HgURSxw703hr3Yh4NnDuhvIi3RT01MepZyU7Kdy7ix2K3FT/iXjzQIXxjpko8
H1jlEXviDXuEhNFnfIERRkYYdoV8RJdVR3pWkb7cEokLolJOKEAYL6iZrwi9ufTk
oDA0l6te/pCRF9uzXCCiV0q5ZQUhmvRRXP4oBCIoMsJ5oU4zoamd1ObOt/9HXn6a
DjRpq9exDSsCVpngGKEoh42koMmURZRajDOQnDuBjzAhSkRDVt+9z0aiy3PIFP2S
+XjaboPVSELpIjctlLy0fh6jYhty/quT/a0EdRCNvKDTm+71I2NAaOSNWUFgN5Os
zRUkQU8BnZFzDYkyMb/OtyrAmRsGxSv71Ghrd+c979E3HTh/gejZhPjYBtqUF9YF
47P9f0uGGzxRvqpIC8kpIuMV1rgEWkK4dMBVe+gfXuKR4u7pMM7xuERStqwHFfY6
FLHL9GQ2ssm2JTGf0ucXf7XrUfz0w4Bzi3lDO9AJbAIe+Ufkj5QHWXCOOVZYrlPt
XersVRuQacKY2Ct+f8YU6y2p1EW5Cja46+OIwF6irrfTOQOYc56EpzjC4VOsc48y
8GajjD982klFtSgNLcCimF7K4a9NiCKusKrMq85VjzELtLX/t3GItwHLUWPpnHqX
SJuZj9Ha4f+iOMcKPnvMvrIqa6ys+kURLctpdwC3CQBqrfoYImlXCix049PtnRyl
ufi1jS6W8VxQwxfYMIdRCp2dI5skibWKZAQ+j03+GmJq1+J5L0BqZ42Av/bNW/le
C9rtwMlXrDrm5GAZzjRB8Gr6EM8j9U9BfWhkK+TwOGQNVof830F3y7/jqIXyUrdU
Q69EK8xmKRmNp/h9eBw2UcF9M344RJsxJ8+e984utkCQh1UG9fBIClUxOXpGoGRo
9FL9ZsKEElgOs0SRhbkR4daoX9T35NW3OX5S+3E6l1/d0ZVrMWxvId1ZFt9PSpns
d64G8gEbLrdOHRqbt6WRa7VXs5LQvsMcWB0BbiAByTmhiEYzp/GZY1I3bEJZ+J1w
ivsk5aqJAB/WBeK+Hifw2MlmJ4HucbnbFgmaolf1MKieD+CRT7vGNXzwfjRr+fPn
FQz31Nya3bjRrQP1leRwCunaQ7opzAuP4FZR8T301wFF9wgFnjGissQHZuc7kP9M
LxUILhRo6vr9i3IHdX6LlKrdrG5/pHdUhTx5krnh34UKWMM2ZIMMjJpZsSffrphx
L+jUoxvcp+RqaCg8VLIYvxbZxwR1Hw9VvardnAUpS61vngj3poQxD50AARdd1WRG
KOfVlkILUTX/hwRa4JC988BVQ9sdXvNzvXoga3rfPYh0zvHiIKQ17XF2t9u4U5pW
0fS0QeeXmRzplCVXI81Ad4Ks/z1YsK9+bZXfZb6L5FMlxhVeQimioNherMLCP9Pm
omI2jkbLw8GfeUQzLYcwAiYpPeYkrZKh4Bvcnns+SEwuFogbo7O/xOasaiSl/R4S
9IV0uNMCJGvxbaq+OG2rT7KdsHHLQ+TUTr+lfGtxIzFup/AVdrXYRk6U8gWwcI7A
sLvbjb07COZQ6KW4WerXrHbldNSk4jT5mSulK6ORpCJQTgDRaRXAkl+YSOr0vjnN
yx3gaTbhioNuw114unH+ZbwXoXg5dZ9x4Yb4C5YBdzedb2igpkxJGlZY47UM7IuV
O5/kXVViyoYR4XcyC5eVysODsdyAq2SdxmfrCIOyWi00K3uxJvo+BBvag+U2t1C/
MBaZDZ2s7zYwXmkHi7s+/KYamuw/6OdtQiOWj6gyzjfh2XvllCdn17E4LgOjm/xu
tP64gHp+INsrxKMkJBWqEXLQY5Yv8ctwIN5/3ylboYiCLblWKcB0IE1wTQpU3yf/
mKwVV9diMlZVb4KGnmxjoL5NPzL0j41Kw2Q2TBNTvIF44vrYDH7/T15bGtCLWAW/
2nCEE7SoeMO4jmbQdrcqxawvMdobO/3uzKYxA1iYdsxIuomM84RiLuww+pOc1Oa9
6CkBLsINNFk0B7ItLWIS6fv+/Xe5t3JVFcnxq6SuTitbQunvfhrefrOFK+MW3wWM
ZY57UPTV3TwmFuO15QkqAVuxQHPR9nsa1VfQSfo8lFN+osE7/F/ens/4udTSb6ZG
iBKMSGj06g5oXa+6uxP7tGMFfpTRPOidCVMYMhmKo7J/oO72Nfn7fg20nCkFMU2j
f9DPf5yGuUCE38gSA6Tg1Ph4d5XZaSc9F4y25Pptt68AnEZqAGz+JW/wkFAQ7BnX
v1T5ZpXdk65XOXOcsUEzUVek5esS8STD7aDk5sN6x1q5PQQCF5Gk6pJizoOj9aZk
/npye8j5pCuEo8sqLOaop1vsGe96naiBqXnUxyGLua6Xt67FEBLRCZuQWux58XOB
FfUotFEtKZGakT2Oa6BUDXs5x8rEeYZGx0KfjzfYVXIwx3nSS8zS57jQ9sGGV7DX
UoANsA9IHIGRKfaH0nR8/vlypBBo8gd4mc6B91KYb8p40DQ49MPjDX01BhGy7DRk
TmZHsuZACGUmSsWl5jZXn5rRoLX7pgCqjHQBq4x8L4I5g1QSyF7bdU75aU6Dh8Fp
Plk5eS7CHB5ZjntLfMmL3OcjyYfhH6CFhg9P3EgFHNst8tlxboyNQKVQW+sBHP/w
gn80hi33g5v39uaBZuw5UsxmQmtC2r9kGX2prxUgcispagcC9m80zySxVSWR4v3P
tThPrx+iInI9EtiZHlm6I0Zo+HUrbfT6VCh1SojBiXnE6bqzagst0yAHu6Kcbngs
sJTp8s3F+nT0WTMznrGsellpuduGoFYmDc0cU3ltT0fAr4TKnVEXbFeIeHJk3QJP
waO1vctzBtiuBU7tasM/kOZopTh/Ey/QFH7ShOINdlT49Zp566kKRzN+OeKeu41O
hCDJ3JjmSms2crO89lSFz7f4StqXgsikXhXXxyCLSVwtLDr40emEpyJWtmyljSWa
z+MUMVnO/ypBhUKU+gI51wzq3EyW9AK8rccAwBU6rtJVrB4V4cfepvc8f4ejCqSV
O0NCsRNyRONN6/BUgJ5q5E0PdzITB8IUwXJIXOsGiZPJ6RUfdBzyyWB8UVFFNBxs
36CCXksyKm9ikQd15heIqBaby+CoGwfavrjio/hUW0dsJOTRH5O5TwV4ayNqtaZG
D9Q3DcFkhAywH/ApsmJuFM+KhEyrhvjWEwJA5HBYwybz/m6k5oJ516IDvXmqTcrB
QgMOoz6zlBAHkfDxIGf758Hb2UPI0ZKXXHOULyEYgnyaclpJklO0/Xe4jqXG07Nk
H//ejbX4ZGhq/+CYu8eLxpK5d6L2rzskwVG2lsnLBm4s/uggILrzNNUV25qSaxci
BPRuIrwMM/4uJxZ6K4DM33sUJJAYTJEVHU512ISfDM7BKETglz8RZ0ixCGuViota
mu19UIStYztisV1C47saC54fmiBA9fKtNL26a9ePgXlvN40/A1aoEv7EoSk6yzd2
+sFDyXzkV+E5sHv6a4vdMTlcfREQAIxDBz1r3vt8H9ujbRHgVnYuq2h2yacmyUVJ
Aov7EI+kpOdpvm5IaUN7gpzz602u9FcSuMGWh2jKwj784qBv3kMbriOvB3/Hovjp
CJ8hFkAXaTyhLD+yjR+dQg9dOymSBzqsP/ld2y+8d1avVHX6goUSMciNOWlOotLN
inkX26T3PCrjSm35Ht9gmq++WYC2JndTiBvL65zoTSJXCW+epVpC2grsTd6BeF8R
DJ9iIPKvi0l7T2uKP1t8O4AmcSKwyg36MgH4zDNu5ctIAxcbJpbcqz4r7b4DdKPn
Ud7LSe/u4B+xIBTF2BnND2pdFIZWQGOC3xb6ie8+91ZaMc2revCNXj2xt+MiU9dH
c46LLse3xlSTupB+FHOZdRIWtHbufmZkkdbiijdsQ+ZKy0oTXmtOxzOBQ+siV1KC
79nfOunxZ1qP1ScEyWuFRUxa2BX7pCnLU8bVjLk3ooQDSsZBPMXgdAEEbYZmkBGn
KP7/FHee3bKOrbRdo9nu6mERbHNdTG19MD2dbOI5SEMDwxuA7L5Z9U9dZX40C2u+
C8Ni0KT6en5B6jpOOyOMQO+3k9468SVBMGyExK648R417JDVMoClpfGvQeh6N3oS
7DU71tm3psv1fV2mn0GDQZAozi7HzdZU8t3VXmy4+6j+0xC4NZa4066kziwLEuIH
92GQuIDyjgpC9aeXMoTHBxIlP4Qb8125aKrrQDmRJVWUvaX113JU3HsmAvqdgyMj
DVtCe89iKq7br0Zv5rJfc0AAppMD2/Rh4VOyjJ8UGw9CAf7mP4nDoUVf3/AzxttZ
/cyT5qArqpoMMlBFe8a1YJGQHqtWSllutSF/9igLTWygMX31stJhTa+5YLf5ah6L
2ZXQqDCudefeH8XI3YawmSLOM/O8XhA+0M0ubTqqbxMQ+Jp7PlAVgWWWiluB30qA
IDJTt3wbb6HEkiuAcKVzQ9yJiBB1a364o+m0uI10+1PxONVdGImUCMDpK+6Jxj4E
LDhu5vzuLv2BYYox3xq2utuFsfpUPU/kJLiJlKqBB5Utjvk3FXZWMaI5Q5edi1PV
FKnNl3kx3J8gjmYhdXgA0hE3Ns7eK6/6vS5FQYdeCtIHGlh5IvYW9V10fgmTGAoY
3sKDyN2NOAzLdl5lV/v/AlyYaqYSYS3cIIYEwkoLTuMTxmtsP63uSMKyBYTOtUG0
+G+UlJFYZCsZygHGbQbXUOoRnsnS4HoqrmUs1Ugf3hSZ/2gi6sSTOX6FXJLvaxJa
WTag9/2uHXPFOTWcw5+SvfbgWx9EUgrx3U6KHK3yB861UTP/M6HZZSLlPibq5Kox
XBPAXYy19QaC5uqSq8F4BHvGKDiTAAQbjFF1pGUxlNBY8iWcO7bAvlIFu4WvyUGy
R1toSXWOBbH3Ita+MXJBnwfELplFU6fJt9bLgKR6tKwcf3bj61HlmpQ7/1sUr0YX
YyKOVFaQ6b4V1AVjAoyLj+5JGrkIRHy7XLU49mSzi4l9Bt4Jbg/nHyoj/vAAlO60
nNmxJnfqw1nT9tRPEzcdpi+/NADSD7/mx0bcmknIkOEZSWxgLsNh5RHREuyDi2fn
hfaYGSzHG+7aN5muN1TpDI9/IOUb6rRwb6WNzWG0R1MHajvcbnY2BTfaaZ+KUmo4
NwHfDb/sAmns3a4XwAk5cWx85vCN9FNrdulpdB/m0B74M/UElVck1PxMPsH+jIDo
u37kFen5wPsZxKSd9haBbbbeDMYWA3w5pfHTl6Bcyj25PnLJnyN2F/ciUAXjNJtX
TzIDq73Dr4dYeV84IFyffocxp9/qBGQGpUoK4M/nOqer5kLkeegaS11U9jYYcWeu
n4aeNwyd5Sxj2RMc3OE3j6bbImmDGpNJ7GoqppbOkUKOz/1q8RBsP60UzDyI1QtQ
6zoC2jMw39SF/U+T712yLDrpBYD52a/qfsow7SOr6W8BnxtJixkFWLvqdvIXArLQ
NFrcFhz4ErUNWGvDKfkxTLV6fSTenhgaivWyKMcj+aId7870DACVO2TcNPfZroac
dfO3/+K471bLjqFnDvKGi6q5lPiYKkvfluZrODccepDw3YxcM/FoH1E0NkB2p7Kr
7PqibEM0OJpxoCoELlihE4cB1RA4zZrULiGBGH+RySxIXBQHWEKhQnlwALvsFucQ
DrLEYE3KqJH/xvHZdDzkrwJ5Syt4mUL34w+ZvvNTfCjNSpOY2y+XAZ6FmIMc6BLp
spswhb3wgdAFTet9ZBWgJ4nrjAusETXJ0P1/22GYmCpIIF+gOUyPuFG4nqL9/CWI
TwtlgbYXNUsS8rNeiQ2GYo4r8HaGLX9GdCqF+9tqNfeMJpya1QstLwPxKeBs8ekc
8MooEN1GcnLzKOrnVQuQziHI33S5qDjXeatTYxqhX6As4q8nnxQwA6yWL/P0W+YY
yEZrswueVLnEfD0ZSV4TSn9pV9FONnPaeU8td34Me2XVXfyFUzxxf44CC9fbHaTf
DSAWBYNZLOr+n/jQaiAMkuOkBJE6GNgJgLCLza+YFXvcamk6uQogKNOl25CFPH6O
d5uqDj91QHisXrifLjavJ5+2dWZ0rm6ZpLn0qabUXkxv8ldr/RgBxIBXWcAmLk7c
CsYRXymkcMaJ5uOiLSygaiih4aQdgVTiliyIjYuCMnCfBpM6i1mF7SCvuL+WPH3z
B53q3dSo+YtolTZjXCiF4t6RTk66YAeSlKuJV/qJRAMnkkmT/qRy11RW6nNGEkGH
i53FOGFgel6Mb+ZgUFQeowaLA9sZjD+BqdRuUdyAASdacX/qm4EgLjtpbgqqL0Po
9aoN5EPFlNa/pm4agsRDT0Esoa+mJNMnh+VU0HKJXy0xRbBL1oLOUYM38MQtg+1f
CahKNVl7Dq3ZakY7U8f0xaOD+OCRQ0A42eQLNfK4u1Wdv5I/TJg1Go89eYDaPa1c
OKuDdAhhzm/XxiI12KzesBlgfn7aEGy1qGLkBX2dt+15ldE3pBRQJ88CXZ4IRNmR
beq9AFBH79rwfw4svEiDizhk4q5Ei9/AQwq0mG9RUtrBA+34Iz76NC98vYeiSWT1
R70cfeYMiuKsWVjgqktCHVxEBSs9po0blLSrvcdw9N7jgIADwlt8rHkusVy7dz6q
ROSQ1woupnE6xckY9A8prv2kEimiJM+yuf+aLvKYABWaIRr1OivPUPFKI0ztIyDK
9Yl6ozR6J1aFcS9JPf4UAKMMOi0xnuuo8Oy7H2LKvPELGEzcOBNK95U9J3t7VcNV
QkBTXhJIxN0aG14JRy4mmyZAk+IJXPHL2FYd8G24TYG8uOLECzG+i9+yDfgQU3WZ
EYh150M2IKu6tuZi6+iIH3NUUoV3q+5yNrdl5bQHy03fjnhOzKQxH5+fIzW6jnmF
GwBJ/67tKdJu31hONawl1xG2OChSNA/GmrHvDd9pnS8BDl3U/kTgm0dA/0ZiZqLU
jka7J9vqGpQwlBDRM0F7KSLZo1uG7MGv5NiH/OuRoYS/S9JK5KjnUexyEe8CsO0K
UNNKO3sCehjX3G0iCRjCsEUSd/fH2in0kfEjkhAMhEGzAxTwAH1TVG84Nu0KPnHa
7h+lD8mVI4Y+3LqFZemm1rmq92krtzMyNM5YYYP5v6b2BuMi/xQMSkDFqjvDqy0k
RxCCOHSfVAWSy5gqZHxUspYdSsVuuBEkKNtAKcNlBW+gBMaXe1pkQMEp7HJmTuhD
YLp3ZdorByVWnHqFsAdj3XKhwqk2lEJNPEoYk6lKl/n3jENw54ZFOO2Vi17z6ibU
pyZyombMKpfH/jHwUIWeGXRFS3PKftYiTNTFZ4QR10Fp01M7v0pph/PrPald7vZW
LIy/Cxhf5j9CcfMOG35tB0QDElvZx5so4a4jngcihAVseGCk8ZGn7t2L599pPd/d
wj7ObkYikvKxJe1OqYasxfmdN5wXNSFVrXdJuvkrNckRLjmpJm5xwD7XT6/q4piO
Lbrc0Y7ciQWuQ6DW7e8cmB+15/TdtsPVRNy6C9GOPevxJGbMM9kNVvRekKKNcYVU
jHctZumE9OW+O66w6DMbfLaad10A64EeWqjZvVlpzurEkUUkTlS83FrbZb9WLnY7
807pCf3B3NqFAMfTG9/EB7c34+OKqzKnZFRjSs493q43pLCkVEM0mJqiZyTLVc4Y
uBj+p9oC/GpmcIC+nHKDHBIBqKEqDeGiWs1s3TU9LFYNTGpg6zTPSCO1+VBfTgKZ
V2YAIi5gP2raofaksJEA3TZJODdJj2N9aRYJWPUSnhGq6rShevM3bMDVOaU8Q9hK
MwQtbKoAyGZlT7tMNbmFhymJcjkpvZs8GkEWQM/QV2ZgWxY7BLKO1JMk0LWXeIZj
8NgowOTqIrMmIhl3e4abdH/HgcWAaKkIdKfisdt7fCaarT97l2rtWVk8SZMF3l8U
gyi4cZ8z65fjzxcTqyUrM6hS8XcF6XExxzPjLiT0kGLYs46GnPQXCQTjviQR4n3U
PlENhObgAYf/+0CEaAam8f47ClNI5H0JydmRzPWOK3A4KxNlV1FrV5YIsRM4r8Uw
58XPOdOrUCapALU/fPhx37XRDY92k6ft1v8A3dbHJNfZ+NsgGoqZWbg6AogDYgVd
dOy7LYUOzxAEfnq3JAr7q2o+SOTPPsNnOoQnauUIOOl5QHnX49yVsrwTQxdmXKwI
eIAsSdovPBDQ/ROST8ct1cjYN4BnSsnqMS9enFsZ1UCLDfn66ftdofnm7KpVhqhH
nWozrjLUKCOMpMXAEMQOTmfhuuE3kM4WsLr5W6jSCaetFBGEOQETFwUQ8FqMRU78
RGmx6EKLgl9OwkMWm3tbMbovmHZ+2g+r8Gh5Bd0ZYVafAHSNxfSjFF3REwgzE7cx
XvXUayFrjThmADTIQ22G/kf6l2FjwogZ788QKnFTK2G0za+IuAI9+NCm5tajMLdQ
i/p+C5YK3cs2cXQsDfwJe9uG24C7KwMqMNfYM12KHVYTaXnlYd5UWJJj0Vig/PkH
AMX5PRoj4B338qdeEzyNsR+qdcpJkkbAZ9hSZfxCAo1vIOISsWWHQJ/gzaqUsVlf
YQAPLQASI5K9zVM38q7jnMauk3+kqVmbAt7Eo958bdmzR4NFJUXV1xLa0PwsytPW
q4FlS8r8bYZovPTd/yCHp+EzY2q4fESi11iIuojIF8CBbhWeaLf0YNvCIJgSSxSH
au8xi2jskpIQfhlJAWgfbZGNvsGUnHLwyX2Ihvxu2tiho4aSqMNCxXKhDi1HYcQK
Seq3+DGxbblGMkOOBCgU84ZRnBkHWDPfb9oZ6yzd4LNdRBm7ETizBegMmun6q/ct
a3/zIxC9MTZxBlFeVPRkZiynlSnFtwet3AQIkJjgVMohn4/14knGtBggezMg64tD
/CewQrzHMTAl9kaynTHlcLBvl0BbjvN5LP5Lh5H5TL1KVIQ8YS9T0+E50yv1GuZ8
SQaPWdf5nLdF07RmWCU9bkNmulBF2mpq4nRcsv0BVyFxJfDRuBirYDfSsIFsSQ29
n8LQ+q9slGpj0dYCCDp43fJskhaPEw4qaAO+1MT7VJ88qRvBXgEEbEonZrvCQg3Z
ahaxJ2hsOiKB2T+C3IJ0EayymxAKbLfs+IIVpKgAeX1PfnW8Rfo4/JvnxFBbt/UD
CFuMWizvZ2Sl5fGn2O240YT25YKcp3VJH9481f34TgMa77YihbLj+IjCTwsCTnDD
BoXLL6Yq7KPRy8S5Vx9fg82k1Yhrwfus/GQtIznTz6TbKpkMa4ryvqPneiXnWfUV
OlWJ3mxxBu1h7k2N+VBtZfcrk/hN/sfg2AGjxcGgR9YzpQSKZF5Az1uu3/SFKn5c
kPRr/JaKAUdYgQjIh0XLwa94ulkIoK+dTaSP7vUNcB2xc+VGFZ/e2WLwxh5uiAeB
mFPAsPmAFvKgAUBAsJbXWN0aRvaPMSZddXzkBFHGF13eNKcyeAPMv7pF8eoxkP/k
LO7o1Nix2PtVYwWBqrJm+w1lDs11jmjokAYCFl0oD/3GyFqAM2TeyWZg5LAZvglt
HATmyxWjWbN5atg1M1CTS5jyNtqH+W63IGmUaLT1FX40UT6NVjNCZu6ikEDruE9Z
4wz2JrDRhXsBGTBGS7Oy27QQV1KAcmTw9FmnK5Xvl2LOu7nuH/TccA5V2m6iaJPx
ilR9PdoyJTJrNAN/xwb7wa/gfy8sMNFrthJn0ziqYAe1Dvz5Jgy0pM2GivyLKlOh
/yKQRHTtF0tumjmXcOH9yYIjyP1lgXcO09jTEYUwYnAmNFnLngVPmP1MxhgxJts+
pXZKylwtqb6aCYHk5dzk4htHeGT5CM67OFfYVP2zbJupOAOUZyYAvLxfMy+Dfd3W
0WjiyN32343V/h6MAMoX0CvDy58ZdHFaVH5VzmU/gkdZxg/XEQTcVaLpYwpy+ur+
LpqYOIK+Uotj/dpqvPgdmy7bfXhLHcRTkFutLXD2gH65NsjEjabtLMYu99VkAWGg
vxSvMrw/fGSj35/oRHR1IZp+PnpC1rxhXKgPYz0hMfZUQ6V4yizZJoqJX6D/lefo
f5yCG1DjL1wm2JXC1UL8hghRmzKWe8TArhWF4qq3i9JogsP1M8kr+yb1ULcae3RW
ji/Ik6u5Ar5QcdYxBw4dJD8rtX/SEPxWA0D3+y3sRIGtpfs7VcMCFGyAHA+/URKL
lA7Wr27sgpk/4FY0GyVxpdfdfkuRA54iTTDPYiYft4bdRM8WaePqq1U90Ut3fg+y
0sXfvxbCFCTmsJgeRt+sTXW+voHYUfHQN8NgHlHPBh4VA9MnWiwaT1UZoz8OaQZn
m74UvFNxSrMmP33b+uV+sADMuxos1rY0yBDVbuC9FvRRbKIcIiOJJGnUIZzten1E
W3y88O3sD2QUHmDQsoEDzee0anqOe+JFBjamG5uWg5MbevjquasfoBsNrboG7t0b
Yg/qOKhu3C8/nsRVd7xQODvBsnI0o6k+psYjbiNANRfhx9HNMA1gExrEdaMGnuYF
YwgxMG3LDzEMXebQVge3oKiFS6vdV9Cf5GHBg6h9x9tJgHWFFtzf348GW2bv43KI
uUOnaDfPRmrhy8hSo9L1VDoXJ6Q/NRI+hU4/XB1cHSYXYJ+WkonCPDItUL/oaaf8
VA07/6eibM0O7g4zommmXg9DnhyhMNS7UvYZccmX7bJ1tvLzaBHABIeyhzst8rQi
XYF9/2xmjQ/OcOoyBcUCSunRgCP/CMWjaG6fnt2xQ86b4ZrNflCIWszyiuuTGux1
MlNGkxnFPb5neoANeVgwQfV0aAH0kcmufBsp+m2oELYmnFLiFzIeK5t9P/sGY4Ej
Ld3vXYnoIoS8zWYCUAFYOZrxgfJtqf4v+i9gTdiFWsBx8eOjXLqozBraPmnj6uTT
YZ7msY1Pj75hlZp2X+jcEtv0y7/z84E0SMYEHU857kHqwyIoTerW2Ve7S2WfBicL
tWSeEZMC8on1IFkvr5QQz3T/PMK++nQKxwd6szxg/eusRM9Z2ryf/U0OyYogoAWT
C3hYeesrhCTyZb1DXsSRbTGfdnbjkUoMSfLGCkCWiWsG1R+DNDYmdXyLVqiH28F9
eYA89y1nSgEpWPI0FIXNLJeaIKNrPB+vPhiaEbXBwGl9KRvWzb7N/4tNFI1W/sO4
ztm8pK04/t/ZIpskfVuSFG6LztFuS4t+jmvUhTEIVEYLkVuNPR9ITedZ8/MmaWf0
I6xJyt5hVZPvwDSAXU6KHFuD1djEY3KcR3vdYdyi2gPl6ae6u91wRhU/BNKYb7YA
KCCOVMyi7OU3OdEVAj5LIO7WI7c8w1Nn7JH+lqt4P0spjC67EntcNk+KLpTEXzsh
Ape8vDrxP43kwLklJ+y7jkrQUjlFO1uxIhDHAxDT2j2+MOrZba4KBZcs5c3YCnwY
IqIW+IqScOuSYxEMJtVGEu7Z1js1cZ0R96mE8/MhsfWEvo4Cr8MUpVKcb2jknxhx
busDHAf0m8RpkQMg4L35j2R08qfIXtn8ssf1dZc6hXKEVYY4/rkba1ymOyqQ8XBe
zCTMCan7wePNlBQv+LNVyX1j8+13hNKTYT7hK9QQ3qZTiCxE0krT1ThH7WEEXzWk
rHDnbACelk+DN3EQqAG9SLVX+5QlBzIzGy0ZpmfcQa9DWrcmLBqf460KZMh6QzWZ
jJJLGeNcm86vUWyXkG+t5IaJG7BqcbQoZPb+JzvyRL8fu7+CApscHp/HUC5SuHMd
tSi4M73wbrmyj37woq25h7w9bYH80sMauoRzNqwBCnXPz/5jw3jyVP+/mh6TSLv1
Lva7S9l5awuHP3pp0VcOLHw9YQuITqtNWhcRGMuirsgbiZ+6lezmICBcV6p5wahU
Q+C+xrqUDA10ahbA7DfBejAEgMz2zW58P20PwV/wpWcrFaNhVuPsU/yxABr61noD
V5eZ+W+obk7UEIPzytEj9cp6keXPCu3h0/hnmLf/WFAKCo+cjPnoUPA9okFnYMvO
jcfD3tCY+WsTdahMiSVJHA3ysI25oqt4h0lGIu2x8Q6KoqebFIZmpSisDuoSFj1V
U9iZgQEghvAk9x9bMejdYF1z2lonYPaWFTG3Qsq57xgDoRZtZiY5j4lYC6t286p4
5Xc0yTuPPFUnSo1N0ylStjMswrvmFAxA7ZQl091u/S7erzOPEI5vPdZXrsCkUZTA
7M8glET2WVGH7F/pFoek04dCi8qu47paGVTnFuR8qFgi6aD2ZEyaOPNxW3Q6JAfh
WTeEBOtWQiy4Rmjcz+gVb5dRigxOIQF+EOzWcYWGwbvOAaRPj8aXTNlCvjFnBffq
Sj8EeSUGV5O6tmmUxAameVKL4GPxlQu7uRg4/xnw3YSJfVxCbtZ65u34DLKrGC0z
yOP+17gFdcp1U9/yy6IX1adl+RWYQoO5kX4s1cZiCaUoobE6dr8xzRYu2POwPT3v
2Lt12hHxZQPKRlVI17pbmIWDHkWoSAZoB5GhP0rRByfXKgr93PR3ouNuy465fZMi
ppryGyVxSVKI/xUwqIw4D29IhXG+jZd0PpOIS0RrVgKdLiFT31gCro5EwvhMWTDd
zwGVjLoLiDcDSse2lxNahZtoFfEbESwi5LMmQCxqT/I35UaIeJmKjGD/UQXe9wg7
xvNAWIHe+JtEXUaAJxBFDY6pcs5G+hlacKwfnVaiZRLTrjqn9V4YE2B4RIXm6KTw
dpnwB+J6xfJx/I2M+B9hwzBPPJSTCnbvG2UOEI++NzxWos1lWnthpF/U5l6tjS3n
KpWr5bQYbN1w4ECqMRFNJm0RPXKEcr36Hntnk9KdUJQdHPTdvR2J3BwOBEIu+Q3P
m57YnL3eFnO5mtP9Fok7N5V8O1S+AR2+Q0AS0takqY5Ck3AJ1iajqKm+v4hn4jWt
VgGjb0HSObNugWDWw0pMDf3ZpcddTTle3JYFZmYRVkOY+P7F++753sPpvfgsqJ+p
wjWX3QrozjdTIV7EVqpPbmYz2YnF1kfJPBKhrRUCviBFFto62vGwayxaUwuuAXY9
nrnb2EC5D04+nRZHP5cbmcMcSvw1zS2wGLY9RY36tVRbdnwUD0Kf2ycjQOA6EgAe
qxZH3pnii6hLjSXfAvqQ8oGY7PadEoj2a9vpC6FZJE+c1b9g2kOMtRVSGbdYjXKq
3HiiFB6hcjciECVOOeWW3eov61845ooN0pxZimOSzMIcwW8G7HLBSGMz5fJQ0ZBh
HW++/TNS5yOm8Bzdyw6h0CzoPcBDhMvuHolhSC7ZNrhQ2tVe1zTdepzncapeLNZG
5muIJKMhEj62YRTfPt7uPPXWMDcqzbo309Jot0pORrKUOcJjRa3BLH8460WsS3d6
rgF6N/+QcLUWcrv6SQEByKKOqOw/ZD3ut4A7HOLwj0TL71NY1KmxmJHq8Q+0Y0OL
tB0fcYp0d0mLCWYZKxwMrEcGGxokHKFCxqLW6yxUlwjvV8FaLOxnxD4J9VmoYMVW
LKxgjUDOsZJ2edO78vHzcRGbug/75dVr+DrV/tW2DnNt/R6X5ZdPTUVxvSOqzX9Y
Fa2h7aeSg8xp7SXExPjqlmfyfogPJAp39vzhCI0xH4kIBm5rBi6xPj7dbOSpF9xX
mCSDlkQFAzWJLAjWnZgHknldPSfXZrz9YO/cxXSvFgKI8O4qaKArHqJMAQTA2A+1
BkZQ0hThL4/8akxAoBgtbvBdTeS8vkOSKIZOjKxTA+737Ax5CCCVax5qwZWTq1xA
k5UxG8JQ+x3atQm9b1QqtAUwa5cWaTsIEIL5fNAHHBgR0EhBhMGfJpjmQec6HAdV
G+9uJ9OX/ya21DdhGx7pqte3i2RsguUi/4kQWJShQ9HIV6t8ThLd1Z81qbitL0tC
TfeqAl8n88HiTsK91wUJrGvQENni31YyH93H3bLfVxHJgl9mx30i+qvtectia0lq
tfNyB+h7cXOZm9U/s/sxyRU5W/fpXuYdLYCiqr9X1mCUlvt78UcJRliONdcCMDK4
vAoyxSRQCE499OIP3pR35/Ee3k8q65lPJTWiMPLk9Js0Zp83AFlowJ1EW+NfnTrn
+w2+A22rO5Kq0NQ00jbiO38U3LTrECJKr6YC7sS+UOavn4NsQ7ws6Uz7WUhwGiIy
t7UWyIfHGKCLRvz8q3XVSxvkBp9yQfbLKj1uGVBImfZl22/wAfSmSPdDPH502w8m
AtphkdI7T7NuWIahvdb3qyxFDavT7xxRzomtWfzdk0wtYqz5KgVu/me5UJYSnqMW
u42ZP+KheVwE4gBtYH287crubFOxi9bXiMF23Oxo20LvBLWy8KVixRi9RjQpR4oE
y6aGnA99YzjtSnYqfpjoI5BAtaJ4VYEPYSB1Syf2KNB/HWhkBd/4yM4LTD5fKHHB
g3oV6/DnHodtli36h4pUxqJfYsYO4oxOdws66fqUPDSvbScv2mUYa5v4dNu01bhf
YESrX0d9JAwUmYu0GrlfPMW0LzeQOmFn0OL+RptSuPfqsR7XZP3Jt5K7SYzqp8QT
bkzZ9ClzsOSQhgAVUdnQOQO4OCwd/oSrQan6xvTb0AJrKt9Q+fozi40piuZILyDk
EqEN/C1ZyyAr4W+Y8ageqyr+DT0A12DhNn2bchs+Bl3g9vN3U/JeS5gR7+NWJ/Lz
1IdIAWYdYC1sQVOH4xo1skO/6MiU2+a9Y94/ANXiF6xkVIHZXJPbGdwniQx4tk9k
Js1P5onLGPCSEvg65r7dIOCQL1oLwfxUnFUmWn9Sz68mYDXeIS6skfnReagGjJy5
zHUqcBtYOt2WBeyXeb8WzQlxlYtfyATH+pze7k8esj+zCL3oolY/riZkgfyKk55B
/kxHH8gMnnMEhDVrI9HNtqNHHqvVsoLr8FLU5+l0AbLuIC1EC5xqUFMNkmQqw/rS
GbmGF7pmX+HV1ZOQ0scWII7IzKPTpuWRpxEL1LtBuN4ILBO9MSh9dV3ygHpCxdyi
88MjmfOcQ+e9FqgOrqHkteUEHRGqr4mhTFwu7NDK0cZhpfRGEsj1mOrKFHxbYOuB
O3ZmJoCgDzahXbd6VTil+RdNZ98gAY96K0WMZpTe03d4Uk2oAOjTN5NM0So4Qj5Z
w2WwPi49GL7+xWMsfhwHUyABA7eOG17td8MyePwX/lBl0cT4FHwehjWu1KbyPQGy
u6Jt4wQllH4EFcCYiUYixlHc52m160dmefq+wVMOUU7vmsFkFx9nX2I/E5rxhH0z
PYVOSeHWIcB2HAfqQNP9Ale3ZkVO6/OuttOqfPb52/fzvNVtRMJynBzkvafe+WGv
bhzPAjMm9YOpgwCRwPracIls/z/EbOm7JOOtpO+Xkv0fIc66v253nubTGPn5CFp0
tkiL4Ysstz1r2rOmPXkG3wAAYy0y2/xomOlSTAL+Tcidcn85j+NIfDnSWGFCzPdV
oKIalL+xVM3Nv/fpmDdOu4XH+XsIayTsCSA+Xg52rhxxf+8SrFVcCfZZjbIlhErM
hz1MbpWSMeBsNwF82/PyS+nWB9wNiOWToH+ZnDJu0dl9aJEdyOGs25D3P44S10yj
k/p1jyatF9HCvxtD+p9mDnziycHQONTXtw3ICdluFXukTTLZBRh2v7Uv8RNKNwIW
EfvPpLFGc/O1ku7uIuPwk5vIpr82174viyvyug/R778NKRnxFkMXgEsTzj4OEgKO
qVTQI2NmRZphGIPBc2Ou8SuigBQxO9ZIIZo2f9kUn7Pic3+yGcTBuDNlLO+5Xqp+
bEjlYuSkStiGod1fkLLG4dDkZhImHgDCCeByYOMhGlPZ7paF0LsRE9evniCOvZJo
NwMFa6k/ySbKiTQUskEiDtx53igZAWi14l3IqyUCDylyKNdBNWiaYD3IAGp7/Nyx
v/rQDu8Ah6QvhMvUBud7cZLprq42HnjnKGUOoi5PldA/shaWlN3obs206h3XYUGM
Dh/C5tMVl2ylMq+uX+QUm305mr4B87SuYGPXAt2cD+8YMWKLVlpqCVz4e9xGWQZj
Swi4cvTAz61wufhGzUkNgty56BuqC1FYgmuXZhb8Uey1V9HkTb9VJzyYBzRtDySt
pQnri1y2mx37bpKdiGbnGbQ1y16VpV8szoYyXlls81RQWdy+BPTw2UwzGir/L6ZG
x4xfwUOtEPBcqd5z2Khjt+9L2w1VNy35Zl2t7jb8Jy4oUMggR3qrONp2e/yOI5jf
G9IOc+xDFTs/NPQzcE3IfsxvZIjBTPGkQYJ6aipUBk3ExOfwqPENuQSbDDAzJYTd
tqq992ojLXga9UQq2VaSQ51kTyQWZyXAQSQaaIe9i9B7tvHDF/g40QnJEYz/1Nhd
gKBwus4rce12leFg5iJMunp2ivjc/0dRnCGmkYkpg81zO6MkaXY5My451m83Ew0k
rSCdbv7BT4LFkTwaovdCDwspgM+BsFJzkZAX7N1ZwKMv050Ar1jBR1g5jwlRVCr1
dxKexrMBvOLt3yyo70vv9oPYpmYW4CSRBDlFssLBvSKRUi5P4K4Q+Y+XPzFIPHsb
mW1p8L1LXXugKarC/DPNTSgdJJGAQjqyG8VcE/cI+VNzmbqHfnAVcwneDc8tKrVd
nkzv2zOZoSL4zsJEmM5fxt/iWIhQGFdJDa9Q4Rku70Ota0eeKC/NZW2yFY+qZril
4QOXh34j1R+saHGYNygXbc3ZiXFCmbSBT+qvhlavXeEloUQ/MkpRhZ6ps+vmua2P
T5uukQ00e4M/d0zVq9/lqZoPWaGtwKRZggCEDzQd6qLjQktHmphSII/pl1KBfazP
3Mko9oHPajOwX/V8J4LQcwjl6n649W9KBz2pFBkGlG3X2UG4/wYZbdC0e1bfJjd/
BjmWyoxXUZdfiwsgS5wxHuz8LMQsLVk7FlHLngHlf9kdpsaOyliKptcBXNXkLDjy
QAU1GjvY6ymCFcsJLvSozHOIhWpceLlnKe/23Meg75uPNbi6ZUW0d1RlWLEkkOiC
9NtN7Z4CN0H+6duAv2oVeHk5ym7CnU4N2jtc+OmqhCyK9g+nQm9+Eq2Mi2nwmIuy
MDubkXtrA0RUg9nEe7uQc/5Hbkt6xr+K+RxXFuxZObOhgu+xppsqykyAHbGRckJM
DUj8hzVd7cXxTZVEjn/Th6+ZtJ1bixsj/E7tYEZiZ1APfLhFWmTnIKdOhh/UgKOw
7qv+s+E+JgFL9UFwvA4LukZYEY2a6XzX3zGigU8JOczmL2v5K5Np+eCf5Tx7a1lN
ze2MZCNFVyIwVMV/Z6sq+0H+b3GSdAd01FrI6j6egtAa2QO3sTDVvW1vx0Fp0+Bc
+XLtwVfVbPdr4XZL4P+MIgrly4ZlrcMYYtCO0yYRdEtK0TBHywjbDZYJaijEVC3o
KsOpB7HwmzPnv4AdWMv+k6d564c7vyk47XxR2/OaeEXI53Of/tZDJYcvmj72H193
cIthUG8oGm/FBIoINtDhY9xBGNwwIJyjguNFGT8hicHEOVLcMqO/QbIoYa8iWJPX
y98r7xDBhrU2rU9IVFeyy4cxGj8z7ZnQeA+2+Y++n67ATQkv12CqZ7irLn8mIpBi
wmejUAy5pxyLxHnNKBgu4PEoNAXglEiS/S0GBpnH4w47GtDOuYLMptNGbwfaGdF9
OQSCCkkpDO8oceD2FhDnAytYfe3V3iYOWGeeUcCTIKTy3B1LPaZYg3qqmBikQtpo
yBR02QXPR1cTvl3IjkvS6UeFB5/lrfPzCd41xBnbLddrSM9xUXYuyzGMJfmW2cen
Egq+VDzhEoTdcqvfEAV937xsczjui+qZcCrFK7BNL7rb4ZphQFS0jzACEmwDOWUU
NaFCdnQW3L6+moioqwYi1KsUAnq8XNmnXP44h2pDYF4BlO9O1BtxydCmmHXDJH5K
wIsxkluoUrdb/5HaZBstS0pXyVB0vBXeJ+YL7+PAqV3mZjtKjHC0S/vJdHWhcdw0
AijcPQna1XcNYE37YHU9W/2zcQZN7LEQ881GC1R4FV+J/9Ukuc2E2AlvXMKDxSL4
XgSFY1WfzcrABIw3VY5afsSEvs6LtSa3BlQg3LuciO/JXAOD5KgC8flbdtb315JD
K8CujQErwxN/78PBzXWCTJx0RcEMOtddZV4gYhjQT0ar6R92HK9kzWmW0Vk5HFsa
q7ZeFBgj5fh6IpjL3CQ0ec1osth0Sn9OVUI/Glr5DwsQc/PfJ7+cY28eIVaC6Gg3
h+ST1lQHuJICwCAs+2kd2KGsW9XVrxuYbpJ759bSUMHxFWjlFd3zriwkUGi4z/UP
egtoB7KSWCJPC3sIVBxazeTh+/DmnFcIlUYd8ZlobFXwVyKY4b8rEvMIItjgJ4oH
CTqiY3tJ43JaJxL8yuQ4KW69Z6TiZKCbK0tPGlNqCA4U7X9Q6tNyCEy0w3b2g8cE
NPG49svd73vd4r13VMZ+IhCJgUWjnbN2Fpmwztx3Bg3dSV1FQjLO+txUHnIr1lF2
KqDGTGqY/+xLy9G6QgMAJ0L9/2BwV9bMBcp/BKUOSug9BfNmsOj/m80X2Fyi42Al
We6bE5N3bmlNf68ZpyS8O+bN2VZwiHCbH2UWMgZ5meWy0pS8FyUDrnv6cV4L0DjB
nDEDCm1Z7M2WReZfvBpGRiB9N7rIdq9T+ITbXpuZBKkgqLJCI05cIfa5krOo6Biu
ugrIbGZXv5KDV7vxm4nQJo6S0KwrgVqCEZp1HgQOel83b+KZ01TWrgAkFaqLqJSu
mYWyTqCffGvtH1a/V1MOnkyo7RMrZ/MqFQPBda6Ll4NkLqp9f+GkOepxK7yh1GQK
pyWCVd5vKVgi7hKdsLVvFVs4eTX/TroDMaHTKUERnPcoFRqyt9oZqcskyA9xXKEI
rOIobIWVPKSUxde4qt4OTiiYrOhgHh7W6KW4lzsmK+ioB4iHJPbygYjkoOotb9L8
+dVL6jO2mVoRgNvIvxcXLqz5cWx0TKlIvePV56gj0eQ6gtYMojX+HbC/3eRfk/tZ
ajVoPp+5jTiWn3qB0kyMDxn7yw1D8pvGzrff1fhZKi1MxUz0BjFDxlgoQpetXBKd
4km7HrAqEzetdYsMFWnmjxQnp2oFMiWWmuIgbeZUsABgZ869H5JzzogoZ5j/ARuv
A2RwOULxV3eUZVkyXsvDVnPB+GAkA/HE27O+KVtKBHOz7MM1MoG+NnNSg2Dqr7rF
ykwPvrsuCc2riQpeLBPB8jkRI/KiKADvR5eGSYtm8qCnqwJG2rOE1jJpx7dEg6ec
poRXM5hnnpmYUq9NwxkPxQodqsRrqx5G8Vz+JlhFcWqZmpHKOzrf91sSSDuR7tYz
JfNCEMEXCRRaLvY+xrQMSM/3x3ADVTgRjo1k4E8BntFESBJDD8tXuf6F/gB2y7pO
OwVmD6IPHQQOZbvXlV/FXdIev+kpwnXBpF/2RetHF0mjgfjxucbBCiOYR25/IHWA
TlkRR2RxNOJskdUqfYjkgEJPPiVumw8vYIKN31DCqnXuHOu61rf/5uk2Px7joKUk
uGyOGxdSqtjByAHmtDarx9Cr1NuFbJykWAKzqhmCl3gJmFzhQG/M+kI0KLJyWHCr
Gjn1/KhV2Fsm7Y9mE03yIphUpoQFQxl1hkhC826YbfuF4LOLSY5KFqfQnA3cl9L/
glEyQNGFTEnrVT/vaFSjYWoooQuKW+egjAJnErips0i8x0zp0nxzbdOWUWldBn4b
HgNpEPjFDeiUcysf2VNo0HIwG/CxnB5jHRv0BjEDkMbqkhXP+lEIZwDZYarcZ1Uf
TbLi7cR+cpXDJsFGUrC4rhY7YVMco2JalwSk5vTMtaFjQTYF2Z9jyviHOELxg4C7
faaN0/T+fxXBr1+jfOEAkzMpypW73cxPps+0OkjYO4ow/JlbC66NIOdARFc+EXWx
jnDF7LGFRtjCNqKVJkSSpBFOj+nbQafwZV+bVDFfb699YgdRgs1hcGvilJsyM5bi
g20Umj51tgmm/Iw0OoWhwqFFZAhs+nkaf8Bc/SLXUBz7pPML8uCWdKJBeAQG4ABK
C2reqtFM4BkWIJB26Uj2/YeES4uvS5lLJCnircfoMX+2Rlp9P/UQaBwq7R0K0ZWj
hDjZEbfjSVfpU6c33xRLBrAWgRC2kStGwKoM9K9b/C6G/9tSky5lKBFWJIBQ8UyU
kLYQJE3FcTVraNoiEf88toML+i5HJWGYoCe0GbPn38I9cTICxVmIz6RXGph938ak
gnFZd8R0yVhINhCi/yT/GDtpzF+U6QVxwPC5sbUSHSeoDhpkppqynCrCEspDbVMT
/CBPoMdFBTK2RHPSR1R3yQkwe3x2n7zcrSTxe5ENoXogxV3HaAAmgWIvLlxHk6G/
kyTDIrnJBXQbrxJvPj96SRQlWzwif6Wb/M65j/Fs8YeZP8nPVBl/aYA2wciO8+Cv
IPIaGBqHaJllHVAGxOpKsXh7pDR7XM8wAVKQ8E1JhrZus8UcNpmSXktF2JVPctgw
IeoqfRP9hJkYWWIPvSrgrYzUfjG6G9vwiNGe/wGJ3F4I1jpmyITIdcn4Nc98pl8E
VugdNrO7+D6nUEXOOeYeRW0UNy08KzKHviOCj1m4C1sgBwArl58majiIYQhOw6Uk
2S5RlzPMOMJ4INwYXeVtgUM2EnFFtU9iMzpQVmmdZRSWNaQaZl+z4sKWXl4hmjDe
UTrM2Z4hjhG20NHvLQFRI4nRpCd5XjOmpv369BqrR9fcCNAq2YSb0OH0CD6tl8xN
cO8NLI+cyuY7RrAyAlZ8NQPiBjOmWIKqkFDxjtNpPZKiGCrpgt6Hi3seCQ77jluC
TBgGEbtSrY7ZALgQjC/Fcu0hl726Za3lYmjBbKyCE5gUrietgurLgYMswf5nakbN
f/hiUagl9ly+isfjKvHb7ZuD+RDuqkyoyUXB+hO4bej0x5YSfJ7gQT118F/Y4YTL
7JIWhZ+KjbBEN1N2+jpjx89HTee9AUCeP39np9a6AsdcX1gR5vP+WnPPyjBj5hzu
dTxhTGV4JVtYbG9zjNEgejybUaFxftY/FAnatogZNhlaWKIw2FQkwxebmYo6BJoX
3mvvIo8N/HYfVovXELyQ3u/+RksDzd2/sI8lLFJFTybNBO4USiRadCPX35RfJckg
VAVcDlqG2sARAhvxZyVZv12Y/UxY7IgwbrPm0ooZ5zrvOeNgAlkIpur2eBKyHmyI
Q3nSQ77ylV2ahtRe814gjstHI44XqaTRxqYC+mYMbmlqhYwyi3EUaXDCVVbJhmLc
xmZpt1OQAwYhD4xa0Gbt0fy48bp9Jw3hVdpk/DyezW/7vWBq5mG471eFS/YWblPV
E8VwhbyBHVhuOh0/yDWb8EbfzbYcY6LWQlK0RBxse/Yvpr+XRinNI0EM+YTFlBqR
Zs5vT5bXirvWgOXPf8BTReR7cMPDZttVl0vV0UbesY/HePg6nF8HcRiJGXpdfuee
6b1t5fS9s4Tnol9iCAdpvGosCxcqp7Ds/+W1U25zZlMPjY8qF+7G9Jipe16+dOKV
6dd/DyXO0KU2vH8IXxeodu6BDbe3EqL0JxmAARUPteirdPvOQd7kYH2cUcASJ+qg
2GR7mK+YdimILMuMtXsn72shS5fZFd1xX3p7hATrHCOo3ThmJ9ysHRy3ix7Z7J6O
VMbNA2vI65AMsqCq3vl9/SYb7X0Z3KE1B3758gWaEbowaMxF11hRYu/Y7T3pM4t5
y9RBC9nJMI+gLpaB1No0OXr8199FYhgQpjAvh3CySuHlkFTcN+EyMP7/9aUiCQhw
2IYSVgbPUvsdU/lKxn0TdW6dU98L9M1d8PgMH5wdDftU9vk75pmOEhihoCywMwmc
eOMbY0STgIKDyp2HRUKDYqMrXgy6V72zR+H6TeydCrIfkWHyGp7VQEwOzZvvKQ7Z
V9yNLKMzuI7cBC4/S1/fAA/SqAVli6mI+8aQJ9BNl5kyfy+kA11QrEclX3BIivHt
EgAjWUgBoigX6j1/GMPhVTNJP15Ym2+3b9TlJo7PSlypfOQr0AprKdvMOicVAoMy
ePFJZB4lKOgfMOzzNVw2SntVgr2SFNG02hKBIiFxdfqMC5Wl7ZaplUcfLuONaL9z
ONeHjn+JEjgf74XII6XSjIqUSgy+KUIHQlWATn5GYyez1CjdL3HXjDpSYh1adQfx
6+NhomjANf3LRiDQjV7NUrg53Mns8ag8P/2tPUniQDPXRy4K9r0MjB5p973NvsHU
dIflkAkXkxZBj5e/VodCjIFHeunMiPPtypXRx+IVnb3TiIxN75aXmchLTEqdaDQU
EFst6pMtbCXlZboux6MgcZKOetRnXnx3jxJkrfqQ761S8o4HHEWzMv1V/Xr3I6Bp
3ufB8zQ2LeADkIoXFFr244tT581fRa6UtagpGO2faMJy7iC922CL1qtSV8Wtphe6
Kbzswc8O8xkVVFHrcnVxSBd+bGaI/3oyA2Up+QOv1eRaJ4aiNlSr2qfVn/2V/SXp
Te/Cp7vA4ZV4yGLUnMI14xjzGXEPOo+1/eD3kpcOs7UnD+1P62O+ZwqMNXUMQWQS
zFeoMxKQuRbaSy4t2yCbQxZ82BE5QQtdY6s7vkXA+tQobbtTrf+7yZaKutbQh58m
Fc7e6AYNfNYc7P20n0pKrKhRdDIpkp5eSI9kUQOsFh6uKlxXQSxvcrva855eNPQI
e5ROikPhlJpvfW0M6NQN2eo52MT1iedNY2BV52wTqY1FgFnUrkwexvczUpHeVxcH
TqBKibuVJc5j5wXzGBVVtDZ5QFj9dZW/27TPsGVRd5QXmwgIUXqXG5ksdHvObXGw
9evpYnsBsz918y2JLMvMF9mfsdWNEPNkH2+evJFv6aqIuyHSPIx7UdVIX0nl/nJl
js2BnZZHYFz5FHVd9m/zvoqc6t8r8VfZVTHUKnu0LEZLIhEh7UnIK2YCo5FAfU3c
Mm+LQCR3nBm2twz3Q27n+Z3zKkxkK00WqTWjppk8PRrUT3gxwlc/T35NhsmStU3q
MAiheXvI9j2aH+yhVSdhDpce5sUmw0sO2SZBMolM0HzJQJ/UtWBLDKJMW9s7KBNI
xdtsr7dAyTBaSOOTdYUdFJCLSkqEj5rkjIBEaYDAdZWvfLAWHwq+V+jT196GiHXh
tTFlqki7H7PfQuin5p1yFb9kEVnATasa95GLw2+F8Lpt6+MLWt+ZS01NJ3n+bxR0
HpeQnPG2wECX8N+Sh2MoVPzC7pQI1B4yIiLz38erHGOGlMifQhrGmOPIXi4a5np4
O856WYE19d8h00hMrMr0YsavU7kiLRORB/90W0vY9uk1FBNMotUOmq6U/dTapyWo
TAHXkeXphUyhpG10UWatY87gD0SNtUChceJQnDSziFRYPGc8feA7gkQFQEqptme3
svH+QrMk4vCtnDiBOdqgBum3Au+dkYCcxraZDNxb/zRJfsjxt3ENnl1vq16XlsOG
d/9jUUl23pTLSXmBRwLz/sUAHZlkO9GHuk/mxjF60cZFgYPa6xXA9ZyarJF4w/ef
PLfIOpl2FxzWjqYk3ZxoDJUC1qm+6BSjEAw/ZRnHZY9SHA5M4IjWIp9EFRrA9j+/
ewF0yCnh1Hz/HKoHg8jnzn5c97Yc6bZj3cSMwlnuqZwmLhdZqdcp0YeiO3h6JisV
lEBTi8IbljLudFL+ttq2/bbSScKyru8gZogj06Zx2P006cqLezGu3xLbveeyVnvp
B2jX+88Y/sg5OWMNqzA7+/FOw27ap6md5kLmEk67kCa/NgllPUYkBfvLyQ1np8gV
USPgx4pWBE0zda2EgjEnmFxBpFi1kjQP1Ruz462qs1KoYI5pndcRYtRQNJGpw/lw
hlrtnNJSsXU29bw6eYTX78iFp6oFtHEsoVVUyUQ7RbmdEa6q8F8G8ShDwh1ny1Gz
gqEJo6vl/TbbBICUIR+K4lo9OjdU1Ju31jDssy29n8jmqon+ffqyAk4KpCJ9Kv0H
N1WwxH2qTkdcQLDt+XEE5oolmop9xiKYoXotWprjGwx/IuZAW/aretKzXqA4hw0h
IqMlgJDbVodJiKJHNu96nkU2nZCF7a0p6D03UjLVj4Yd/skoDr3/amPwsU1VvgPP
ZCSJIagzLRntbGRkGzlXSLgBeH3QuQzIDrPEK25OhCpmktunfbasj2IxnuGIwd3L
n0hnVRocX7+g7GYU7UyDJZWDAGaJtPLQz5o9v9sC6dPoq87pFv3AQjUqisXkfHNs
49FuRCXNAREoCy96Dr3mjWTLmKLNAMOVGyeGQWBnm8tckqFG8sGjOF5xr8oNyHfi
H9cQIm+Xug+g3BLjfC3ZjJW/ehhH9yqk/ofkxieRbYqhDihR6O7spLqGcmv/KVaW
/x85dKbU0gprZt7dG1yaOiVrpzYYG+C46Q8h/7bJsGVT8ivYqnzZoWOKF3JuzKZZ
h5RbN9wz0qfYZKvhUTG7SOcaCjCTRq3mnfDV/qHnuhUgNqaPmoJBzc/jWDmhcRIN
8MNlc/BdIAUdYKQStfexRlThq04JZUoa+abvXBK6nmwHYJG9zyE5bsU7fERjJxEp
Qj58RHqhmXuyG5nRjbY3ICnRRo6undp1Hrev2JafUoFOtn9a2xsJyQJNml/0MMH3
yVGMWOeFkSycq//B0bx0Kk/X6M1bewUmeNES3iytUeQVYeiCvxqyqu8U3Y8+RbhP
P3IPNMzocGYHckDWqmXoiLbum3cRYh8fZYAul4gSA6F+rkYmDEyepGjYqdTpwy/8
DY4oPvpTLRbXHRRtH3gvmlOaXiz3a0BKSAZswiJFeHH9lax93HJlBcYcocp3/WwJ
7lO/HkNcnMFXxA/yfqpi5WmrGe0JCFPfDQ8rDnidbjxEak2uwge9iwXkxaLaIfog
8hBf18/FqBSpcjjVuwFeOePnrmZx3LdQ0e1an5+yDfRtau3F90W+q2BdqSLPDSvW
bC+uh3Sd83UjL+Ld5y3/Qg1Kd9TPojghI4kApMMZscWkhrLuLCNtBBx8mX/b59cJ
ZBIHcwSj/NdFhLzWYuGPKJaYdZPzl3NdfbJYUJW+HauVDOBxCV+rPRovOEUt9Fpq
IEmxoApWmpaFWQ90LG0DeqPC+FU6e2pyTnNFszc0R72fSAExVq1lvusLnRo85+11
0FxkoFMzzrlzouc6MkMUudJFqKuvBcpyDITQ+o48n/aGW2ifW4wiACukiX4CmmEk
Bgswud5ww0hqmlcEAvMKyz4Wo4JuwGTP5MFm93IQysrToN7fuFOQ0ZCHeEX+c4hb
N/5xUBOzg5WrCfn9TL1ZrFBsJGeMmGBBbf13nyQXi13iT0ks89K8SMywpmRSkSGI
oXxiKOtI444KP7Eksn2yYAlJZpUlpG6VnTds/tjmvCfbB3N5f3Iad3MLF/NUp6qT
uZM+uR7DHmTc64su3juvFuKueXTsHpcvaA6prs1hM1sL+6Msp9VrZPvQ66hFZ0ON
NX8FcjKskuvyEBU1DOBwcagH9lWef2+EtbK6bL3YQ6z66XadKVPOtMEV1bBTPHZF
MuA1icf/KAVmCcIufkkH0HkQuniPUmhoTTjCBMvy5FfhjuOi80vWiiBm7CdMJGtn
i3+up2CPNF5VqOjV9D6K74Q5BqBBCrcK600gIRNzRu0IHge2B5yoyCKJrl/0XgN9
5OZWXDCJst5wor6dbi+Yf+xqSHpI7f2e8rwdo7itbX2esqPy8baQTLGDWfUgDWhg
BMxLUZ1QgGIt8J6UHaXcOkKI6Jb/2Vru4SLHlBaPzcI7jYq3+StTT4jg444AjD2S
EDscPx1qdfeWaVUNKNapbWc8AJ9auZ8v555SsqBnVAnKAKg+NhkbDJag0102VSSy
vfocuiXPYijJmMMiDOF8fFD16uYZchfQ8RhmlXl/etVkqzsVBuvEWWidhSolAscK
Orv+Lmq1/0GlKZWwi8sAdqUlsW38XxuVFXgjlIyqO07wZuyAcYZNF8SpNJGajzq9
hFaSF5pO6LMEcqJMI6kBo7LvrUYomStRig3Y3J4IU1VBPB+K+C2ltmQPYpOp0Fb3
Wa+Yizt2X1QFaVRWvM647LsM3su34P8+A83GvCjkMhNi7xB61BWjSiw4qQbKdm/4
mLkJViZQe5zRXua24kmeFa9xsrLsfEhFbiuKYqHv+ciyywAXFyw2aan3cw1wKCj5
wgMGCNkpBGwukc/XSPp/HvtORN9WbjVT5wY6ZAkW+qTkw0GA8X375prbk5ZjdeEv
R2JecIqnBES+9lb96XVtGFFrlZfIVs21Q8uK4X3GjW96+nQU9fzHfru4qEb1Jrd+
hZDsbU1S4nCGK/IN0pR06KcD/10tB+bq4WUWxnj+PFAbeYSgBY4VFjITd/ddI3td
+IbIwYbNW2RG7oFZ6dXpIlqhFb0BqGqCDV+RpUy8uQxHNII68+x8ulYfs9jzw5zd
KBAf78Nk+MhEzfeMuU9eQF42q0HneawQaQnFIAQsJ1PS5O3W+O2yvRmRfhL6cCKt
ns0vU52DOVsJAMDNG/VmFuVazL67453A7/QJ4Opp3a86OyxWeKshjhiJp6irU5cC
AekPNCFmil8GpqWAzpyohJB3cHDPJ81m9bySPSv7EmDNg1bjeVd3TSnS1rIIVY1I
Q4yFa4BY22sTAVtxeSGWNXyhpBn5+BooF+GxKIy0qcYOAm8TUhKwm5SNHpYQ7LOp
wEP0aK4BI/k/qyc9hhVqdQE1NaCYQWCuSpbQszj4e+GMYhYDSa79UeX4Q7ftx6Gd
TVl9SrxfSMrR8knY9gKDFdeUpMQskwYtmD3kqYY4JpkgZYjKMmSFhbYMBVa2h6fz
4giRuRlxtpwUyVoid159i/rWYQpBgbR8tXdF9b+q4OOaju2Bdq4XRExfOzX5DKoR
C11dYaGWp9anhCJvBY2p86sefqeEPrAWtp36qdYlOBq4qrE/7dkDurJBq9wmoznO
xmMvPQM1/fOJW0keJKjEGPSL0B1b7Z0eeP6RpDbmoO/9xZSwbQ35JsEF46h+2W2t
KTB/ToPhXU12oA8btFI1EV2df38E/lFqRf5vzy6YYUi+ElzoAoJ+HbUJMgjlHVKy
7W7gdUf+Z0THTzaxBfBvrHQLEIMSe94FaHPBioR0TB7ky43i/vl2QcAmvigajwWa
5aL72mePRk8ntfFeQvj0Wr/8DownEwFgDgnZQdT9m0W8jbKo6H9X5aEnehrrjibY
kzbrxDFeITlHrGEqDUhpPKzoWmEvrXtCWBuWW9DfNrRZxR7NOMd15j+8wN7giDV+
X5fHQpv+jvdnV1q5wyKd+bfCi7VvpK5/jujYAllFdR9Xmu7oG1O+BSVfZMGMpcsV
G6P/zBHipjknSzUlntQSIM4yQnPfEftCcX5DorKfS4W21wNO4ifH0N+EMnhVyX9S
ZnrunBsT+QNmODLf7Mot/RPxIQfN3GrsCRekfnG84K28UD4d8j8tIKzA6Jltu1nV
SOjGgjj/3rIPtP4+sC1WJ/AhG6QOW4vEUIiMxu+nmlvPNuPbHcJrxFVW/ncavuae
D9jqcd4Rk/+o6632XpGV2SLa/Z/B5cwcfemZ+c2xE9L42W3aJr6Fe/VZm7hhe8uH
47V7CUAl4n5WBgz4+Wp7fSbSq2QIzdbU511Ki/w4nSXX5jFDSww9Q142WE7dUrFf
2J7lhN2MoKyjKHRDTjeV4U8i1BbN6cjRNtRBdLiW627LboW0ACRxDRduYYtxGTOz
OkWZmMjSuxapCyydbRXlfyvDGC8tALw7VBIBamPyhkRY7eB8ZhOx6KVx8PtMSKf0
LARKJAnNBGpnDyCUhSaLukgane0J3aZc3Z/Zw9aOmMIwPo0nN1VFDffL0g0VKvkL
Y9p4J6c/gRE2/tSRWFu6SrU3Q/fjB31kfASgMmLNFvwJ8vNxeifETnbChUeyL3jT
bng76fDYlTxo/sP4qPByko57i+MYYdZ30bXiYyczy3gNWE1FadHXtBU/+2CwTVUa
FP4MP+SS3WDkcEccpHSJJDcrvmlR7ZSqqh/5ywCTSsxJMxW8gCFKuutKVFV5ZcbZ
Y4pEcuWQBlm3RLRsQSjpIyfjAwtNn7J/f+TVMK7dqxpsHOGAflFxkyU1S5RFN3GM
Hu6ELk9/uqqDnOTvPK4xyIoDzwXi8xxxHQuoxOFfy2ODe6KxupXBEpA/94Jrub3S
M7O70CDWfYe15vfxZEcork4gKNP8y0uY5gIPOT3wocALrYRlyVt1TPS0Ce6+85xq
sNvYHEryEEh8VOx3yCk8/h5dwp5ygPOMVZRXTvgaFZQtE4hHODo9zwPs5s/RHo1D
AZKG6EO+fljfftjtIJH6OCwNve/KTs1k3Je9j2SZIVLJ+KOsQg3rTHBsKof+wLE+
5QoSBAX19awEUt/LS9KfKC2hp8/v0B5VW3L1PqOboMDvR0HUqkeScSE1SS/GqraK
dyiPs0Oot77zkxTnY2ZCV85E8lM2vHI/zyzJrouiNWYnMMWPzKSVA0H53JTqw2Qb
8S7HzHWHvpQ2Jw/E0w9PeuCuRt38UNmkYM0kzTb4MtbGW/UhYao3WbJ2liXT1hMj
ioEa5+8MX9cjV1lVkveL2G+rOIoB+ZWmXAiFrhdl7c4WZzA+JfJ688aSLe5n3MU9
VNXE/QzJJ9zjwMUYSAKT6+oBFEV57RHqqvhphhYi/dxW3MczEl+LZNgauQf3XdqX
I11VaoW4CsssJkF9dGQXequcWSEgo+OOxnvFgRnjtOkKellUILhs7bZkdDbAawO8
768gkVPL60CcGBpNuBsxBXsNktIwRIOZjXwzpW5v2JHUOP8z+TuiUC01dGY8r1Zz
zBsLK/XBf9nZHcoOJokd1kwwTQzd3ZZPm4gggMXLLYWZodcMQDWeNZ+C2HDswoDW
SQ3VymJllbV39eRSu6ZvuJppS+KZwy8tYywRxdeBEOKyRLvLZ5dWDCwBecwDGHXT
tPxFVOr7Le3JbBrok9jXJRbjNUSbgg6LFLWRDWFKsaMm8oms81CmMnlhYVYsHZJr
Q3goOXydSQwa7DFHECKysGrhh3TY2H3N9SNxtnS9yk7VGCFya9YMIrmWJaij3n4G
2hS5CI/p2twHd9hDsBZzV7StsjEmSpmxN552PqLV7TyAJNMMfzKXLydj4cpA6Lvj
ikwWl2xe/raM7/dO2/M6Bao/W9CV8dgvYCi8xHLlY143yngCoNqj2Q5dGaDmygT0
6sPSviS/9bqpfuJfA2I1dTVemG7qMZdhRiB2uB8e29Hl5IQUiDOp+dI7C+7aYXPa
HHp9nN7PghC+xCgLc30U0Y1qrGsFdBudjnvNrkABfKZJpPdEjHSjEokg6OPoGtWw
AIH3WGUCaqoA3/tFdtWEe9C2ax7yksbGN9rpLngnE4a/aM9vYM5o/rxkRchXovLt
XhZZ1gBp53OC7W5uWcQwMzJWLwv1pa0dW7ZX8xvhcN1RXa36Gs+1b6gL1Xx5Zy9R
m0PhN8VEOKE+2zNJutTCVKF+/Az59DNsDi7h0IGXi0KqV1Z55d8Cax9KgTAGKwbL
BgbvggaIbzOx0hjhiuzYCdQMCpiG6CFhSe2EeCRNQVZ2wcSz4Wk18SGxwDB0HQ8K
t2W4PyqInLtPrLDkBT98pq/dIxdG9Ple9q0O4BprUMO+PjRtt/pw8c2H2yQBpx+r
Nu5uDEKy0Hv3CWZpbWvJeP9L//F/ptXaDIbMC2wOIEE93vFVCnFt+gYg0x/EH8j5
YjMCqiTXGdmWRwsE7n6EPFmnHekzapndbSni7ERcIZYUAe7+Ecoa1ibP8535rcIW
kiJ+7JhmmYNwQfXwWF1tkJDrbnSY0lW+kS7K7dF7oUy/TZe3yzukQ+PrxA1sznXD
7kSaIDu6Eq1dJpnWCneEFaAPzajyoP7FvZ2hPOQfddjQ3MS1il0C0WIC1NfhbsSk
sOFTfmuYrSpB8gZC1CuBI76uiQ0FRJGYxUBQpkQmU0DpsM7Vx4rP3dRgvYnk2rOZ
Lj6jdA7RvwdknYelgZF+PKJe6hOzg0kivUtCyqJrRiorGgdvYxTdpWfkqy7rfzUh
u9Rn/prBqXBf2cPOdj3CxVXsGb+NYYV+hwOY0oMi/9nMNFTCFcvMVtPw2crN+CaN
XGV5F2f0xeASqBF1gUx+szUuuyTRkL+vB7BJGn29tJ5GGTZgh6mTMjBWTd7lXSma
r+rGF0L2Zh46jTQVDnBDqMcQ1L1SXIhzfHqx3fUXegkQYs57R+45PMA8nuSyOZ14
cTNiyB0MufiNx+dApwxYgC3KgP4oxhkJHafmzB8+rWkTzJFvV7AtufJEns6miX83
oYgUkFGhXQrJWKCzlkviCEVNBgzTZI5MvHHV4CMh8lQhbPT8AAVcng1bVXwjzGZp
BS64oRe96uL2eSLA8QGRX237fL+/VklOMkUCs7tRyeU9+ejmHQrqYe8buWeeNhoe
lbDyTbAq51/I2FUOqD+z1FLNdSCrfbFdTFZV6R7eVBJL43r9hNFlLQipBl0c+tAK
aBu5U0lvBcUjBfAqwFMZDIxJmqA3gEK4O3tg0SXohbMFGo82jnn6G0q77zfU6dLn
bBMHJAlDyZh/AdAO25AR+S2feVnAqMAE5MHRpCy6DqANHp0Tii2fOc7xi2NR+3ho
ZN21jRyjcu/4+3TbM6Bw/YiDzf2wDFJTttAO77zLaYlRoWcmlMRZafRRbRIKwd2F
9BebqG//Rb94Ein9VmMmgn379mqt1kMas3nbZWrxwqLvhvXXhWGXUusacbINeklj
/wkXUxYWvokldxg+TxovaLc/TBU5UqicS+4xs80lraoP3hkE8dG6aAA0ItagPiQE
oIO4ghhVGKDpTlnU1ZxsHWlQJBPw8oIFp5/9WQnaSV3erVXtA/FsCt3n/qe/+apn
jsZTTlHEaWjGNP+/fL8DQq1ah5WFdcPg4xx0RRQbGRN6RkWHIOK+QDBHxNJkHTxn
YW1khMdzXI3YpUYJf8wrsiUE07oC8x93+pcXMs4dsv69K3KkcbEtmkX1mN/0A5Kj
7eX4gnTcGLwcX4nhz8V+987S4LmKTCwUPg09gjujfFGiVSaH04TiSGyzbq7QAI3p
bZatVuYsbhTpr32zCLJpeRYg+UUjgoP+5ooi0MUahRdIJr3Qt7jCqm5qPoNV3D8a
LQY6dzwrko5NfvRZBcNk0iGzjMo2uhdfKwdm6Y3mLsjMBMQwuSrLsA08MU4SvyrG
A//BppU0R3JXtYEKRdw+MeEql4ht19PeN9mizsVIptub0utv3HHIs2od+DzxYVbC
ug7aK8L1KcBskP5P/yASC57XpeEgIs1aZj6VUrn3vLIXkV0CjtjUkjBxl3x0T+px
7+biX7QSC5Lue3A4CWIpRXqgn8wLvNYqdUeIF1xQaf8tMuhfgUEz4gCQgmRlmeE1
tgPtcJFVk+1NZ8P1Vezr02g/6tZdKtdH5TZs0HROtoOYW1cnhjrGkkGdt2squotf
BF98ogMX0IBWGZifqz8KvbjP4TEB1QsQJ9AallfCSiNxX9io5pgB2Iv4UwmotSDk
Kxy+H/Dha+KhIxOOZty2zMbueEDMkwwB/Dp7Y+QH/+kMiYsuicdu9Lt+SF7/c++z
Ur17vBkB+Q8SKMV17WmCS2WPHZGvSeAfsER66wmwFzxjApVZPnbsGajJ8z+n5ZXb
p58l1rGUmaaZPrLix6aswORwsgWPPIoq/MDU7Lfoor59dsE94QEXIToDHqASic4Z
xbIO5m137051PQ1BERp6jFwtGS4c1SYZ9G5EO4w1ER0QHy9BJIPrYwY/bONDVM2W
Sau+Z1W9J5JWTBuT4q8ElILBhjP1vwwJrCYhwI7sMhmh/b3xxYpgcHQAmx8wBpmF
gUXBeR5XGcLX96sCQdUe0itZxo8T+pGs76xFcmBpUXuDwdxASEzUqHYyJo3yr0Ns
joOhhaFQVm8ixXuBIr++FN8PH51dEjiIcySX2HAGMrJzOyDIHkCaMHyrwXGV6k0v
DorNBeWaSCqpIoo8bZdmh48rwE4+4ymMr2LbQUe/S7gXh+0PrFjxOFc4AOQKmnUp
g8IMMtQLi0NkmVd2rnj+veA8LA7I4/x8EsjbKjS0skYyVY//rRfXyC4K4SixTe9m
uMyt7Pl1tKJ/cZPDYNS9PRgExqMc1MroF4GrwTRK5NG+YoMlHOrApK2PIKNAc3f4
V3yqGoYscGrBLOHorENpgNxxR5i/z8QsuIf3kNgmXAAevEDhJLmAUMIdZpps4wCU
VwBmIlE96293bjsrwy1pu6MK7ZwiZMXV1OXjQCEH3/S7ms24/WjiQxCJkvN/YioW
KJpQHir6i1b4jp+svwv5L+M3+0Ih2lDS6BY34l+FzZXsnaZnNRwdubrBtqnzJyfl
bSLNH0xr/p+hDAO0dXyqDiuadu8DByn0S/fw2gosFn1ufMrb+iTRKTLJ3GyXznsA
B8+w0Pzu7KgeYiES9UHYPzAFNN+/yptTZpyFiwI6TSwnfO1Q04N4m8ko019R9YkC
8dtnTdOmVbPh/mCFFFcGvvIuDzUiIZbmN7YoFLR41oGqvl1BRTTHOwPfiB9yBK2k
7ndz63/Mt4y+WvFM6QGl/7PpZhCsmatELqa2nZTTs7fKyk92+nXKfnPs3v6oh4Pr
0O4aaBAoQOSmBivy64bbMM+ERWIaDznoVtM/YJgTi8NsBt0r4zrL/hXJhfeP5ED7
KdseYhYZMc4MvBVDSttuZRDTqpKuguF5t9D982qpSDApCc2TAPsLEVmvA1SSnpI0
q6YqA7m/AyUfKK1GPbYQWhmeL+LpL4WaIvJvSeIIrMV4HfIkxCyAGTsFb68f+n2T
orOJyhVb2R0OA1BdVNzH9tyvtZxKn820DPF/c2OOKQJyK2RlqTOUcrcPtBjowN7C
sUANxNYBTMqG4pGi+U6hi0mpCCODoh2FdU68/2pI6UPsA6NvrjZoy1R/4YkjjAtY
OiazQqjnnh2Fuh5fz/n90ZPSBm7eo1AYNAaYuTAPIXk+wDp1rPo+unClkxJ7Uhj8
EzNhWnOL/KZ5RlDQBg9LUh+dzOijrDCltizdrwkRIVnOdgikV7ktEjkrj4BJ506r
0WfKC9fggErIjfcbF8wSY0LE+IY+bpjkmDpvdRRABaYryZpdtXha7y5xv5SEDgMc
ehjLAL7bYJ5D/t7S/Y1x/zbFYayGk942kybCNBuNSzu2WF/HtpMWcGXGalZhuoS8
1Sc3fu4UvMpFS3kbtCe8zikXWeY+usPOxi1PNV7UNTtlM/TwEJFnWRHIcHHAZtUT
/Mx10bEcrOJDmK0+12/BTmzL85ocXjcVa/0HN9ViZC5l7jKmvLPqIakINgK1foig
VWcnCb+GD7Kr316W9SC86hkra5+sVpdenSjlBUVZD6O9K+3hGohdpF9atqCalpY0
6Wakuri4yAGiidRNXPnjsJkNq3/hcYKNk86frCDQ5HnmfbaIBkNwRFXa+zAHHX4k
+oO4/lQvbZ3SAmxKlARd3NaCB2wCi5M5I6quskUiTzvezaYu92z3fpu7qYctYlu6
7Q7WJj3rRjej2xK7e6ZerHaFMsVsIxPwD1gKf3yuhFbmTuNnnA7CcAsvyOgnxUcu
NNainOqeVLc5hJBypdzahxxTBtBeDkLjr2KH653nnlRv9Mm6jz27IO3ykRaFTbbz
pHhH1CfINUwte6xKhA3FE3+xDO/bcbGkEfDm2vFBWXv23r5zp+kFvZopYTjj8cNz
oaRpMcsbh38DlShnmgmTDcDbTyvlp/ERWE866K0kjIduJWdDpiI1kPwwxjz9ythQ
jBu0hwlyOTyNiqZoRe/TZHIJo4i/XjXWaqpEgW4Eg9bbTLBVtEHu/0zV64kjbTt3
GxGg690vtkiGEcCzSPCyyHfv7UGs7K4Gu4hS0xlC5DpNzo8g3oq9tijORHTujaMf
zeAiIUFgEfyz/xddYgtH1U6reEEwnXXkU62ESRyx7L6GQQ1NxaYj+bWY+lLQgpfQ
3qm4bP2939KmzBBg7//4+147MpgDSWzjJDQCzIbi9OCqZNPwIp6qJVD/Pfd+8wAG
F2uh5uOYkMXvPxy5ritKDDxV5Mbja67vuPeFgPnRYN84DARn+bgNFKn8hH622teF
j4qJF0O07YU2eQ+m9zdFE3nGT/yTTUKSgtKV7Oh+MAKiCTtqtycVfAHC9A3Ei025
ig75OrnZ1shVGdbyNsctiLhfTlqB6mqbVjq3wLkkU9gWoZj35Vnc47XSjAb9KFEq
8rMex8b0lkfcZtyLKMofL7YR7WXNRhDcqFb7Y+TcIQIKOkhXa+VTGI6lC9GzAw8q
bOvJUNWoCCpA5THhg782FHshTRKe/K8liZfO+ByBqEl8OPyXAypOcUsgnznmUiFz
370eePNecqot/3ovoS9YFBo3o5AW8VKYniV7wJCofPCocMCIYGVk56T8iVPRuKyD
pFpe2egOzcN2KiWGTUKPJAKp+i680Ur4cK6DcNYaASgTLlz0+X+bfpX2pGrJufX5
5ohCPG8EBHYwR5o5anyDZbPABDNMUZ7q5YPYbD2lotQ4mUoEYhimOGApC53qxxl0
FvoZINSC70zM1bwF4D2RqsaYELV/7O8LAQzv8QBn4d/xHOS7RLQHjRQXkK8Vs70u
v9N/8TjEXUvI6BJgYSWOypb2KBeyrJSRloZbTqQwFW9cVIQ0KtMCA/9kj7vLLkdf
T98FGbLad9Vf3UCiqlnRxIdVgH7L4uLhpHwaaydmmyWCDI7CDlzXM9uNGNx+lop2
yCGF4sA/jTI8dqsmOUjzfoJmAfkZvoRHCSs3YtycDGAOhZu+h8t2pp1F/IkVP6Mm
0KNgC6hOHIBJ2QW7npvxKCJMI5ji/CSsGvkMUOTHgqgjyD+SEPTjFNX2w0BNLmUC
8C6qkFhKCP+XV1U0P/V0+5Clz65zuoD6UxQqUdGnP955hl7IDenWrbV4nRuZOctV
juobDQi1NMHzqo0Ahjw7QDK+92W7HzOzyVp/5WjqBDOtML0uJDy6xadCwpLKGu9e
drkrew3k8vUkgDoUKSdq5bRo8Z0yfMo3CSgeLH9DjywC4aOloTL/W/aiq1LSQ61X
Dl7Qu4scd7vUgg84ztdcDp5wb3or7j0fGBS+yMdxj+uu1fBoJC3KAPBjv+bQx2qq
iey+aDb1w7bArkpEpgID6ssIU4O11xhFdnywiYp4lqWL6zvyYmLTfALlBbSQr/Ig
jts1Bq15kUik4kVGe86rB8u3j7FM1m0F/z0USLYfc/x7TxUuEs41oNqtnz7pSNjo
0fuDhKk9TUv94k7kB7IJhFqWXOxjxlR4qSPM5P4zn8ckRc3BOoNJJ6VouOjkBppg
A1NZwEPIlIsWTr5DqbtjbYyny1mm4mZ5JdczWKeukX+SlVn4LtBL9jEj+It00lnd
DSS+q34HV9KiuKYu7pXVse814PKDZQIG7AXs812K7uxJjG1+musnRTUi75m9/t1J
enTwDf25mTQsm1avBI6XG82RvNf7dbwKQPOWfN/KB6i3Ke5nJUPv3uGFA+mBs4RW
cJeD33jckENw3EuAP5tV2qfgCLN8b+3V80sB8bhbTgwy2AA/jeO12WR5ZijaIgrB
4kcv+Kf++6Qw1sFiKRQrD1YE+C3Kn37SyKQeQnVBvUIuUeimISjI0oG+oRSerkzH
taF8eB3mhb7QawXiRe4VPrPPSQatmZW2EFmLVrpY8jzdlMdoPSMSv8PTyw3SLq7Y
mFQwDlExFDN+yDySiVmA5WdHGAZ0QYkKsvntQlTstSqBTXkLDq905UCSR/O73zln
VMR2Zif3MUTzf+/2XDRKE6LuveyYPHKwxTbdUAoj6qntmvjb2igoOPasLSXYmml+
rNdM9nmuOtzP2wAUgqQTZQ52FQ1S0DZXyK0tzt5jbDh0gdfhJinzvz31bJUq2gsg
pPFrVmo4ylwFEWHWHR8RYnBkTbdyBe0AbCfL4PLu563tK/4O1IzO+KVeE3wUyOSK
/dqwpQi496e2Gqh+eVlfKLkZ8rfqyutYRQHFXkLLUY2lmn0Ep4V+b7nDAaLj06JQ
H1CzYOmlQ7NdqAFK/7w0IpAaqw3Xpj8IAXpT/aayL5QEDQsx5XFm2+DuasMPKRPd
b+gCpZxfwiNoInoUK+0K4v/5QeOxcPs1FiobsbjivuOcLSxBWM3Yjv2JH9dgdvxp
JBJu86oUDZ975GeaosrLPBH7hNCvYsRxEUpO5hfwz5/P5q50sIBqUu7d/9jyko9u
MizMvz2ecPrLcF+1ONeFXp4BtS0MWF7yvJ8Sxf39RmWyAHCRWXXsimk0XEQWVJHu
C39C9YF+XW5sWPbK8tkau1LqdeauhkAdbgz1Otvyy7iNZ43eUtdZA3yMSKztISUg
XffAqEC4sPeURw+ObPVjQMmXkrxrLX7m47/Aa0sOlBe/QPbH7faan82MDl4Yo+SB
aiXAXGoeg6fnKIIy7O6QKLGp6VsnqRKTQZTMf7kxb5EqD1PAvT4MED+P0opzTlGn
4kzz2uoR40JsXX/cPjiKZf9OyGuUxZiAPAbQ4sKbO7dJ95C2HSQ5jSRDJTJM+zaG
jXcwcB0EcM05Kuo8y/K//rexaMPOn49SQZZTrBs4C00kaqcGZJlp5B1DP/0gO1/n
qE6vwSZzYiNhbxuKIYFzGnkfE+2VcJWiuT+SCChTkBWTygwIKHN00DXlnsnF49ik
jblz2DDmO694cfW1hctQLazh0be2b7w78+gxrREKU9Xy4glUAcf0co928qPYVgts
2IMrcaujXvXlaJcEypIJ2YkMZkxaEHQj1adqtpa/BTMst/L/htHItFc6XSgFKBMC
HHEljukx077Vl6jwo1kkJPC0Adz4Jc/9fSzG4XdychEYRTIbnNMM5COD6coS/esf
l5l0aHwxhQQBejzBuFLlawX1OtnHIWTmzDUo/X4fDoRv2D/qQjn3KiN2MlaR/bRL
TaM7cZEJa/7eqfuo/aOhqPTIIsrRDh7qcRurhg8hKsQ1pK/hOiu1aY1wrHYj3CpC
wq8uHtlTxl1MIck+F4CSObWUCcOGG4RbTY6G6tzQb6N2YVXgYrzfYVAFUlrO0OIT
WSWaZqeDyQLgGTrQQroereuqnyRYdiYGkWc29dlF+wUmcRwQojZh3frYwCKZNB9O
YZIQnkCBi1AXYRXd/3TIfJxEcf4DimXXb77J/+AG/EKzBfL8IXO6Ys9dwrpFV5an
JfpDXE4+wp1ACdyYtrWWcsXpAxpJDiE8KL1WSHcp2FVP3k+sUJzlYqBP+htOe3sH
+jQMmJPiS+B6tP9AMwJbDJjZfLt5pnIMQlyWQLnMaRkX6qOMTtp3CtbcV1Y+mUmQ
mzhXr7FJCO42mb/jB9Mo1Zo/7BawYzhH7Jc9uHxKA4gZNNQ3k0VOBEFBTLXHmM0k
yUu2EdONU8vmUCNFL/jBpmEdJjZ0t97AOOJZSseoUGkl+XB4l7uGJFCDt0+JsSj0
Ruasy6OSk7hHqQlGdqGf19Tzk0hlW5qY0DW2Te8arC/GaLU3cbdhUzqWv9yeQpTj
`pragma protect end_protected
