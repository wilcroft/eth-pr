// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:12 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
X72t0/5himoHKtf2+1Oi5BLUPqZDdF8UQQ97q3wtRU7oo7DmL94EiqdQsKL9n6fD
ZnSIKuhNXwEOlG2WB2+VucsnvfqKmxTUrEHKh48gsM3ToC2ir57elGHhyDntFzHK
C+nJfC7SX+DoTWxglt49qdFq/8M0L3ep5B6+UUJqjyQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 23744)
HHSB6qL8IHz452sJ+ToHwgnHEKZK3WQtZ17D/OwPnU6lBYYAgW5VFjaRuqsuuX9g
+mlyzoOVpPT2Vq6oINiAnTD1gg9rUPCGIE4L7ThlMR4NS9oFpI+iGkF5arRQtFGe
huG7IcgP09k4qxmdB0bahyTQIJGecYPRAuYWOAtdse7qriu5HXa9j3148TVZuNMb
MO2GCFozpZqYPz203/DjL1+OndsaWfS1TzPuC6Isljwznvnjga0d1TVrzFLx1Ws5
iQT3OhwJeXOrcniELzGJzXJw3M2+8xwvq8zwKgr9xv4slmlhYkwUiJJ+7joN1MKr
3DQnY5ZcFIGtWv6cILg0vL766RxzkG25JRGQh5v8H0d0AhYfedAxAFYh7B26PTLF
uDONhYmdAUS/69AHmK1FXzIusvFY0sZSYYps3sJ5D7RoL1zPSYCaiFLa5ketOU6f
U6blhGvFSWVfgT+fyVpsaid1JOg5w7mTRrZ0F3APAa0CaceFsy3reVkKm/UA6fUg
f7Bibpcv1Mcqd2lB8baE3Ap5ZPilld8yWMasmEiTQTXnaXz4DHzQZ61P/PYBWDin
X0CjWI8iQV2YMI6gRYmOsrUUl1Kyzban1wWZ8b9T9rs1PbP5boUzfetOJ3ThSmbV
XGFo0COOc2UbBgX3UPZFBZhI1QIYPOht9axCAzpU9vcwlCEq0Y+JTV+rFAgjRPJY
E/Qec4I3L1V+jIqb+xujiW4Lx2TSx/INQhEyLqD8QRlqUcEPNBtagRTBYHTbjRcf
DP+wN7fHNFRmobbV+UFtdrHUwxRKhKYHctD//SMSrJWc/JgIBJ72nbaQkmH+G9k1
nJ58q62wRoy5qyznULPR8nbAzLtQ2zouZGMJHNp8w3ikxMyvVvISYszPlwmpOOtN
VZ1iiX/AShvAwF9uHxoqsHc4pk5nVx9zeVlSBf4iF0JBBRWSp8g1Ju6eE91DN4Jc
EQUX8jvDKa79ob1OGi2o1w4pV2fxR+v5PPHJzAFCvVYiuJswNOPzGurBXq4xWkD6
458RorVvGMc/0X52CH1RClftd2YxIpL1PIrugZ+1KQ9hbxBqMaKZGD1yO5y4KdOP
7WqoB8FHgIZmJmilpesqQeYcfsQKebb51R1d8/stDPi5hb7h1h9jNIuXjNXpPfJ+
5g/4+36pRbYr49h4QMkPVF/QDc0dBrD98LEE/wTe+C/fgTukFb5W6aFA3OO+PYGM
fnoqmTmqxSrOd8RV50C2HMHUJ2ipSLzfGX+jwabJPtqe9v63Ml/V/9cZyD0zN0HU
f2KPNpXZ8rw/84rICXeS7oiQWUF9ZbSerCOYfxVvzbQaMg0ceWFS/PHJkVj5IJhV
PwpWMPZGwrwp1X/JPguW1DSvYRMT1VeOJzN1psc420fyFhrxZQk4J9xtpo/C6Fxs
MiiTa2cam9yle+1WleCqZlSidJHMqVwGi+X6DzdNtQY3nd6cYcEDBToj/kN7orik
/glpbj2LaqghrIVdbx/1dNOwcZibHPMqcdDCdxREo74S/vJjlblImR3+/xsShVo+
U7GJtXLf3RTDlpo/WDj8dp9m0wXn5suB9NL46cVp+Fh34bbToK+5OpULSB7RFkVf
nKIXPhrohMG4SGCVHiYb3WRSg71HMBkexOIpYUkechGACL19Y/0XrMbPEl9CiZqz
y/j1dv5RIiK4SgYM/UjJ+57kYWG+mw5ijWWXy/jkCfMts3ivaBxWsEb7KneyAQqA
ScxM92qqGTnil3qFgR8BK/kGlG//wP6F8I+cz0EUydfBVBOkBlTbSYOEpzlir0g4
fOD6115zcsouHCOewITlHvGpR5qSjJdAMzfoo7nj7AXXa5W2fQBIKChYqEg9NnIE
iQf5+bPZbNbnTWkoF+XkT+nCSbyHDZLHXG1m23ldIk+mJwFIJHfq62SlQkfg/ZvB
65q/yHIWm+lz+3N7OxdR+NwWYfzMNzL92VQWIK+pYkeHT43NgC+y5C3tPynqXM+6
m7UqCQLVrw/y1GJhUeC5M0xQ5gNNiSUiHx0XQRotfc9O2OgL4CnnpJDpIkYHchLN
BXK2wJpAZb8u6w8CaFa4okIVNquxFmPrqsQwF3r4ic4Vb2rHJoFsT9TLupT8Gg0J
X4LfFfLXUvhG1lQGaZSXacHgwipSBHdSrDxgAEeITfhfxaSX+7g4CJpry5fN574q
SKRVZuuNB6MJfCTQQfUXgbNaL959U0wiZgoo4AkB+dpv3YQ86OMakryk33eIqqBk
lilw0Qlqn5cNcX+Pv6ixSfDFh8cS2yJJjcqqwRWqEgEQ8qMIiN3vN7dumshTrbEH
vZbO20tMPQPZZ2WXDVnzz5mM9CtZKKEhFpjtAIAk0bzOEJiEaLN92ewKTJeUvHne
eFMD/10TfqPaZfX5yeSNrepajeFhQbw+rPYgZLAI6+h1qojQBRu1imy8VJ5koJxF
7iHmlIFXDV25wml3CiFpfs0uEeqtt+V2bPt2rnqHfv6LH4zXbyx5cuYHTTrWjUt7
rRYX8ieyqv39l6/1Sh7qey5F7s9BHNlxuzm6Ptx9CgKrpqyDTrfYT3AdDgwMjtR/
+7ovGBkBa29oWaZ8IP2wZQfAAC0vwGlXRqnFhUshhVh5Q+6XDNenlJ2owhbdqVbe
injyd7t0wwDMhGJSYXPhoMVKmCP4b8gqDqd+yYuDOud2eZeq/CYekqIuQrU9YR9K
4uKzQ9ZMMYN2gD8if8s90nBXTrRCZKph6fyizJ9R1zgR2cL2qT99kfo7YY18kaGc
YZ6auzCkteSUh+5h7iK/jxkrd8C8lfjC67yIqraVFGmvNJlPf2GZletMzmCzQFHZ
DsL3/Jqk5DwC+UpnFK1HF51C0lCS6bR3hf6GiQL/g5jAPrpW6aRu6LLRIfFjB6p7
LA3HliU2OWL6/hCJmNTpozbc3Ww6KgpS0LJAAlVuf7ft4BhNSr7ESlKSYIOzcRiG
pxS4dEFn5AmuaZ4C1VRRyddm+/4WydTnzvO1ug0XmlKLesHXKOrOVAwZS/8tp7JU
0ceNXscGdtXBC2EQrWE9PapS6cTQweAcyitAfh4b08W7cb8oAs5YZtqGPFLyw/OZ
ur2jp7advDwGD4hIS2pYC8gs3ih0nA4iueqbgEX9DObkYz5KzBYyQ4RuF/ZHgIRA
qNKS+soTgyXZ1Kzoqf5MHF/Jd3qd3MaFkOthAVEao4TAVOp9Tjc24twHw9NpLgKj
3/hiGDdnM37SSkAI5o+aJY6CklIuY+KhdUfEJNdBDHW8UHPIoo4i5U4TKJk300ep
lurutvgvKWAQyJPFmke+/I7IObKMkks9lLFW1UCmGaPfBhC+Bi1ePerxKzCmEC1r
RB52rz4YjHzFVvJo3KcgUnvyHG2uBhd5Ud+C/jLSRx01r/6Vrct15kUxougfiEUY
XqqaOSnd2CjCQPKNWXQKWOG8HAcpaSkRQhLo5vVA7nXqisa5AsCmyCdu2D8QHTkU
e7qPPJG6KfTYj9nNx+MeoY5rJCYoja01o7ubg2TlZzisoxcf8oG8Xi93X06lU21A
ELl1mSI90+XE9vhgERqSbBUBMzr+ZP2nZRiZqkqqmImwOpHI3XRb9xGGNN0+Ts9w
OiU40tn59+ycUeVEqMl/y8saC7UhLyDrwYEXbjMHpXhMgSEEFE9JRILTyW5CDccQ
MWVQbxwXFakdpMqWQlzjrN7OE0pGO8oHwprBpFHpSblLRAG6daW0mWOKZTxFIw9A
MWWYUbbznDjnexx4NdpJEuRBu6Cil2s0B3NKxLYwY4LdYauBdyZpZbwtOrm2uR8Q
XxQWV/hRMS2lTe3d72HPkPxD0EgH+dZJ88WeXhshnYvstrPPbCQmqldQY7XLs0F2
7UEpgXOQQDLBdwGE16pdP4WyOBjh1nqRP5IDZ/r7D7Uwq2PjMUznXOWnNFtQ5ODj
VYr8qGR7MF7SyXmLqQWFhSffdzXO28umudurHx9RiZuHfrlUraWBg0r/z/jublCx
HWi4ot8snT3KWYJWCl+9JN3kws3Wk/DpTFIKg3kcK5zU+4PHH5JMPzZuto84ZJyF
D9oT57JylC8T8X1uJMlJSi8q1hgIw0DmyDoupAtbrPaF4Dl5sTdDqBdfBmp8INhQ
s/4fEk3e2d2KcGIPxPBnw0EWHaUsz1SgYFdvDayVPELh/rxkoyyg6MNA9D7JaJzE
J2IWyoU2/RZEKIJwiPigDII9C3+pJxSYDpkwMPPuEAado3fdzyHKD/zc6oEMGhgG
14P9979N0iAON8kydsLg8WmYtm7tfuQBiDTN9ULjl0tpr8K44HsonvGInxZNu97D
ipnMh6bNBfZRUW88bVzFaZRKu9zw6SLHw30K+IZfSvbOrL4EZXKb9cBWjYZ0DqhX
bTSlKH0HS1f+OlEyRpLEplhTUfdTczPP9DNnloe+eOTAgX4A8Tt1IdSTJ4fVRUik
W0u+3n3lOylV5r3/5jUjlxuKw0rb8mz1QhUGQKw/d/szTW5MJcRIGR+2N2uhsBQD
uVPGAyXfcN9xa0MUsEWR3mufcysXiNpW+A6RVPsz3nuat9kaLhtBwilYSgsajo1b
3Os8yykrE7CVdFc5HS5xysPmK2oAW7wBdOLJTsJ81getmlVAO9Lq7D7uLMbtt/uz
JRsqYBqWqUtt2GneHH+hs6Y6Sy3dXWWAKDyC7FBZFLsAhhLkOp+PGCkX3O0C60Hg
Q6rXPmzk8pxELSQ9f734/xZOHaDJUAdXARUKD7AtAO7M/vHHvb434Wp2sh50U3EX
zGTLnKnHxPDOvAr5lhbyHxCQtkSf35B+8Pcbkc2yWmCoekXLvNCT44Yt7BXfoue1
jqczK9O4Zp20J8r7GTPcsvcan7d7lLOSFLxZZ+FDlzdgoXo3iriBbSoSLc6Nugwm
vdm4LivM+GNfMtEthCiiez2RoCNyZj8Kcb+Xb4FadDoWHWJqAAYQVCtZ6r8Y27X7
L4tJQA2Jr2y0kgoZlOQnknmn2QqEULed0ATts8ZJEIU19uAQsUh7+YLoNUOjXVZ6
8TBqeTdDlRA1rTkJFgleSSctpcV1rtq3xFD4rrVmHqUg08uV7H8fXhCWoBOng91/
nZ8yi6J3or7n1fdGMMZCNZ+pxeOdIAjJxX9xSC2Q+sBGI7oMJpMF1kZ+T+cN/fFS
j4YeMY/vazxttGojWwfvDQt9Si1PTkMfHfrhh60Bzv6jnd2rQ29huVXo49FoAlhr
HSsYkddtnKE+UWgSg08lGFarDT7WaKg15eHVItsRt8oA0PKBAUN1jcpfwr2LURzH
Q6D6t9YZ3fVdyUjvk1h3W6v8NbUKTBI7q6tIZyppXvjuJNn4HwQTfuMBYY+Z+a1V
93Q+nHjScl08lhmpCKhHidF805m8vPBMDiYq2U9ntEeLrEFCUP7U7Fy0VaLR/CpG
95+IzRuRZdUnaf5x9KHJexrLc5m6V6aDBBZ0H4dHEmL9n+4OT+R+FsWEoT2kztm8
1vQo9UW3uxdnr1/kICqNX70aLZYFutQmkyJrC/Iw828zjT7vYxnoM8cBEkGLxEZm
jCXQr9GsaYzNh+y1cNvUIUhag6CSjzHM9OjI8o9WKp9Hnf9Nyit205tBzVMFlQxT
M6gXlEH4LFCYqPJzYILxgQoM6n9zBj8N3FCBDDFXijPV/dg0c7w1WISHOtRtP69c
LTxBEKz3E/BLyAU0FI6hRsFYeBe7KOsFLhj4S6WPBE6g8pvY7qfyPI0qyUn08pnG
UC1EKRrXp43YufeFp9QLBTrYGspric2hVKzP3kivpa0XB+tCSZDUQo2voki7VSuT
Yqc2SZ6RYc1yXsfwKz992l1DrNB+GGkadChxM/+byIqovAoDtmS7ZpSN42FdBdRn
4VhQLMHt6SXO9QXBzCVHkPkDSiDfejyaIXFaJiQ3Tegrizm7A9uWl28LHG6srn3O
nkbuMDVfOVxtmFNV0iS36QkNQC86gy4K2Ik9bZmfzDGXZyM+lkk5LSPi541PYl4m
e3M7m3uKcpCW+fBVf9a6VnCq+/ua02ugoGWqAqUHoPE44RuJZ0U+sa/DJ5J+biSX
zFm1cH+7jI72eYpqKa9RksptJLerpubBTz8gTjlzCyyJXDjtawKjH4f0FbPYg2nC
HAAfo7TLNhBL0CeAtY2isXAE7KsHJ1TdTsP8Y4vaJHbYxq+W6iC7ZefMDSUK3WO0
cr936JJdOGF7pX7MkFAWeodmiWQsCBsyze0oUbF6KqrNcUy3VAPrTQ+QZ2b4NucT
MnVuFuCFvuZBfAN65acm6FTouxeNGQMsVjpSzbZnVN/xjDxxgqpFd5GqZ7ZtmCwB
dd5F1y8TbfB2HUVNLm9I/8RZsDr3MJWfTFpzGObNdSAKuGf1UZC8wNbPX3Tl/VGl
FQnHhQ/B4E+vx15xO+6Jl9STGOZtFmXCEOZe9KMKeC3iHXSEafoGTF4MbJEjrQXt
C/SpU+jzMVO17z3X5pgsDj2Zyoyr4WkIegedxMitLiUQXtyZDBdH9j+MI1SfNoHb
tnQP+NVm140gvjt0jaaBGwmKU6VWH6RVezJGlfki6ROH/qaN9Im0T09Wp8/bSKMB
0WBY3n5NP2ne0OLXcRYtL2XrrCrc3I9T856LhIDzJOKnPUUyirQP+duvn6cUVcg+
jy09TXFfeLqWtIVbG0AKew7ONHRPIpStsHEWT8mEvvE5YUhC/+Gmtb2cBIV+aNUf
xKs+goh5wo8jLYgiqgNOV/DsvaC3eCiTpAdntUXAgIswU4hBRusd6gE2HC9i7JxI
5KpSxufU9yx56O9XFfE/igBTvKNfGKxTMPZdKOXuVSzZlwWi3vHa+OMm7CnCS5h0
szgUCg/9jsoQirEQOkNh7pg1LDeJOcuZ8IlLQ0DcSri1gSRjSI4HAZ2j4hyxgihi
FNs6w8RzBhysE56lnVkgozLk7teOR+MqJ9BT4sEN9rMk9UX6Ra5kUQ4GtSwgdt6u
abRQ+yJ5z+nyArxbuWvCG6aTOLUSJPl3q5V9IfGCoweFYSBbJHeutgjekmCkpY6+
3MSTiQjg7mOOKXokmkCPIJolRjYbpzAO1ZL5toX9+7Ym4yyPIP3euVR95JaHC0xQ
TFprj6/SCnOyLpfvv4MVE1ocIyMNjDcPP3EV+xZb1fHs6d3D18TpjHLKwkjeXtAx
bFBHWdeS0n9h0RhaOzD878BQFplgTweQ7xgge/Ib4tFzckFcTkkzBaLCFWGdfvML
FSzj56WW2UqQYD1SqU38rFADUaWwv8NRc2fM2VP/fBdL63wYybcp2oeqQHvIA834
WkwdVI4b6vFQVu+Y6rHgv5kyaqLlg770SqEx/Mi7+LIvvuaxTNNeXzEENHXTgRv7
8uZ/tUPJSXOPXxR6z544+vpVMtlvxMSNFpoHyFiceR+1AKFJZagxvb+tcXqyw7u8
37G3WkkwA5o+vCtTHUM/usIfGo3UEH+FX6LT8JK5e+rB76qZuIHvhgd/G+4rl/XW
CR0DPDjxMRFQYwZ9Wv9WMkwpg5quYh5wf4H4wU8iUzIMUx0cBhSO1ZEG2/m9pArD
0397eL3F14Mepc4IQPUVDVq9UkFcrae1b86qbFa75ZgamL4SYgTc0UpOwIEuR4mx
luFOgPQ+BB7KPz3LmJt2Fk/2QhxJYu6ULEHf3B3JarAol/nK9IH9W3puWzRMimVW
ZDwHBzOPZL0RXxJF00XZH10BdWBOl2630047spgHEY0pPtLGgyczxQbGBMVdrP3K
t1+zmHU2S85b0fh5NRNSAGa9Mn+MZtxSua+1grqHS6VeLLTy9GCFYpXLgDAK6c6X
WP4/uSIBvxDknUTm16q28cbY8choYibcbYVx2AyTgfQZVYyriu+u7q1bbC2W6qwM
4WaveJh7yfoKBtUaQtY06CwOhuIbCE0GJpQx83aJh0qaH0Hcoyhv12OLSiEXaUVx
czXRh/a0bI83kiFSCLwVCMoqhKiXQ7+eLSXHbkK7kBbQEZ6Zo5M9b05IpWvnfAE2
TxvvgJGRJCLCQsaelItAaJ6UK2RAVMiAoiC1rqnesgcuC3ToZIPKtlLsLDDNRry1
HUxnIaydqNAeryAi5oN1X7qtMyzkMujpKzIfiSdPYUdnSBcen6yVhIoJcPYviZf3
EJgJoizZPKVTBXjTIGzEEEzauuwDle9pShazyD3o2GzoyuvVaH/JEM0csYzjXJs4
rZFqRW/F/Iwk3l0A5XCjEnBQgi/8rBVbgRx/S4EvP836PCq/FxbjDOtg17ZvKIJe
QMoFOJlEYa/QgcgW4eupk4Lpf969tWB44NG8ZHwVqtIykbnhoePl4eiJZNVl4xxJ
QaQF4nKOFuZuNfrDw5NH1hJY8T+GAR20/OlOgQTvaLCh4dpzGSnOVJow1hUZg+q6
8gpbejO3Rk/F/6A/GA0/f7JTWS4HayOv8XEA+0XW9I7/PM4jJWwqvL0uG4gJsd8q
0jom3sHJ4VOfApgXOQfJrcBt5w5Repsjp8clImgpw5b0KIlCKYyX6hkapG+PDKRD
q/lUJkiO5TqJ4mNKWlib6mGwML65TPWrCDWtMKW1j6QZ6fK1WbFgzBSd4sS4PTfw
opHiEAOtAcjrfn6FMN6QhoJk2MLigG4pMC4FnT8vnp7SY1D5lF3dXTCeY059kvca
W2MA/TUX+HLF9Xui/v8b3Ig5E2ddOy83227IiI6oUBi5jmQg9STIWpxbjqNEVLzL
3Aqa+AmRVRtYy7oWS8jT2mMHo2nwRu3a55cjedgf58MWYDsgmZfdQF7RFwP/xjZj
5diIKGX1nApLumWy4r8UzSWmUIld3Bi0e0CW6eLOlTJ2gw6/XX5UJZnVQjNrHdD9
1uP3q48/pPdHrMulEla5Ho2auJkmJBg32UrDsNBTZqWX48xGFRHEpQd/HCh82oGR
lo/h7zLJVG+MVWzBjkLf2SjdgdLj9M1N4y+n20alekgsdjPYEHPzZu0FmFq4qqpe
t2IHVFQPudsUWNrRQCH91IYYpxFuJEElqDzJEjv9CsAuOc5QGZoVF5vogt7C4eq/
OARwCGCCEWe1JABJQ3yyAErRIUnq+9eyQkeghwmnt3rEL9kfga+Mw6JW17zxfNe2
5+IARyacnM1cUicbMejGeWcXoDx8a9+k+iSy+5AMaPcNSHu6RwsA08VlJvDt0Uqt
KYrbQYyBVw2A6Ugaj2rGRMzRg2+xDk6ILNaNN7/SOHBRQeDp7el2MTc/yOZ1wMOk
is3gymLKWAOetLyqkWrMA8S4xKhHb1Ypn8qgBlW4yON7NTm0/x1tDKZPyhmQ5ifU
PpsBZcSUE8g1ABdCM+P9bGH6581zjvbajdWOC9eoBCdCohb5AzCK7y2Pe5jEwwjb
ncinr9bWN0mR+5tfAHos0wKORRdfadWgK6V7kTU7667V+7NaIfSDNLEIR7flD+Fa
0O68to6TNXS9cViNv7QkE1zYpp8WS+RQNUsZkmWh8M8REKZoueseXcxvSBKlFZ+m
7b2rPKxLMPXwhLrLvLfGHsB9maS8JhJdeYIf1daNpDDezfOGHYWQXNdS32A/dhqU
lESAjxk9MPwd4ejhwEcnnJsM1IpNATsqEeahw5irtg3gEmX9kcyndpyKQWOp7K/5
Y/vJYZJiNYZ1W9VlZ1vS/xjBfRBzWWQMXIM2GV8lqnhJao6miJe3BamwiuuKM0Lf
utWa2+7Hc+NYvgWWP7qxrGj5LzWy4oGl1vkWmuSdYjSknlQwpKuJNOzAsiHPmU76
BR2Fn1oD2tgtNR264gEDEUC3EDbQruX4oRUNkf9cMHP2CsHG5zv88wcVea8BJG8I
oA96T+kFFOr9cMA+jedBBkb9k5gTM4zW1h59XCANeIqNiMkJwexz9I6ZsvL5WQrL
TQRj9TdDcJyi4IIiAiIrFgQRRERv6Iv5Yfp5HDELVCY2qZCNMriTS+Rpcs2fcQAZ
RRQ1hyECg63czTVs/kqt3U5CWXJYmKlc1I/YQSceDYU5GBmkPiEdUvnmLwclOVhw
nqJIYtpBFRFYnHDwXUsPIMP0uMvuS/VgG06IELcgOmzOhoo20xzZvtViY7Ki6752
Lmb7DIeMwaWyzRopXdeV0xJyglPj+UUOO/H5uzicCQQHB2Zfle6UMHz62bvlNZca
LUhHDIDB0ph4GoJa0J2LXjr0CjdH0SiNb5/LkKY8yyZKNmqHIh3OR5M+dyC/Vsy9
CmEc1/BZWWttmR8ivMrXP34wteXAjsw7+gSXgVAROwKktgvIqVX5UwJzHFAhIxdf
006ZzOlO+8cL47LZvroTLhaULcBbhbyMe0jy+5a+Fv1cfRuY2VAiEvQMoR9JTMOx
Vn395kd5wd3mJKrHEWaAPCZq6Fr1T3E0t4WJLqa5D/7Yuz3beSTfdfz6aeZXOTgf
wEZTpUVZ5mLRJ8iOge1gt8228k52/uYQDugdbpvz71yaTOgXWW0iBZEECGORGXBy
tb62O6J/jEHQk/8pndlnuBOqAUsqtWmgucXJhXlpx9czR9qnKEDs0IFUv2Wo/B4i
aXF2Q10E9xbZ/PoOr1CZBYnqCEGm+ZZadQBe6ZIA9SsWIXwKLWTBRlfRb4psJ0TC
5n7BJ5MprZrtZAIPkbBtLl4HSiTads3G3WIh41jVjCn89Gv8cfB+vW/3+hlU8Gc2
czaXBZSWXVgeFImIeVwD0NS0Jb8XY5BkyCc1bre23KxMVsiN5ojt2GVAsEnB2Dm4
wMcmgV7jg2M4fubTr/xN2fbVZFe3KxwsKcw/jkw+UFnJ/17RXu8aB95IehpRtwco
Uha5gqCtUg5LOFA/JS0KSTwS+tHoJJXBwskA9JmGpkvDbrQTq4JbjpRAejelRzeC
c5k6K4cb9sgOm48t5ADintc7X/o233iWsOr5K7RM5oKzH3707iX7bLCW2PdxBlX+
rnZwExFyb+Ob5CjhDJW38FW3EYphV5Sw4VhtST6R7XAh/mCYGVln8XY2lwlBIAhB
+G0te0kyo7JCJiIvnK4OPunn9EtEE4zM9scPhsykCBe9TpBIxDcW7tnKKy2koTSj
G05LG7o4VosAg4FuCOa9LA8lSdhPey85tfoCBoQcV2aPb+/8sdC5jiaTTfLDswqX
lxlaAoRES0ki5vND93JsnArHPtEsJ4zn53ZFvYgkBIAUOyf0hMxO+U8LRigk/873
tru2j87QU1rD+iKeyLZ1dNq54Bx+/ORul06BZ1VhVUdEqwe99STdnGcPCuoF3Oua
Nxar9gIW54w4wv5bG+Px4i+7hw1GZQR+I7p9PvI46elcbSv2jXZ+YKrCe9C2Eeja
IvPQJsTySAAhLyN+x6aq4j7FLIrYOouCL8LlMjQD4EFhOYzQya33zSAdbSwuxb2W
Ft6LcpG2amh+tqOPCM4JXENrO+O88tyQjX1ZO3/zgaOJdQWqPWidTfBJ7n3Cwags
EWR/vLPW915++Q0AF0xnSJIZkp96UHuWi4+/OrSlFQbQXR8frPRSoslLl5RTGuB+
bXs5I0F/GpRBmHn7aQZHf57p6AM0xyHJvdu5UWKvgksYk+e8hQwy5JTDdBnlT2ub
6bHF7p8MAkhICSitJi0K/oReUjkmfwXUGtqkLyEDDVWEnsXplivxeKdtexSkuS2h
flqsPYHQPjtlJMENWf9dpDLC12hQtYgqftv4JpIPzhKf0d/EQjwG0xjIobQlS/zT
Zx9tR5R76/IdhbkNYp6bBx4kOnN46ikHTq3QigmqfYIgnV5hO8KWRU17rqPkn9nr
ve41v1cfQSZMVYQpNTVaMY0ROarZdlgVki/8nXHBi2rY8BZ/49iMCHVYsAEQdrEA
6VNPiMGsruLGJ8j5rkKWt5srntB0Bh7Tl2Z5M7stgGVfA5Id3rETKBdx1HkXNw+0
+gtoW5589SAhJDTCW3jdfyjx75U5v5YVTHhYq9+1DB7VwATxRXM11FNyjC0Ma50t
A+s6A+VHeDSkFiP5dKHsK1JjNQTH803sbiag8PVlNkBRaUnqVRLNl9+//TludJEP
fFerh1muxMqNw2W4MhxPKoXb62Iq5IS1KIJ4POw2vt02dow+UwgWp7SzUkbVk9OC
Ji5jRk+crvwHqZQFCI8N7iPYXyxtl7pZ1PKjllXKl2uBAbEMTdodtl4SnEkKQgkh
QoWTcz1EwNl7xWwsdLgprNhouXaAYwBe5p1QSpjTz+1S0qOFDmTGx5+1xxfMwfdR
GsihdhfY9iifcv+Rhymj4zSf59DWoczeXC3JSZim523eeG1Hvmr5CcgCcDH3g7w+
jxmvbOmTPcmip+MXL2+euw6+0sBFOOX/erP3fZVZsyn0EqtAAlKTTNSzoFzC5JrO
u4e3vX+1qxlkl91616jQuEucg+gQs2y3kJ3xzYCMInYASQnclcuQge2b18EUx6nH
FINnrGIEtccDnoA/PCKZkyNomUEVarER86KsJZfDGInghH+a+HE1AsxdYjdbXVvp
q2xT26EW7tTNN5N8yh2hs3xz4O/eht1vmEciGtE9yarfDWTwsMiUCJttt7Xd+OBi
ZlUKcS+dA7rPKfZIlPCt5JiKjRu3Ldxx5K9TjIJ0c9wAjP3ldtEdHzGJ58YUhZMu
SiI8um+3A+MqEoLrGxAAO1lrnXXdS3VLq1ltARpnxRVu5RnzTQjMi+gIzc71lqyt
m7OZZvzUWkiEWYOhMxI2Gv06p88FZPCKZEU36ih6yy5avgtVcHnhv+ud7GiaMu2B
fyc1gCAp3K5dFQ1Nr9sPY+krLzrcRoGQWdF6SKj9hejM9ZjNGMI7YEKpmlk40sm1
9Lmsu3WuSLbPcEtR4TmXwyQvDd3Dej+cacwA/wwN0IPGGNf00Z1ITgZri5dUg1uI
KcocCJGPejtw1tNXU1jbSjjjUGucyQjwj+BGYOE1tExSvtLm2bnMk5h9rhq7MNUh
+gcPWibfqd8yEL39H9pXKT8SNOOx/NhONKR9vGXX0NeceFLotlkbsHlYIxaigD8V
pYIeYBPF1R6yDsuNqXwruCYF5gZRLxRzpxmQfSSgKKnZTTaIV5AX2G7LkVnD2627
+gHMwh4FT05ln/lpeKEpRTC4tkEFr30MLYaAN2Y5hl8B+qtQZyIK8E236ja5Dc9B
goRlUFIR1VirW46JtQvbfzXOVhz9uRsUOZMs7MkC2rQDGHZ9Iql6rknCJSsIuGXM
BP9n4sGK9+njJrTLP+3Q4SUQvDQiJbIoj+XGQwUMdLipxt5Jz/r41lTiXdYI0k/D
5IwxfR3Ng9rVvxshPlt4aLBh4p4aZk/WTk4pVNsoLydjn9wAez7+UeD/4GIUL76g
DOFEMT/IdsCtZjfiaH6eqhoM9vE/l+c1ttgXXzD+wrQkgQeHUnpO5t8N20buUuVN
znr1f2Iniq+Aop6eC3I2T6lV1iAkn5hkP2yTyPCRPqEs8hAocUoHFGM78uYOyS/g
Zo6i2+kIpmbQLSHmq/tOu6wwU4CaOsoLw+obeKG3xmxwRyVylz2iP5pQlIALL7fs
Py66uOI4N3p9+WZUR4loFm6nBp80AXkeWrq0dw4wcBY97ORwLn0UcdkgdYctDpe6
uLna23xTasa+/gsXBLmz4Oc0pZmcPkQfQGMJ32zNXWr7M+B83+2cVG0o8yiBHLQW
hzE+rh43ZP0sBCyXZoSRGGMzIKtTbdnTGpcjLDLVHai2/994CnotzYdsl3mtcVrW
nYdTWamQGVaVqMm/D0fd3dAdi7C2xgpOrJ7qjMLEP1+iZeiiBUEmpnM2/3//UEnb
YXr4tMLFrWnpyq7YsnjUCCSI+1Y3FMoGzGguST7kpzokdrN+I1qmRfq5AGAZFAF2
QUx0C3M0ioxlxCtDawiWKnIvDXDedfOXd0fyoazyXZrXDg1eII6j3a30b2API70R
oK4H0NRrrrH7wX3PM9AqjlTm6ZfnZ/s37ycCwh3ahy/+CWdw4BclDNxqWbfMXLLb
5/yIGueAychCD/I5Fg9DIIqlmALO8deMfxEr4ukN1J1C58vpieigIiPKlwx0sPm+
hai0WvttHt3nnnNT71d1kfpvNYlQYkB3dGfmHDSsuQdwz+cb2ztFf+LG7L+OlRHF
0SLzY3l6nmJDVzsbcUo1ccGAeGAx4nlaBbHgypOM2YeB0B7WMhxHCH433k0+Msjm
goHLv2dfBHxqy8LtWxqd3wFIPtRPI7p1+ftUHUVfoX8f4L0sUnUwBp1V2jFSItr7
O7vuiJs7EwlbOEg1fh9Eqlmet0V5Nfd7QtWNDdsqcdyZc3jd51xfn/4Fex+uyjtM
AbUaPtT6qtsTG/anGa8b8rbXtaZJcRcQ/zmfCLvUB5zMGe1tDOU83AdsRFkhgRmM
jT2VnosvIqV6xcOtlAcw82xZYXK8mpVUeHXZveTAPbFvrhulWisuK7zb89k/tKkk
utRcUx4hOjhKELWrtHgTpIPFrQQvyBW3QT9Gu74CKrxyVSFp9tRAdxGX03MwPF0L
nfYJhQM/lpsOiSQJiFIGi4j2yIJBjCeQaBQkaTb6py9vKmlsSo3GTPLVlth9/jvb
0lQoaiMITMlQmLvLcavBrsd2vD5JoR81zhekvt8kPG5Ca2A0E6Im/kL3wAbf+Xn+
05t5AP4qYqH7PAUdMc5KrNusav6NwIaDZYUiiab3IVS0sIaOfP0Jg8+HaZsUoRjs
1LXIeuSD2Stdp9hVzRtZhKEybwmuENqtRYFIXUKTeDcoHkI5k6TSdz1xApvbm6mi
CW/nckx4CtJl0z8MRqawJ6/t6wNaHHqoF51QtXph90hYM9CElayKjsV2Bocw5ZiN
wb6q9mmc5lClVSRcAXVmu8qJ9/qFj9/pZWmAJwQ9zwsOPwEqnrmK4NO9YmkqG5ky
EChN7Q2/U+xE3pACRl/4ko4b32paNYU0glJ+EwYSLOH79ruJEwDut5KoG84ItJo2
B4MXng2r1higJIlPKUoaKvdHqYigGfGE0/82StXRsS0P8mHS+J7tDCUuzBRQ9nvB
vqDcZh5mig6uTPhAaEUPMSnCJN40hV+JOevmE6njwWkfCgvDZLk3g61EDj5n4FiG
v4T6GBFeUbfzzazEMJisi3CHUIEcK0Hc4xsLPFbTAIZFN9mi4eR9exzYA9JhF/Fm
8C9QDg+BVXhLoHOjB3F5RemPNRjuZUOl4Mb287mv11Np4Phdd/IPSQ1AsqYvFMdS
Kqike52L3vC/d/8kqtB9qt66xg/QlkBrwA5DWXxa79XUcm2VYOBoL18XesBu3JwL
2U4vNoYPeprkxOtMeh9pCWzLNR903OcUwSbnSs5JZ1/pG6wOR3wkYqgWZwx9OOZD
U0i9qM1ncYTUcUdSNJibXZx+vqshMinCuBma/U3IZfMcRJEdF/0T7WfOnxyZtybD
spXuChKOIsrlqifVxlWbyVjql8WD79pjdpVzUw6LJjvAhUmMvuxKfEChymGLUdOH
ToljZppTHSWBckDBvnam762fMwbbiNDI5jfA0KguGQwDMVqXq9xUjqzXFGhgRLjo
RzmdWijN+unvCwt7x/eUPcYz33bgKSURlXxv8xt+fSevtRnrroANau8ziKAGeCcJ
7dPbVnu7/49UgJpCwu0XHJnifBpaL2GM5WI2DMz7bSmYvkIGvrApXBcWt4+Lzhr1
w89UOEjefT2FNZTw+KuDh/E/WhNL3sCQn/KWoUFhRsZk74fpag4yoaRLR08/beGA
BZ8sESsfiymjvMYrXl75Uxcke7FteS7K/CFv4vLvFbg04NHTc1ePViDRj9yHc3+y
7mKNmd9HvxIjZgyNG4NR4yvGRBe3EGpoO49i6+fZB8qd6e/QO2/+T1D7BFqH4COT
Bp1zqh/gftQPb8vQpYAwyCVfOrkcF7j6pTsSWr3ihdmgrrKDOSWKXL++u/3DUpao
QD2Hpu3/8RnYo/WYzmHjkkMPo7GAlKgsJJkz2jX55YkA3CpzXpdp7ibRMhAulQsm
HXkp8ZOI9q2ce4heMrfj+uqWXG7w9jEKvt/UKnwLfE15PZInJWdsq7JOug9rCAfH
BwtzeLbp8xGrnFj7gv6JrGl4KyXQSeEhHYiCP6emfXAZ79536Ke7cNeXjGRYYxxr
LLy0r8nm2/fNA6XbLyM8zSXppuKwHtv81rnYNZge698WEa+FEs6DEfUjO82Cqldn
waesWkSvMnub1PThYe2A6ePwNSdxI+vVlNSzkNycsm5hMOSeEJ/n/alR+I3uXA5E
XpJo/ubLhPtd3Y3pDM2xlxxaA5+Nzbz0ny/vI1m5gBTsMwHzB/h6UbYy5yNC6uLb
0H6y4EtRHNT9bezrsRio00CDJ3/4Iv8Z4AUlMLQnK5M/MKlIaHccrmJ3JSyfiQu7
KJI56+YR8wodAGpuMXVl2rh+lQFkenVn0VhTq6cmV7/wGxex8QItT6f2A/04L4Np
noilo8mCE2ah/6iXD3+IQtJPJaLXrRRVtxrMP+IErcgjOqhOlAMAdlr/PLuPRVy6
6vljYfQnsCW9bkExL5UirXsA4tGkrhOIboOIJtkE8vZr0QBp0qXSkfTl828gxGEG
T+wkzFPpaVfVtevAUvREe5U+qOZ8IO890hvHe9HqUgss/iSPhJQPfPV4TIQHz6g6
S4zhMCZtRJ6eHzCRsyPrukitPBDsBfmfbf/BhNhPm3B8Om8E4dg6U8ubiRcIDn20
UpR/FikQOttQP7+2W116BMR5cNf8Uio74qXnu1N9JoXypfwZ1Fpe9+qWuM4P3uN5
BjiXH8YA5QinfR9wp3OPbeIBEJV1kNAgygVXlne492ukGKBANZRxqDa9ivdBKb8t
NbmpIt5vBSNIjNIvJ3tE7k7xG8Hvo0z7pK/roqofVymZxZnFuYn37dr1LZIFxxhu
Xj0sXMdjB9K1a4WiKqlOVSIjAALk8eBtcR66pcwcZDWTvD3rN+9rhhKNRFQQUIgf
LTGijT+R+C1LXFAfsrxSnLv7FR4LxIxcb4S+sTdy112+k6iM2xDSdVDFwtjAdCtb
WQaTjsnOCO7oJsRXl/rAebE7Q1+xaCBqnNUf1WWxcK/N0IvnYN5jfMPZGBPOCePA
JbnNsZBe9KoJVuwG6LQVxBsdIG2JXRFjUxd0LGhJOvW3ukiYw6ZN18q/ye55JSn8
9UDn1FSXlvihjjzVFP02Kx13GeAvQp6eR7MOOTOp+bBxOasgHyZ53OPofy5r21wJ
lM3ovrcnHSjtw1DN/YMQXsfCdNlorHkKb7ASqYrs1ygcG+AC6q5bHPpCulOyMaiA
RiNj6QXFIh9iJPoXhL3CkA1tuBiZxxJEpY0ekWFCT4LgQoFC04Fcnf0eVBzN3plz
Y52ZXT4KyrUdK8suj32T6GpzxQuY/bbZf6ZeRuAKkAxcTUKjaAckNJqIN+X5BooJ
V+0PD0GlUkAyVp5+ifSlHA2eZzECfTQ74w/3c0PUVYOKb1LI6n3Rt79F5nz0jPWN
GjPR+eSFlFmGBauPZhEH5l3LrjOXFaK1Vms9/tgf86QvoROr3FYV7ep94WSqJwz2
AlM6MGSpnP5ooe1dZnthZKxFJoBLKdSCsnUvefmqsWBPJEGgHOW9+9izdCoIg8HA
LHNpnUrHsK8tzWvI84t+1ixwqTRzMTMRvvrHbaUVzTLnIrA5cylp9bohcA3QZtWy
NI5iffcMMJMDXIoxIjwHaJOfvNicnFbRHvuxZx73SQzwYNbaQIvxgWz9KGe1BtYn
o42XFOniBgA41ReXGeun7INYG29f1ebidw3j8CNyFVcbvjJ6tHTvVW0wnR1E0m++
GFuokaP4SXQBlyInPNy2qOcIOzYDqdMxcgOoWav3oV8kqpEmOVJ9qTKbuik+AtIt
QzCEx03WqJPPZQbEylMvn5HYZAZfrizLj+5H8WTTTcW/C7dmRXzoN5xPwKMaSAxo
H1Vzn7LRqyztWh7yjglHSyt4mqK28VQu/CY3r1p6JSmRhRoT4Eaian2ddBHp09YS
134oz4v5IPK9RCR0a8x+4ajTT0vkGgdBbGNcgQvIpVhTTa94VSOhMUVn44208HB1
U5w772s9JtN6HfkzmUfP3/GhkqrriLvozqyKnjqUzhKUH5lUwycWbUQJsqRd5Rbp
8iBfaiNZkHXa37Lj/Ock9fgwEKG0l3q0IYusU5kuEjNkDfmBPixoGJ3DxkH5ftY7
NGMtvIqgE3OiPYQtkS2DdzsLG0tUInhfnFwgUNGpP6Uits6vzf0pHIgDm61RHSVX
0xqYH0JeVzb71rxgp9PzD5gQFjFbH5XhEN/8San6GBYJUzArZWIAgCsWuFe0FpcF
0PEU8IIKRid/cGzVWGX76XiNQN+XacXRxWDrdMhMF4uYW1rJJu1/hRVJRWkHNLIY
ZJTQesFrU/Nb6mw3SLcJQ5wYQUoP9kVMAvUqATuAZlxHoYANB5w8g1SqRXK8hogt
CUuDU1j11ohtXIik3iP2xjKIR7Z4pj8kVrVvantR8dICxICP6bJ/095iZ1t+AfjY
2nsCL+x3PfVkk6hdmWiRK0d9zY4GgYdNgMcWrC8SuYGRTHHrLQhQl2wVsSVSsU5g
cN3Uw+wgd1QXhUq3XUZmGjdEoR6E7PA9XBxHdXtc+fz+0fV3l7TeVpZKuoZEBz10
aa00M076cheTxh1nu7Nz24qWYYkWbBEWJ0lZCUe27TVFI68b5M6tCkeJ5uxhSGM0
8rtrdhFqAFfvKuhu0BaYB2PhC8yRUXBShjLD/LquOKF4yimzJyMbtCcXepc2Wkwh
e2Hwgthz26J2PCul3XRo9nyo+jvw77YlL3hTKxrD80Muu3uztZU9QzeeYq1t31tA
MTvuMZb1cl6gXpJNTtlBh6MybSkgGsP85GZ3oQm0gQQfKpJpD1kYZhQYeVgLT64h
HfDGnvoD+UBMpYJ1E9hYNoctO3bUKAO5K53sqnh/PqQVyxYq1tWoXMXGwrhHH59Q
eEPi5Ao10N+i6O3f0hsFZcdDpUGRWl7vI1eziOg9PvbgCr2WQoZQ7FUEPFCQtbDH
4G5MOb8MRWHlOdz5DCIQdk4zi0PwW+vOvJWUHNdjojEk4uPL9m4cjjD/wVLsvyKo
lxS1qKikOMYYZlerT1BnT4K4Lihh43mF9eLOh7l+kcfu8GqrjCiJSzA85XjmzIHm
RmcV8bHtMZxQ7685pvP14OpbW9s1T/8WZprbQag0p6RMazQJS/OOQufChUmrbo3/
jL/XtWkF/FUu9uTqW5T6lf3h0JBmTTD+bHd9OG2mce7VdF+FnbaI1lrf+wtNgie3
DoCaOQvlk3qYggzj3KKCexo9JX4nFVzJGU8PHY2YMiy9VX/0o+xyxD88T5j4/wa0
b2dOwwZCY7q+JyL0JH0xnTt/bsuWRYA4rWgdeBoM0DJJBljZCMkAxKeUcVYvvzke
lsFaeNmomsBk0P7899b8ryIWKnnmvJmnFyVSFiuK69bJc2NRNUtoc2zq+eckANri
PNah8N11oU9S5MqPUuByXjC4zmVhFtZllRHS2SGDNRUnoqXUxKEEq9/LL7Cvi42K
UUXIFkumdOhgu2oVsRtaU7PaQhAOIY+VsV/5XZtC6Jmy2x0ZP4dcfBWz5/2eBds8
6iL/PwpzkP/7j975nRWr6vBkoeZQoa/2pA9oNpD2m67u8Ds0mihP99FqwSkfXb9K
S6hkf6Mn8f/BdU7qffgUVB7L9iH3VHYglX1F9yUVDCGALfzrKNClh8jAP6Wa3PPj
cqM1C23Gy5apvOMCfJuFxDOnEpRUfPDmYhwi4ZL3MiCyAg1cs3PwC5sIoRX8LQoa
9PpNBs7aqgHcAQPx/nQuevxuyP/lL7OpdLVrCENJItl2iDS1EOkCRq63cXefVx/3
6M4FHhH9aJhc+Nl6pOK5gFqcSXpCL4bvFc0MbrBuyc4ORx6iKY3JLllUwPebk8KH
/h93va9c64QgCw0NX45gmol/3WUSHcMsfJV5naBkCNyfE70kfEx2dVSksFBRxJfp
Z3SzaZbOgG+jJhdNZtVqivlUr9C6gvrBDZxWdE/cGKZiOY0P4I9GRSSaK9vcMbOB
yN8IGVnu7HjxFDziMW0+j7Z+66l6gzXl9j+RsiiH7qssdlNax0A/1QAia7PN3+kJ
vYVLCs7zuaGtTzCjtrhC0p6QIwPFCeO8onbOYfYjwZFUikG8/Ud5w5HBlUck8GD0
CKiwHvH+TC5DWImqXOTOWQ9no7p4pkpArXkGOEhLB76oNEXKtoZ6BfHTzwW5uG4m
dhH8v8/YvmxzcQu/n9bxyyRMWsHWe0vwPKScnFP74e5ydqhtsfB6ER63a7kyI0LJ
6EzQgUDyvSBMlbQvYbhX8ZnJvMGQK12fTt8+ykjWcoqWGG5QlPGPh+8D9LBY52r6
E6ch1UrmUU/U1ws69zLqrLzG3Ioe3Xu7px6lgqRbeN8tvOqXgzMW6wTdUrL0E0jZ
+xuaZHl8hfAdg+J7Xj+/YbcDiD/mB796rJfQw687MwCALhckeNYdkgB39UISinYV
gdgBywxDWnEXxs05V+vVinoQU7W/kvv+OTSrTXFT15pgxsGYIAnE87WE7iqsC3+H
cXW+1Rz6eeNY0uU9pg/QAeZTzeIVQ7RNAPzVwxkOgKEkXVXVTCn4Oog38WeY7Q3l
tVC7Lnzgo/1x4CeFoRVd7B/bqLcb5C3VHeMtOt5tXVNuHlAJutBmD+lGiKncFJ4C
JDAzqsbwIHgtxw72tEZ4MRt05OHqDRukSIlouQ0fZm63k0vA0R706Q/gWLmlDI8G
8jCJuhkEYjwW5uRXEpsDBAVJbYFD+xYERM8hc70YDDBdNCWbSKycOpqxqVUsK0HJ
gqhFJ9JDmGtUGWxtbLnDb/BeYG9N0607aeJ5M6qNXnD8sMBvHZRBhro8Wjjv7shh
HC1OofUjh0GZSfOgkD+XAETGmImZcnjedBxTofscArOUgDC/FpBYZzlV2lN9Kyuj
rjf+ma6KIMrcXambPCbr6eosu1mYcDC9Vji2nleG4KtDVfNPo5qPY2GwDSElqRU4
cLizsj7asNUVe8qNy487kC88Ox0+2OxLnsOzjCh0p5znyX6S37HXzVtdr26ID5OX
OasBY88GrgpbnNxNFVxx7WeiPkoWvO/F6wQ5Gsjo6IvbvDk2K/kC4TvIH2f5XJPJ
XzOY4qhOb+btnZvinCAOGLyHhN/DpG1vNV0Kzrr+YCMNv0yGxzO+CZ3oj4+xVg0N
TMo9tbTdIkROXIFSOrpFPD56UsNtMD2V4va8ndsETV6TM+FOc21wE5x1kfRraSK+
tx+AnZSMbwcutMw4p0gna2Stv08p40XKiJGD2w2U4ejAPv7Py8wQJy3rnqb0edhG
YydV3Zer2vHWv6dL3sI4wtlFHbqLL+6zKUusm9E05B0XfgalSv0l7siBZIIwkEC+
59wb0N5Vb/CW0Dp29vh/+YdA1ZxHKJPPhO326s6PydNkHEJqq52kjb+MInrOYdrQ
PnjtMCrsE/LvC2uAGryIJyq3PgfR/l0ifHysEMu8fV4O23/5EXO4rWneNE4Y9QTF
voLbkX84+YnMJ/BEor+Wway1tQTEhhNmgHQmkrI5jTurJCMr8GsH9+9eCx4vayXr
ooVzDbGe+nq2/mhHEF1J5UIxGhZ+y7zjJviIKEQwaHxVxauSsj7G7r1mA1Mly0jz
jDW1crGsb02TSB5aRXlt0AGgmBtowmneWrxPh4BNGWrp0PN29CZlDRellMx91kXv
uklvNZGcK9qtGID1cFFIwRW54nvj80iESNetMkm3hyhhFWGK6J85J62vi1FOPtYr
YQoojtkbdfTFbdU5evmSKC+njUQH2glnS7+cKp3ImE1dJ7CZ5mXfzd4YHV2CDT91
sF7FRedJKwJC+nSPHtMjBjLsaFyR7G7tRJEiNSEqraS3d/MlvlwNZpFy0XEN6Ck7
NnhAqgU8X0pd0LvNq/D58z4vTf0GeAUUjnJ9alKczw8/AVH/bizxGaTFxXGmd/hN
kVrCxbyypSSNSfEr1PXmBo2NuY1ipLpY68kMJ8k+ah1e1xyU8wbos0GeNyvd6AZx
r6JsPY9N5buC4wtXa+bMo8pRg6PrHPJIksBBm1wfkjZvryDgfIfbE113P3/yh4+w
DZQpEQrEsv/CwwkxKtf4RkFR81waIJ/bU/dFGDoXfCl+uHB9UyK9CS2dQr28Mry+
P7jxli6alachfz/ByZpSEbOc0WXw/OWAZ0WmbpTscy3ud3IsYnNvxkeXZu30z/Vn
mUJl8sCbKNFrVfP9TTvQKckBzhAPEZrPHZ0woK8/R6uwe6Y3Y+blY7p0hCJuVzvO
9+C/9i8ClAvQwUwsjBSMi4nHT5CU+nrwir0IgfPkOhKomI17Y8aS0xc+UgRhEiHS
dg2/gAm44rKt02YOt9+NP52+Ve5qLq3l2WaAhHfR6a+oA+mX73MKypC/YvDeZ97g
4QPD7UzFy4qqP0LU6ug4RpT/DVCYAZRI/lkkU2DUDqtLZpkZ5XQknBRAFoc0gIFU
4/Plbx6TxTpsZmk9KpzzUqKXb1vjsyEyglN1WfkfLFKUkkiWjUeLF+rcaXmXze9Q
pPur3rUgxdHPFXGVEbHxkLS5RkOTWpnwJDeIG3pyMIX0I775yQImqdJl3GVrme2c
fpkerBSu1o5n3CyJSCjyjzv71aPmq4mWj1C6GbtdKii3K3W62W8AHTA3t8bL2KSB
eFSgED6HmPxHkuMMdc6F2DzGjDP7D554ElYfJcHKaozKWcaIdbeVIJPrsvSVtlBa
nKpvo49dQN6Yj1RZkklc9RAdeyFABk6bBQHROKoMiWtevUUTr3zUXLzwXQCyMVSc
XPu67TrUq6gqwAF6exgHQhXCVXGe8JGWXJSBJeCaeUX+UHWBurJlIxGnqbyWRh84
597ooADFSJVTeb6KiKdGyfZaLmFTnEhy4D7R6eha/o+7GQ46E/Y9Cn3MV5IVGBYo
GPf07yH3AonO/WcBeOjXd1qoMb/yYtgEcnuSoow/e9pCiTrZoqvDmZgTLaOCbTQO
zpBls9dwP1YeowTnVqUwR/MmqtbKDwo1cjBDWWxQPYRLjxhvgNFQ4YwhdbXLL+pN
HMX32zaSR0NP6HvVQeO3WESWJhogCDwvH8ao4+R/m2otiNmUAnCQoTysTChunOnN
YNC9RaLWLPyF+SNK1bbqQe7lBZTMXHQKAJKE4dsVuKFCuiK7snCoFBBK3EGAdurd
niWuXzQg4gp9gk+VC2oOD7R8Mn6las0/Znrd0HK+GpgLOBjh9emXySQQTVm6Q++B
eGtpwC5wGBfRE60WcETuXbcETqcE6U62MhNKrADlDdZCJulg+Apnt0mPuFWY8lQd
zQlxz+BEyJhQsPGhBR8q7fI18Khl0FaOptnI+xpZ8rXAA1eJz62pwheU01fJS+Fj
o/87NLiCYvewJq8IwBsdVWxM7Ey5KLYDUX3P3sYRfYlNBb0+pBKbsURdgblyialE
zzELRmqR9DcHUvPyzhneW2c66Eb+LtDCT4rh2BJriPTYiugyFLFvyk+pHu/CGdlD
xui7h9YFypmeNV2fyabWBSiNxLcf6jMpC9a74f9WfF0haqEQ0f02UARHKVncpFup
RafiVOrF7iyb7dmK35BatvgkS0NSV7bmY5GtCPiVatambs/rk4u4/e+btUSWsvD+
qJoxyxAIbI983E4lPExQRM+Qv4FpY56aXCbsT3ES2W82zr6WWmMOyxkLLAhbtVGD
MlkoKG+vmDA+GyZGjBBHH+lJ2gfHWzU5b3i3lOn5bJJpV7p/QQEnQ9xokhLfbrcl
F9lCo29YVHPJyn/6MwowrPS2LjvcgojDPud/T23dzxAKiaMJJHox97MXuRHDs00U
SQWgzbj7OGzx1YNl94TgYF8QTMschqhrUYvOyZP+TuQIku5RX7Ghm4tWoJo5Xteo
7Avf4slmbywcsYC2WY7NUe4oaZilWPBaBifKjZCw8DTSQlbKxBPFjaTpG7TmaT53
PrW475SKSt264gSh4XWxAz/S1RGpH3BIeDoXAHIXMg6gzSAilFAMpgYuJ/gCvmos
HC+hxQ4gctmUmFJvzJ5UdS7d1ubi4iU1CMciZAsmlvfl+I72m87M92JUt9gwBSJJ
gDQt1jaBpWtAQCIo4djyW0paM8l3FVotvnXdCah0YrFQMZs2rsrwxJgyMkUzWlHA
wVbSr7PqKEknSu0dngyGOqhiZXTbTczPzOj2pa1TY80FvPucVdVdSTPWsazz/yZj
pc7wB/5ECB+7Nu9iNGarIvvEKSUsHNFM/kEtTK8nLEKvFv0TDv4pXRB6Xo+yjlFR
/q1cco6cGt0XBDf34iDQyHH40IJ7UdNK57xhcBBV/OEfHI2WMD4uqZpAfRbqouEL
US9NEbdnz3QAmgSF/xtxbfn/QCbR873aksoXJl7eq0KXVFpEg2cpUkVR74POn0gC
GQlATrEbMTehiupUP1ynEehsc+P3uOS2kYBr5fVwD+rgG/4YACJQBzyLH7Sf0sM4
4Sev4/K7sRU1168xvgdMLamRImPlgD9U5v2qQtuymAaz5m4a8Y0JAwqTUfKTb484
tmaSHDsQ1AIhTYk0W/3tkVcYHANQ8myMibHCoGmybyXsCGvmhqaQkJaYzbxNU+uN
J2gtrxSeFU3J1kWiNf71dkmiDBDnT4C3yjP88B+a2lxS5WCl1N/W1VEREoxpZJEe
EzKnaZWkCDdD0uMHIvSJnSXEoqnIy0ZaY2TIg4dQrLI//FLAyq4ihAlOIGHRksiS
IJGiPSsMogOD5uAp4xezs0apZeVZHBlADK1FMGhVbcdIBvV/sOM32vGhr8SdZud8
6J7PluQoPZlBvPQ0Jam/05etOaMnWWS5Juk1golIQIjOzMKZNw8gzc+0yp9fhNMN
40vtgsBgcLj50cM9ie7l1wdd5FzOatue9dnQ281231Cdyn7iPZVtfA6OC7r1EF+K
nKX7Y2wFKsh+/Ol1rMu73VOsHyyyORSfyNvyIaNCwHPDHK3v2vdKW5t60fBasnMe
Ekck77g8urKKtohCFKEl4HIZ/p0rtgLLPfFRNlvp8fuLCBhq8JLq/EyMaVQgJSf1
pC/I4hT6+krcLC3kpV+Iupk+qUwIBWxzXEL4/qJaCtKhI4L5DtJLo9vWOvtLg/6m
HUbKZ6/jM6yZavJOKdTCeW/Zy66nH6gDEfm6ejR9HjvbO4zpj5NZDWMGxIe8FdFT
k21IA2fHgDZYiTnQORX+Ptxc9q3dDQPWjyscOpK2lQQxCyc55amgHL3iqwIn2ILN
U7SGYODmTjD+XL/GixYGUMJnWlR7FzeAHq2pOyLggHXeCq7yCAy/KCxDk3hFjB2U
FIgfKiESrOaitLd3kANZdQ0SL2JVHJH7sKqHr8ecFgX30QFUgiiTo7B8809FLd/8
xoNJVWZlvg99JvGHUGCTEgdphI6M5Q+ddbBeR51AXT/ntDwEqYejHQXXsX31WG7/
jeR9Gu4s1T2WnSTVXHbT+tGT1nXccabcKo7mgAy2YyZwSHynu0O4FebeFSNA1F99
jMpIaHNEt9JDoMDQz7AZMXcadvTk4T42M2b/gtyHMUL4oXloDsPsjnf4Fjm6e+/8
6JK61RHchcQeZek12pOcS2I/HnaK2GAw2yXva5D54yn7f6sjfkxvKcqlDkWXzFwW
W7w619dehjBVtUmhtMYJEIAn8bFFlAQ2d89UbPG+Ff/AEfQ0CAOZ+wk6onWuIUYp
cJ1k5UrXOsq3c9y6+b9+ATBiHb4anfm2GT2kOjqba4M8d0fQlx6MN6n47vx2ElTp
Mm8tV1Xqe4ZLCO1KcMzuZsSFa9VC3E+0Jy83/byv5PoCWbk1LrXvNLUNSGfjgzfx
0V5XQmfXyUjPoHtJTANjyS53VBzpxmNbPApltuIrm390isjL1+9eFy9aVHs7wZry
BEWmgnCLEJTopSZZESo+rcuLQ634ffoVy7gu3oA1+xAOAzyb3cNaWLR0+c0KpPCD
w4TawNdhEGglGYg2kixuHx5x4RDWJ2WUm5XfmBuZxmaV0e2etIPpXfsU2r9ZLS4V
vNds5zoior58k8sjCwDsJMexUyDOTRFdnCbs2Gggi04ybhVGsrw4p4xd05phkbin
t44TXxHD5UCygg01LkjYykBM8DjujgA9OFBe7/GmQuzd5qrYu8qTxA/zDrzF6FSQ
CBetuINSqz87x2pDYNeqFD5pqWLlkwVr56T3g/FYgnV+HGObYpdZ2Sqqrz+5fDeK
xD2pbCEUbr9WmBLVhiAGCX5anevpVaHvfkMck9J1Tx4jZ9PS7U6t30UYrMGfdsek
QE+TuvOM0/WCQj/K2H19i2fDW13vM6wjIMPHr8ZwN0mvZqGsHLvvV6wZHNvfbO7v
sbJ54a0Ebka7LLolEhxcf2qCIi/+AsB6ej6s69PxFTTtPg4GYzIYAoa8y7zuJ6pM
39kp+LscHSRYhsFDE7j/0PO+T9B1diOz97aTAjqg8dzBFQeOqbsXzfAITfyckvIr
/D4ojaDo+6zh+TCo67uZhZnDK6MUuEv355u5mLpWayhdy9OiBxM7WGdybSyKsQ6+
gvgu7gBvAPYJzJHdLmvHmOjvWrrAlXW8BdffSYtm0uo+62zGhRQ6X3schFtZMMUl
Sli8Pwj3hKtzGrn0wozHzil9zK1TDwphya7uVGjMa1yY1cQqjpr3QOHq//LfVe3E
B1ne7HC54L2Di2HpSPrdLzATpjsISDfWXsxfvjGSPhVjY8eUs8jkLv2Vh9hHly/0
5dTBYJLp4teN2AXXVApk70UK5ATDsPwteUn+MdTdt2RpsU0tXtJtjBYywUQCOJWH
uGZA7Nvn0ta71DRk5hnuReqMCphDOKE1+icwxttyErXnnMuG2co1db2iTX2P0the
U/jAAeKcgk0v8+qPEQburixNRvYBNJyDrUN600M9KJ4Hxx/8y9eOHGHbzWTlOgxc
uCV5yihXN0j1HJNwv4VfIOub2VPE+iuTUSaqvf17zLJ/vYwkDUoGx7BTC2h9TtUn
+NUvuf8cwDSYWdYpUyxR3g+AtUF7MuHfJmfhhwZWJY+kSjalhGBQKhnXIJ2plb9t
+qKXTx0kzg+6RAjGxuPYigOeaonelBYzD5T2oO2kOCpCiuscSSVaBAcBJ1ftnTvK
rkrUPwI2QHuVr9e+Q/feQQJjunoJjetsipWfp4J5s38suqr0IjlCd5Buhimkw9PS
uyT/tzYZtHIRmmDD6hRtIs+5FjKzJNLbWWg7GlTRMR365FoHJ25eWjBVOe733MgU
h8FceIm55/Ou7zc+VLGoFdZBvpshhWqZz4L2kHmF5y7rWI5SnWCb7LEwQPp1hmru
TAomPIeIGmNjCggyArhnAz8Osj+VMl2illr39FlTLxQ1BiDpmACKhH/MmYVuNya6
eLFjegn0gN50H2e2cW3Cd6tQ27SaGploTzvrT7p2JfkEJnO16Vh1ypAavdjLd3Gw
bABeWgUqvUr27ZJ5Oce32cQkUGYtzMAcPDEsFupeheWpQ6JYOaPhwhr1o1ydZ3YZ
XBvX0RmatlapGwo5ZXokIS0DbFG6dswSm9Cnp7W9VdVQG2XZEoBrvhgM0q5GOr3t
mMCGbZ0yS9dV46Uwt7TH74GqbQuS9l2vV5KG1dVAWC+hJRC5DyqT2HHTbkQWZjLD
ROiv94lZPdlbOsqImvZm+Xil72ErmnEtoYXfyZGRuoYboyTph50PtQt/okkOZsY5
CLryfuCS5t6NhX3R0iET4jx+wo07rg4+xeKivfhXsZE0I48OV3lbNsFC1wVZE8HI
2T1Zc6MPeUlW/Hn3QgIIMG7fDGlpgnkUR71LapC1BkzcVlbaYe9Ct0Hr3EZPgRnB
QysU5UGuK/Iytn2i8I54pMryM5ShEHRxZzICbI/Zy8gH8U3vHFuG13QQslUw1QLZ
sBjL9WOR+zKS05BHbxRHMmJ9ujilon8hjIyFIHR9/49lL0KlOcAI4N5FGAC+1f7x
CfMGYQl0df7CjgNNmCvAAXxVUWThftI/v3158YM2KewTbJALplJsQZ2ufClCTXGj
o8YDpM5MhNAxZERs54u+5W6rjWAB8Gx1uNQO4m/QxtttPCvqgVr2e10BLTOxBpp/
YXAIhQsJAMYRqZNAWQOtFmwtkUdsyUTVttLB1OIB2UPgNiwXbacepMqYV0s/Qk8Y
0aSd/aVQrFb08PEd41ZaWMsmOAWsvmluMQKLnIjJ1aOjSmesNZxvK2AVFQfzc1Fg
o+NLgHveaHK3YHYeEBpfZ0VDAUX5JRbMeqhOnBz3AAoObPlE8T5toQOn+bj10fOF
oQlzp/zjiyz8MmBr5Ivqs6SV9oC3Lvo6sUfCO0SynQ2GD8Bst34Pi6kNgoddXJLz
RbNQAgxiz4AmgXHgWmUBis6WDf5DhA4wcvaszP5x1U0o2tY9cC6xQpLU9yBb1xy9
CfQhzmqQJYwjAfCQEa0MmYw3BaeLXsqa8sImg8BoGFDzAPGymrUcRAdaOtggCkyT
hBzfScWKYDe3cBc2rEBi8SoR9Rj5lmxCeK/UZWDzp9sY+jF7AQjc3xq4mGjHCOXQ
LEsAYbBhwEMS2tEuvdvroZ7FdqOhnmCBiNh2D13nzziwfeSOFTHW7qDMh3wQJHki
os99Jmj31mXqNWyGiMf18vIo54istuGWDm1L7w63leYgEDQy8PQVVmpZ/Mwj11uN
eDxGyuoJtLBtLUFUjGdK8sJ8BlT5NfNuwESRCoSZUIseLE3kUAmTVMxU4HQ4mGet
M6cSVZPVXulYXYnvpzKnRANT0GMoGokt6jIwgSqJvx/RD29uIH8NyqsxUsF/Wn2N
IJIJWyPYrlY5dQDsG4ZtGMgkZDXCRPT5tKsu/biOTIILSRqlEQ8fctuDZK3k5+pW
GUPqkbwS3z3nviIV2csjNSKtgVtMXt81iAJ7zwvjZuhiQ0NKIk+Alxba+RgBsczs
hKVjcwG8hAvxlU5OUuMxssLmef2Gdec5ZfbKM4IqHnxbNLtxi5uJIk5M/dl9Wly9
+jP4x1qjx1HpN3B7k2tyzxJTeyZgU+Z+e1fKA/2yF0mTezXWXR3qsZEYhIzlNiF9
H4ZNLFIR0J3MIQe4fEqBUwX8h3zcbiJTjTS1Zm1YLjr1HIuIYpu8+rkHNlIt7Mg7
q3qZFZTKVLqR7pu5BGcyiD9ZqP4gwNfQLhxgxyI6oGlXp2H+mxHFrjufeyplN9O0
Ci51ThiEDpQtFEl4UwxYHqK7OSDWIsi2eHXa8sl1HughCumdcAr6rqbf39Omb4dd
r5EBnf1J/nij1Y639IC+bJztYH/KgBzC8IjKnlFTtRpEQTTxZjbdAfEwTtd6bJud
KuDk5Bo49eWzpui6LOF3UjK6/saewwafROu7WS2JCeZ3Q7jvZbEcTN+mdEOqRaHg
z3giskJS3Hx9YL0wEy1KSpmadjkSKYKTVi/XCESKcLLeus1OAX+NFzCEZ4SZycoR
Eo8zce3pAs/Nhd5d8vfqK2ah6AbGROOFJfJIrasl2hEmm8BIEv6BFYvuIRCvJgyv
dHnwh8Znts1GLfBLuGNdFWfsYjmy1FK5fuuGurVKJ4kTR49B7zUkQBRXuL9Ar7ky
vSIhVqQD/CkfRpfhvpBSzWICSoVcTMGCi3PPRIG70UCbnbJpBcEw79Q4NdPWksVU
ALyU4JcMOhEz++pOoD6ipvofX4bYUxZWjQIg/J7dUsI6u12eaaV4TSgXKMbtglPL
g+p4roQqdWdyLWKp58tcR5xs6AP2xv5npZZ7ODYS9DsDFbn0ZI6apcb3f0fRit6K
yJ0rDpSA+duquHlAQZzS19XMX0lJ5ja3BR1kwvywtVSL67QCsBydelFbYeD7Uwnt
piCG+Xy3VXZmGtlOIHnaf/Lp2onDsJKqJXVY2AR1bsI5YyhJKcSGRxBk+rABh2EK
+rfcQoSLAqED/J9C4yr1fRA0MCBU8n19J1dZVUodvP+JYSKUEmErB8Ew45munmuU
CSaY2ZUiP6AolWQTbj3u+/QUjQXqatCuIaz5LxAzXUyK8hq4c58G0H4JMhey7wN3
lARnUWC+T5iseTvH7mwHQujpb+11nwUNsB6JJIjrOlcM4aFLuWDQEwmHFqMTHbde
E5PPzAVS5DEsC4SfKkFXylO16ynh7dspYOLIE3cIKBZ56XN+qSYq1rOZM/tZDVrP
rXuCFERRUrtHUzOHxUnWp8abfl6Cx8NBPdGzewmyUhuaEiP1iodOb6XLuVW9iZTy
YKsYvDuLLSpRmKm0D77tScAew1BDr3wjZQ34LObmP27Zpctpfyg5Q+tkOZqhSTV0
sSRGIGyD/Zxa4j3nu+anr92Xr4z8eD5yd0ugt4aZgsOwSTxFbVHdwWdpYt8YOAaU
wzsAjveFCWQ5l250ctwujpPUDcZy1zOOw+hqzAyzu5bCOAPt/L54yGH4H6VAZlz1
VLntRRHv+6AMDwmUeBsRa1WrtDCjkEwVUJriU4oOC34hunoIL6MTBd50DHRZfqNF
A3yew/zWs0Ty5Jsx3PaDPk48TRv/bmUbZ1blJjSsrlEZMGdMN/NhzHb1BHD15vph
zIoRtGvJdnJaT1TGdkCKpY6yO8zH7Bwl/tm1SmoG5SfQBMxn7Aar7Ea5qZesG1dq
zgOLW+oTT9/qB0WtM2KCrcNQDNS8RqqggE7UUzG3QrJmvhO5Lls8+djQcvQZvC0D
IBQ+tRsKCjGrkPTaxWPvy48B+VUYpkVYr9tlTzzBxy2H/sTo+vF7GrXCM31aY9L9
pOorVGtsOE8UThEtXsBVKJ2MnvgrD+f7pjsaRZbDIGbPItEHPrFSZ021gq7PhG8Y
7zq8V9WJvYEI1b99N4O52hKyMd9ZqWINVUinVC7LBUfFW7g7o0REs+z55ttvumcT
5DL+OHiJaNYl9Grq2/Ll2UnJvweKBh2s67yA2rn6xpzuEm+7TOBD8oX+MVcWb7sQ
Ki/q+SBMqNPk7QT4+ugL9PEbuAoQlVlx5AYYKai/5TfwE4eim+iDW6RJkE2buV41
E7LQTWI95bo1nuTV4+QaPnw5O3xtf0GTmsxEPhBSft3h5TfWA2a0pmmzxGVO+5Ij
nd3T8HZQigW6YQ2c1Qy7eLQbr8YBK8UPEZ1EAX4363WJVmLR8ZtxJHS+fl3eSbLJ
QVn7jvkdg1FOEQ2sUnBaGL25JfkfEJWAdiMrKAKaLLIZNW++Qcyu9DZ19c5QuLlH
LZOdKe+h7PkrEit78MUoxTEJINvJ1prcuF18ePx93u0XCY/piLqMtT6P35DhAQaF
lbZEOP+Q4GjVhcWGgfy1E7PmcxIkVds3VLzVevHIjfsUiGUm/gSBpS81SV61LEK1
Tdno28P5x+Qcx8EeIfPgfzheb/Uvj3SQJwfKSZmXn8yjOUtjBo3gf3JAHKMUs3cH
yshwy5T6/RFgL7YA2KMGBk4qj0RPjgnZvcqOOm0qxQ/ADs03SAw4DKLJpAxjRse7
CpYzh3wyDOQqngpJtiAB9Lks1p1J2uDb7BWlPvmsDyqjQ70u2h2X8cdjKHnTIuGh
jUc5XngWOIyoSZ/h2uhFmm2vyoAg5FoU8ZaRcuZj+0Zm5XzoWSEogGWpPjxsY8e+
JNx6zVqwJaDLcpI03zwALVv4vnYZBNkrZ50/yx/ePqwH3LmCZLZn9qYwwepoODPe
f2nQbtKtIxnfAh78hAXcqhc6K0ODhSKpbm2uxHHQhy3pZCarkIM1yLDF5qkCk9wz
gA092ILVpAO5LmH2q+ubmiJZ2eZ4oLH4gLCs//zvT5/p5RVm19VxDL/Sp3DuRz85
SmTNXnzduQmfkoJ5YYyQmtTODip+ay7Bq4wqdq+D0EDS8NmEa5bPmcX80YPGrssL
DJAztWTe9dz+xeCD/gdVLHOychpoDpcFm/zGfICcivqlJvbPcdxDBtK9OACSZyA2
KOGjP3ltzLlf0vIhHe5C9BXHjjg9FLkGFaZC8rEVFS4=
`pragma protect end_protected
