// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:37:08 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hiRPtDD3o66y2sAiHn3m8XeUEOyvd1Y/rMVLvKpf5nllFhCJbDt/v4K/+XWtP/jX
FTn64vjx6GKVhLBH47IbVHxh7HZTeZB5NwGCJ2mbsYftDz/kDWE1nq039FKstofl
9igStm/HUYkQb/F4TTo+DqMFO5XZ8a2bLdI//zyfZTk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10256)
MRq0+6nMza22OKdlPaACGzd4Dfu+aXukxosYSR5CQPWnbCzFOvTZxtpLiGCUUQKd
XNwh4naIp+Fb2fKj18QlWg37EuqSwBGtIvbUN/XZO3qfESPPDaefX3uem6fKtS8D
A9LCwmhdkP2T+jsv+MY2DvFppFQ/edfOjh/p5IOmh4hMylxYFWjsq2vqy/wurrtD
FPDdfvl56KxjfniCCYmTDUkx2pe2r01UDChKQxJADw9ZPbLu/fDoMAMdKhK62x4z
49uSDWOeCKOWVt/xjRzv5Wk211e1BqDHDg+g2zs8VHEi7hD2OVeaW6TGPkYZgIrB
xTVTijZFSjGWSsAIJg39vWNXIrt6v8rDwLGmaYSh2x/w7EyvwEe2Yd4DUB6V8vvx
Grf3b23z/fJq3eb7T0s1pJBkbi6fufz8iJL0tknlrS8pDFbByZKslkxvqgVgJagw
s5zNSi9onDxt3YPTEQHM/rw6ItqzaHAxe+Umc2LI0S3HCErL2kkmg1OmAEtB/fRN
AQKitprRQu9zwAMGuXBpD6FbypVov1dPVxFmEvZrOREfVaOMBVsJ/rDVSpARVh53
FQ77KZ2mvGZqB64Qx8cqf9ZQdY0FExXPakYLyZPYyZUw7oB07ETPAQPorxxRh0Px
a0XwyRcqhNfCJdl2umikRvStMxXztRKtZI5+adVYyHpwwSL30sD1k2AAAH31uLJF
/BD2hxO3NpFkIlCvSG8ENM+7OPFV9T+JvAJv9aq1B4VppdhCL/8pLPujKf7XAF5B
+/FUXKDf13ToDoBI6ZohOtnxnwVZljxJcZBPno99G32+Cnx0p9kp7X9/3Xz8iGco
P+N+DR9DsjIMKQpodPgd0wJqvKnPgFXt4beLnEKqSiHW3aS8HkM/kftY4D1lQZWL
2cmP/FFCZ71noM28KKajkP2eD5pJTBwUVE0e8S9GCY8b9CZtEnVAXNymwtnj6lrh
p85wMf2F2GQjn1oX05dSKrfi9VMwvZIp6JouAaCPvoP5EJ+rETWQ6CCpXaRzLyJn
DicAjEjWQkjw/3BFFeLRyvnR6kfXQ62ALKpAoSPoC+lpRqzCgTzMaEenIjiZJNdB
E8vJkc1TOeO0o+NgadrB0qd3Vyyn2UFonacIcBzCETE5/Cu6FhLIwEj4g3s1Pm/L
bVfD7xP0Ojd+HPJWVAxFv5b83+CKUrk5yr1xMEqzep0aSnEToavtDgm9znAoltrs
GAeLjGIRRjpHnbne2ugeQdLKHtTTikPqZz0EK9hGi8cfo17f2xb27l0D5wbsmS23
VFY31t5BqKLHl2XgGea+d4+vZEHyXfdXv8yMY92B8sKhR8B+BDkdHVYuipPVhf28
Wr5aJuJCNkW/1dwEc49rEU63/vxkElZTGvmLMaqJbtJt41Qc6QXQwlDDJh6vn+Z/
nlvbEkuWOG2ceYsoXoLAKT8waOiTITFjUR/SGgOqZMiB4WkFX8k6yYixOoQrYHRv
Uy4BKirWsJ9zcvNYBILJqM+uF1klZVvRjUKLJ37XxOMaXkOfNBJdaSesVcXA5+Iy
HbhYrmZZSYZbIlMglyVIaLqCq4gzKcuBrtAovs4iz6A1qDCmDdsEcywnvqNNreYR
ItnwNVjp8vc9xDJFAAMQOGx7w0EAfi7T2CZN/GAYozORUUJwcO/h62irQWXXGGIL
nro78+Ea5SB1bM1tADEs2BkIgIzu7yI4RIBwMYfUdeIDnTz9gLR5qIXkA5e8rU4k
HMA1GNuKGZzyQ1aQRNLuJpM2ELT27TxwDC55i+IMo6cn2aypWOVczLWs87nkm1DQ
Zu52fC11h61vkQ36CwOWyawyzX2osj4Ao9P7YPwGQVSPLrPPkj49cRfqen5tryW/
w7/Q5b/JYHLjnq6WDUzXQyW+hFhYtvyKWjOu/ZTFeYjJWfDJUc9gaoyVM73wmk69
RBgPv3/x4ysyjqRASHEUfo3YQLcqZAcAQ4vxdCTEmNHTwtsV8L7dtgc4Js7cguSU
U6A0FVPP42nLwo05zbOKTroU8bxjb1vI6xTFJsQEBlOREijGJRcJ2HUIYwRYhK/u
f/uYL1I0apR3cB0xvvntAKuYC31S8Dh0aVYucv11ULsrqafEAInGv15fhkFd1KER
VMwPgUsk8isej+0KsVxcYaahLJ83c0i6fk41RCJhio1Jo0hny7GChT2RslKBf6u7
xF+LnXqeQavbDLv9g/jq/TsWrHjGAIKaPuJGfjJGcWph5IQnDDFrjANZzjugO0RM
xXo8iZ8XWI6YV1tDGA0el9q/lJugeJ8wPcA3vjCyoga/am7zs3ldPnyWiN+FB/W8
q9uBu+O6W/y1XiYuLtlLiXaMeH0uJO/Ic7rF32IOpbwV4sD/1OA0U8C8Hhe3N4OI
sUKP2UFiWFeGbPWDfh7ko4tpfLN1mu5OGcTAcamfDI2at+A4ebkv0yUUXrJxN5Gi
6WdWYiMIX3K5DbrhVUma9FtaXtfB+LYvFcYmFA9KVac/3Wu78E9C/BGTWLp1Fm2a
99c7N+35lgCLcz8px1fhbvNxn2AyV4Rd37+NQ13ibmTG+jjGY3czV1Zljf4ufh7d
UEYmALq6Eqn2W/98O3SKZ3mh4bKh+fV6UmucENeASel4oAHhVKXUELWQC6UV+DTf
5ujQ2VHm6omV9Kgo1NJYutXHZiNnHuqAuSzhzycxj6Dq2GQO9qNMRnWRrfFATEzO
0JGSVQbKc2EVKtLh8zAndmJHDcYS2k/QNJHezq3Y3Cw83FhbVDyFUvBuNKRypIP1
ImuTDod1x/2US22Yps2LSTNV0hOEtu0Ndu5etxVk4OH6GMvDA5VfyFyW8lQufVfB
RjIl3R72FBFg1OdKWqCABLnHAb1hmd4I5C0zO0+C506f4jaiQt8A9IZWOaIT3Gn8
q2fsuXfHS1nZn+sU2SogejJV2r2RlWRU/EPv5svQTxSQ1WvkYS4vXV0OkX22Blaq
VBVZ9xhXGf3ki3t+8tZjOvo1b2ZeacZi6yu+NUsqaz5J74G2h3QTRuUoS8LiJqTN
CBz/oZ2ymkaySe4G4v7YK+qzrN9NiS1pMif6pbZNJ+pk21zYTNE1URTlc/TfayfY
Xr6m2B/KBj69BFRrQFAUg4v2fHiIkrYNHbF9piy4MIY/uGIFOUHwCo+CQa9nT9zx
eRsNWBy8198lNJAKONOzUSXsif5eFZN9yN7TF88J90jEUWOtDwt3IHEB+sXttiVv
draIoF7pHZyz/iMPIWkhNWvLIcyIdQ/OqEewsbo0QjFmG1rpHFa11OJwB1sDXxLr
8N0fK2s/3YzqygjErCuaLdl/0mulKDjd2u0Zj44nthUNkLYLdCEeBN/FiUBTWOuB
fcrO/T07t+LredeuhL2OP4apkNoymQhXF8yeQ25qylsOot6Rek1OPdPvWkId9YZu
Eg2g8iEKH8NEDfRfSXJG+NrYjOAMaa5WRiY9ZHFsuXQ5KCt3dEUbS5ogG1UYPm93
ptPuLRmuWQ5jBb0eQN3YldlLKSxcHE5DVB/uVYTKN1r6Fon9VZ/3TQRLO5EU7NPv
ds2DMfuhuXM+o66KmPn9tymPtTLp6h523mNw84F6W7WbCtnB/vgrAFRX+JX7kvvI
wPvm0tXg5ce9SQ1Eco5fsBvdZvpVK4QKCbGOxXhvKo+U8mgNg7wTaqjh/tKfed6W
DLljQnm9+c6NqsFBGInsiCyW9mmh65QVjjIM3c2DKvoWJADyUQy8XI4/rud4vNff
VHj5Q//chm63G3U2d5ocNeZGFOWWetWc1g6/izVHdKexSWi0KEsugJtZEZ92Ep9w
dRLxt0PwgmNEIGD832bTTcPP92UMXXewMrNf6G8chvvDQDp7gEcv9U0K5IDwYJ1c
5TdiNnuti6D9HjKGh6aBFowT9/MiPkINfCVt2zAxfuq8d8ez+qwuyJF7p0efeCxn
2lSaZYZ2N7SIn5SWhvekDxviqNkYX6m4FonuRGCcCyK1cqmixEuU14xSOCqtQ9kk
NQS5VTWjTC6SoNvl+Il2rfze6jpOrYuNkh7WMZwQHcA0tCQk1qd2r0qJHoeLjBia
/Gtl6I7e98wBNMriHsnFFh8XaR4inCa/1MsfopYeHZ8XlRyhNMa73H5bcQAB0tE+
0diXthZS04EU7O1NIL7YM+nFoFBrvkj4Qe8h9q0FCAhSdeJA08jdQdYoLtIgja6x
4tY0UlhqEZPqQHcOx5m1Or1vHHOln1SiL/vQtCGTtZuHW0ORCUV9oCZp2puxXzBT
uj92CfwBlTsukOrVzQttHrhi1MZG+I2yXPO4pAWUjuMM+s3wMF6JvDWZ2m4DtUFp
5TvnvVK4s+hRjnQHlapBf/XrBA9jvZHRdbRyhNmLomZ5fTJukxd2Sk2suenSutPN
W4IoeSamfZaBjgtzxUVADP2bRAsjfjTEuB95C779Q7utXKOGoTBLJ3bT7RrkiXeK
mMhzlXRsLFMvAP7sfsMIwDprK0SyHhNzVUFi3DK8N2cwAlq7szIQyDvO6RFrBCD0
o+mNmt+UoqgwD97SEWMI291Hok2tvsGY2bECAuoLUF/y5dcchclSq+0/MNJQzXOV
EwGHIM3laY7xu8JhWkveIzFEUzlpu9Cl/fBHYuwEpVwP6XGpUa8aYlB0gA3fJz0w
Ov8z23merFfEa5UrK8mG4VPnebYkn2qghV1XjYANYY32PPL0NsBAfUi1Qc3z8+22
Q3qmZr3U9x1BxO6VWRibtkKU/4yza3P8fcI6yF/mPuz/rHh96imPk6I0Wj7mtLLC
Ye3hrDYx8H0fFQKMQFxLYVZF77r+IFdgk3cNEst7cr7GBJhYm3mZhFajSMahWtaW
axQgsfO+kU3wjmWrbBbDgM7JwJ7vQmAUIUi3jcM9HgjKVTaJH8QJs+xDJEWqhTPL
ka+gQNtjdoc6+B6CLJYjtDoOgBl4TZIyFAxHqX96qqrmXuFRc4GVgaKnliK0uIfa
Ev0dqY6YIeiUc5yEOHaH2mVQZ8PiOze1NI985lZWE6Fi/E2Jf7T6VxWwyeuguKOr
hqeVbAJMqGokdm/3MzmA0pMGh3LK8VAr2aCPZVMlWy3YKP90ANobxsj+AeZsDN56
8vhFTNfqLIx5KFDnxiyiQ2u/9D5zsJO7vyaLdR/iRt/cMc32IQ2r/K9KRr2INxPc
xu2iSt9I5ygplbR1Q5nJ7s8M6v1boaFc/0GYZgAo1//m19Y3ibPo7f7LeyEGEK5G
50g/M6wy0wCzBvqlO1b6AcdkiGJOqrhBXc6xSO/C9VOiIe4hsTztJrcgmpepR58T
F21R1HkEwB+61YLCAVMv8BhIej0HtELGvKXrkk0sMJoF9LlO6zXtZEXP82jun5Pz
PV0BsnPYLxGyhgFdR0tADGx1W4eTBop7QxZ6HM3XITIoD4+fMq2opuERiCQne78e
XUK4JxI21uc5ntbma7GzDFkKby7O1vCY1iQOHZnUWAlq4ZKJ9gAwaXVhDE043GS3
lS0X5MPiAa6b7PLI1CiXGddzGuCk+tlXKj88+3Jjr34X/e019pU6RtJJjvAv94WL
bQk4c5pGdfFQb1Lrxri6RODhNoCTJ+ZSzBuDjRcZns0ImYHsXN7/ov/CA79wViF/
Xfu5szge2bHKzT8Mcw3UJwBig2s3UJPU8WXbNAegyYhpgzJvD5iceexN+UDppOjS
Yaskix97RrZOn/k5DQOwqUFDk3xKlbRZzZ0xgH6eQ8I/GPvy3Q0mtTKDuONidPEH
RaE3U8UxiFGhMaNzzM/Bq/GsHPO3BQA0hZixO2rnoUN3wkJ2Z33HEYJv3xrMlDLg
I3EMUXfYlPAx+UDOJYxMGjVnS+y40e2059cVfrVu8en3h03bcXRl2byK7nFzVcdq
TpTTE/pFPzdPc19qaYAf3Qg7B6MXJbkEJGYmMLl5I63s/ql0Ej7nwK/N7UljVZEh
SRK+ACdu4sXk6urwczI3nqTeDpKtVQ8ZxJ4VWusu3WaJIzccAFkL/6y289FBl7F5
t75bL3n7wyfxz9o8sSCMFr+dRoOYmxD/T9DsuX2NgSUGM0hi3yQCren5XCZ18c4x
t2jP9nceUeUJfnwBWkGZC5veUMfRzam+mwaZ2rlQkjsvSUhgagr4xp6jZxmHil3V
cZFf//trVHungAfeIgX4HT8s928CcaZd2mdzoIQKenhoRl7bZlOnoEsayuBktwlK
aJHeqglAdN7P+9FS1rlGT2Dhck4L5bIDnMTNUdjxpCLj31R3bk13MzOLnLibXjIL
Ra1DqNGihn3PX7HndXpC/FMnRodhWHFU/OqIkvfOj64xD+iZqk/Vr1T1dUhU+qeq
fc8Xei1k2ZcycAGjhiYGehCXW/K2JEYWybYLV8RozrpzDf5840VAWdUxPt4Q63Sk
Tewq+dYkw2Aea9903H+SMoSEdh60bTJcHUUw6BUQ2GcWpRh6RzfqsJlIhFUdmMZN
XCUsA3zMxqvYovNi/sBB7VpE9KcMqkSqQp6r0jamb8k7YVjYAl+L5JloHoYt1h0A
wfC6sOW7EYvhRHRWm/ANY+eqNLRF2+KGkcZQF38OVEip+vT1Ax/EtOaJlLJlJZUY
HR5ydsVhiglNjIdlCns8v8bryrvSfk991PI8+TIea2YDzZUFWCeRJnEjSNk0434M
O/s6wopBrcOrm0jrobt91re/A8cR8hurc5dElenJqObXGsJdfZTCDf8yZmMkhxkB
PkTh/FwcSNi5o2/lbA0dx6dQ49B8K0Y0vD+YfNoBcwFYjcgqrLkZmPB8LjbacL64
6kHGtX4f5j4lSTTPoboMCDoAPxYswB7B9VIyYMyJS7/ehNM75k6BDYYcsHp2r3r8
ygwDtPC7XCg3jfLcZKHulysXoNWZHaejjmpNzmyUZgJVYcz2oBccJWac+MPnhtCn
ykCF0IBCLSYIydhSHO7YLfx6XR+HCciifRljqTTL4yp70VaC9aemknfGVdxls1QH
NGe05aDxZJGeek+RUPWkyxWr0AEjV22yhmOGVih4lVi/PN2zyXIn3o7Y2hhwHMJf
IWiiYk24MwxJEBxPQxLn1KRJA8qSofRh6js72SP3piHO7kC3fE5PTO3/b74DeD1p
YO6btwienBzzkSb9rXFjIuZSuAlsdY+y1rEoxn+aNAoiCO7mgbQmXxrgXeZo2uHN
609yLiyOpRjmMBWesVJKfxW2tX1FdX2/rBqVECZE+J7KCIQty5Ru9rJ6UEhfSQvL
sJn4dvsYQgbOZ0XpB+zUK8YVKOpkEIRb3f2XUFdW0hHgNuACqq5Ff9H6XkeqkhKN
axN4UpViZVUn417Rp+0L7TuxXo1DYuz8CgbAAaDLmHD3iGw3LHlX3cms0ByG6NBk
ma53LmnfAopzyuip0ww/wj7NXSMSL2yp03LeHJ5RWlnrVDuF2cdg8CWgxMMmbYW5
y/7G81n7tOBHdxW7OGTzQ8yFBaA9nmQH7TWbOO656zSyf1l98+DLxiK349jU1okL
73rbHebIfTiHCiWhF74QKbRWkSCkE7YAsei3h8xUsrlNu0CRJ9O6ulRyCT8ohHzy
/22y7a2zDoSqG5KDEGW10rXqCYtkvR8kxnWBFIXNCL9JE5UXWd+11FlBnqEvbKtM
OG3+wN3ZyTgyRr6yurDIqVn2TGx/3jQXCyUZMqDe2RZkZj5H7TZImsIe/jqy9zlo
8E+vUB78VM/j6og5ZAkxP1dQ0rOwhXUIm4vlq2hKD8Dc/cqtom2qxH7DZKQ10/Iz
Tc4L17+iz/lkVCOIMccU02EAOXHAi6Nx0zW5UJRIfFg+mLFoEkfrSgMEbi+Wg5qc
SHf0oePPmH211BxwQuIpSm2H56g8Z8pb1Tvp3zDrAHShk1EYNEJKFbBkGKOpAo9H
EV8/ZztMKCHuWaOtQ5MLdleEZrAfb6vyPNZK4aAZGa9b6KGGH1LvwYJgZ9Ht7Uy9
XDxW0sOI5BCvwEiklZ+s4QkR+7o2g5IIS39MQU9xYVqCGoNu3qL/8uO/xFpf1NP6
+7WD/S2CMMNwsVrwuPnYzhuRNtrxeNVTs3d6+rmx9VMjz1D1VJ1zmsFI5D0VzAP6
EzeS3lV0DRuMfFGz95kpioqCgOlHeiwklantSEAKEWkO1AenRhtAPDBKGhuVHVCv
6hiE6qeH2JcF4xvD0erquF+PIlbHOotHAtKi65D9mtC8fMO3uvPawbDTWYWejsYg
6llFbfZSvyjRX2o2vpxT2ZjMV887TEX2r9Gy7Ik7U4eCuHuOZL1/Qjl5j/4E6W+d
g0r9Dvy5D1ScCgbJXwobzF9i2qfjTuSez+kg1qyNRhQqp89MWvXrrEAuAX1HM0K+
nlFHTeoY/UkcGHK8dFSXVHp9MZQufsb+e0EgjD9SYtG3oRKmGJmWbGHFc5h71SV6
XND4VjM25Ejp7S4IP/OvYqeJUa+Ljnh07pUZfbgK8mc+2BYxT7qdEUbzzlY8G/HK
wdte9NApi++u7xduPDfH+cLml21T+h32LRLs8w28Qu+D1VhII4MSnrY0lcFD8fuh
FqieJhfajRgVkc/hxjfo8ULmyz+uUgKIV3rRV8FRISivgLbbVPy1dYDmYJiP+Aeb
wGegkiE6o77ijR8BWdAxU+T7qnXNNCrjs3X/Q5+108hok0Hd4amTDDBJQmFD782N
uMp+6Uhb+d8BmLFm1wncIEbWB5NuMCooRwa+3VtG2IR6i8ekOspw9AOS98Jg8sC4
zyjd9507JHZB6KAOSCv6g8yVXTEgTRWK2RzXROaTUXVv3Gj4lr4aN3YBzYgAf741
VuWY0F4qr3RvgPlr15V/WouQDEOmi1Cb/ye1nMgPZpTveErOkitwOF5ctupu7pdd
UEv0UacUL7RP4mHx9UJlNrrkZQ7VLD4qB9VJelyeayCH+kLn4+Q4HBVREm6VkVFB
h4mlMb2DC+TgOtRgDYz4g1TDk2OrFLZ4fNqqc2hYxvkyFFfrgkDCU7i6lfNlFoGU
RNk68kL9wO7LkzYrkKvmugldWtz0yKl6vkhEjC26ZmwgZbT24pYVk+YuUlIt/9Af
EauGXD/rxvAsMRp32wdlnXJfD6Y/yJspBYz+81PvX0VEqGM0lwEKlg+lK2Vik7Di
PhVBOqBHRZSYhqeZz0RPxfd9GulG/zf/QlOFRFS1V5BySW3X6z6eFP82kDa50JjZ
FIbnj7ocTZvKmBxF2dv7iFevNEcWi/uEdewZZ7CTVj7bncMrY0bzk3nrScEpxHt+
+2ZRd2zUQde72zpe17vXHnKvGTozJwhTZG3oqin8liE4CrqXyAHau0i3st5pPeld
5k92faVW6XjU2OwnoX9pCBb093nIHxXvKbP4v10g9w/edqetnpiRujaiq4Wj7IbE
zxmD0JCCTdg4WZslI5s+jBdpaRNUmiEOVkHAeQPjdk258H3ikh4EDK7GL8o9d+Kw
ckfMIxnrPfVn+FlaVfCbnKgP/lDFd9lItHQ99nmSyw89m2aJ1vqBAg7lAAesmWnn
nnsX5JW+OuzWKdg8SmHI2E3LFwAQInUATN2T0svtsA5DKTzZAFqaynG05qmfSv+v
RbxyzkKUstJZUFZfsGPN3HXZX2RT+H05bCqTvIl7g6vjX6G3RdYtL1cZXV2s5JH2
WwoVJnuT/Z7Ez9j19PgPd4sUePEcw8I8ZeOIa/tberyiYs6LEY1s2pFptioiQJbk
Hjq++d3XJnAzVLJOYXnYV5KC8LIamc+KlhqDsdLs3tk2rKixC+0TEypW78UlkG/m
9pS8ezS5orU0GNNThps67aMOcCCWyraA8emWP85lopk7h73lrYu4D+IneUvVnbGa
k/99Lxf3PoL4qtW2SfP4f64GTVIMuWDxEQ9zeWlst2FzJSSkLD8gi4j7WOd0q5A0
27MTn/gVzVHqJ6j3Z/JcXbmeXv5YpTBeYT9v16B9p3jc72NHJrKyST8wR25t/5j8
LjwADJHRTgz0jq2srdh5v8Mm+mI0fUAJrrYUebRRR8VRWGxLCcvUTNQEe4mCD4MF
zXzrytgltpAsNN35l8s/M5y7cTqQac7/73wFiQ7tJkqwVMBSj/BZ9KozAUShsmD7
eT0FJcveqoiGRdqDCI+NZ7qRvORjsjmNq/uBzD/mQW7YJvXumzJDqGmWpz0s+DyZ
niSqif3Udvyc4dqwqI2VDfq27ALXbSgppsTIep6j8x9/qX9RTgQaEx64FL0pK7Fo
0XHaZZLFGWRqV1MbyfjAvFX64e0tVS+CrWTS9/2eGzPISZt/zFob22hxt8qle+Xp
TSYC+9PFqSKLC4WibUsYrAsPtHarsDjEgPcHrbLys3s3u/mpd99Yg5Ye1LgVvdHq
xsmr69lVcGQpp9eGosBN/f3A1o/Q4Kvl2SKr+pLK1T/JQo0RQnpS9taWSRnI2YmG
k4rWkUZWJaX0k/I+b/7riSU4C87jY8QCywQK4cbvgNgWxp0L4s29y2amFPjQrAqP
zJZ2rg6l5hZ0fMU86DYEwznwL73u8epZSAAAaE3TNx4hHKmLfQF8L/SJyjIIwP92
r57Aup9i6F5l5y990g+vyzT3bO+cB1w5Xu4IjYYPluLi+9O7P2p93IKxEF0eKIz+
ILEWx5UdB38TbjaZmknQO/XgDGTOmqU65/ZP4MiLXR+qsXTMQdOc0tRB84UvfCSc
zIWbj9RdiDAJmZwHR01kzqN/6N7P1Y0l+k0IxGs3RD+3DYtycKDE7QYa2uqGnMj5
89nPcEUCaYE7Bj/si/ajd3GJUM2sXHXWXcqLEZb4TG0ZpnaFruoVG83qDrJO/lso
UTa4ZJWUUOKqjI/kNWiPmJdDVYMDUWrOxD0cFHQXHlevRtpRZe6lD6Jf9/vK29g9
5a7eDvy8IG4fO6KsdKA8D3aJ00qdO/8FckfMjbdQWvv7WAquM001hzWaQNP9fNyg
XSwl3uBp+VZdH7ALx97Pe3ReeegQCngNmWo3lVjhby9H+eibfiWPOhngWbfGr9Dl
M0VnZffYRpfU8RnGZoOSwHTG6pt98a2LFJmQzdJZnN2gjKm58PoKPL3ypDMPD9eP
2QY9FuRCEB5K4MDBch/k9GY123rzNk9RUCSzNXrdebCMzEqvpZDssMVR98LoMyjw
v1H40DTsVAuYXZyi7b0CzHLYgLGBG97zyaC/v80or4pVr/RqjtopBNeY403clZ9f
RtfDhpHCVPBYZnnBl699rDFe6Ph/8R8KOmUHowQuIc44VihvG46Lnyurw3Wdqjsh
u18ZUZYsj0nq2GwYCzTjf+vvIUumDKXWoqoAPDhkxkAWZed7pAb30ynFmWX2GSm9
efhI2iOPIzu0e5WdG8FLz+92QrySMCUCsNSuxzWZ4/1YdNRon4jt708bVqglajDK
pZ/pTGC+pDTt1TDUcOge9EgC0JfJc03kB2vrhAfBnYWOf+Kq/Vz9Gi/1Kzhi+UwT
BZpzWCcgzxtKIsdOuHKWQ3QkpSiCc5rNZzjJJ3W8bOdobX3ObpDQdNSAw1SWbeQK
OESDks9R84bsUlHeYFmuU1FYe3oV7dqdc6MEGCnpQHey6O9IHGmiXDIrjtqMqNTx
oSrZTCiuuaMHMzRMYieAmJkSOgpz/u8kIyQridH0lbl/zn7+6kPEopOmMcy86Sqn
YzDmAtAAPQYSf3eBoSiyzTm5E0nfF0zi8sJ+7QbCpAjE0kAAV4nxrw0G69526k/i
ZiBzhzeTtPl2YebU19tHMRUFGkLK5BfsJpRxQhu63jLLUociVd8VR6LQdt2XFvv3
PftAS99ruDiyG623LbO/wzzJCz2kjJ+XL+Hbhwiq7SBFKp1SGXXOfgYhWcPnA2GK
gBMqXoqUQi/+uaE2dq4MOtJrfR7ndbqsEkkoMz9rw0Q/AUGKGy0buqivqt2czude
C5OOFP3/57O0Tt0DCIqpzG9IzHKzJ8Pozh1J66l7b15oLY6RoIdTDhJ1fwsAjkCf
zKYBsO3ju0pSZMpkwOoMFb4d8DUZSs45OdeXWTbKRxvWUtLqvShKk0oWE6zr3SOw
8TaV253pdKNR6ChKGk8rwTvnABi3aOsJcNIYVw9gJ+72HT5iR3D3IhGBjueobTc2
5JGEl5T3VevL5VlqB/gzgM3CQRvcxF2kBH4CPAAq/xQOji5s24g6YZmri6XS/4Lw
aUmyeHHPesvRnKf1PIqd5C/z9LjQgCDA6ec866r7ytWIF/MqSVFkbqHrGR/JG3SQ
PIdPXMZEiwbwzulBDr4/HiEZjYX+xrwmESA1N/S7rjy8yLGuRmfvyVdoZa1NoH6O
lk8E58HZOe4K6bl3e9fUqVRTvjv4G9GcvaInDhH/DyFqGiSZ6LNi4psI7Ya6QzI5
WyvT70LzL1z9qv6P3l91/zebuF1dj7a/TpnxmQo8MnEdivMklX0H0lulG76oMXoj
jrUg41iJH6XbUi7myE0FupVqO99qvLWLH84GfXb9/PjUEyO4c+695Kq093Fxwis0
g7CmtT6M50UgXHwvsnnwMYp6PfMEieOC2DIHvf+66WSJlyIEkoOJobdMoOGD4mAy
O/2+UafMXvEdnRXH3PQV1BU+RT4HZTNx1mecSUXW17JqFm7IuFuZqrUiIewj4KFX
vTCXExva1TIAie4yaW5VGttihUhiwwgQfp0mzqRSG8NMQJaqzMOndDUxqcAZ2sNx
XtE47XQ6hOrAxdNER01t6NRXHeiV/su9290UkBMFZO6Ds9TNes6qxrHqa5Ct1OE/
8dgUSr07jIKoneAUU/d0IFa+WdOXPTqsKZZSrOuR8x7TCXs0KfFgvWyDUPcW3kbO
ePHOAimStSFDYo3X+nr0jySxUzukdxdlDPicG35O8yyeFgKNL+ZJUQqAacnju11/
yb7qzyFRJR44AI/Cdi3LSONLYAlysvLpyIRLxTnz/CH3+I2PLGxbTein3LxKIATz
jqjV3rDMet6BaFr67LuMsloOgsGdKvi5O26/pR4lf+e+uqnrGjXew1wbrz+n9Nk8
abEeNM1TyMFLYMewTssw6Se318s6UbP2xrvoSWQEsTr63fhV2OswHz6nDaaGyN8f
g7oZ4T3Rw1CFOGfS4y1UFV12pzACXFm57guFWtWLW0F74RbEOrv+2pONPtu7Strn
B0uwDu8YOm4PxFk8MSD0ME23ntQzfnaJpJRj6OFJMme/JjJdgZyhS6lh6YlDlVFr
QwTDPoseIteWrR7PBz922cR6D38xw2UXH727upueB5FNl1bbHJip8i6FoeKjfrxj
gwHgovpFvzR2KdimlwoVTrFW09kNXJOkHFzEyRqAFZWUJiWmyvwNdP6wLGXPaVxt
qZfh2N3VDRtE2kbJzBlW0Uv5FBYXrRe0lZ8gy21HqB40r69y/z9VP74NEtJH9huo
JZKS+2rFckxBIesPtlGeqISUp8PUDemjLVNXr+K8U9PvOhH30vfcuwIN1hjwwmCq
gE7M5u615HfeHCQtFI58S++m52IXobSXPS8ZwVf8t5Qr3rmmpt1sTw5onWlRwpOw
Us4A67P9ScEDsiJggoKBtazjlvvqP8Zh1BLgHgA/Ofk6pewAN+AzlMqQtdGP8g1A
NOchLddc2Kn84uBr8zE+FseobH5+XCL9dZwA15Pbf9VMj/65dwt5j5xh4FG29eUT
LZGMg1fwcxGcQxE7u6dYm8z9udlB+WSNSR0+Qe9ctVmDEWDFhkB7rvsrZhj65ZHZ
hzM/HhjG+6C+DCwKaaJ8u76TsIzOAQsyZ/YO4b0JkV5TBR4mv7h8EZgh7hBMmbZW
8eoYHy12RiTS3hEkl9JJag32w/nLK34DS759GzzxakA=
`pragma protect end_protected
