// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:35:01 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NxxhXzBBSsmBMOYg/Y89aDJQfCUxR+ocISVEttl4Jq4pNLYAywt1e0oyP+jNJFiy
4pmUhbqaP44bd2tGOsut6WYJKIRmFy2OMdKdEFHw/KcPskG7RmX8klnN9o1QDNvT
SagE7A1tzGk7B1Ic784meApoRuwPlZWAl1YEpwUIl7g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12560)
fENpSaXVHfhuoHZdU7Ith77ve8iHheK857RHuTSx2IVqrMYaO7VxpmsiM6NJKj6b
xbFA25Vm1GX2VlS1S1yK6E8cY57HPPuGJuUENHosyMVMNjTxs6mTxpKQ5zcY6W18
LgxRH1a6OvGVeeQuJtk9jzc6Pr4Rmwvio91HWGisAUY7YCxE3POlTtBW048hJFVz
vNJY/WEHbd3XOAUHCR1kT3m0/ssdNYCouJQKrSZD9rzZxKEAZ9WQWR33Qn45UcGM
rv1n9rEjEMEkoi77khqazOLodrIV4nEMXPdE4yJVBVHE7W/lgk8JJw5oTZERNimG
bahCplJK2e+l8HFvjAXZ0Dwn68HE90yyjMl/CBHmnLlGUDK6EoRqkzEY/d2YX27s
XPwiVPM9uqEPrZpGR2T8irLqqAfdXu4pl2i5fU5kd5WO42DtVwYEy3+x1QmnUlwB
SWBJGiT7c3n+ZGK0TgheitQE4XxcN9oiEAAVpM3L3wI1D42sfaoKnt60uOa41k5A
v3uhaqwTEIYVJgtWXtmwQVOueapcVMEvwo4JnO5BwzHCuvoZCO8JfbHUFiVX4lyT
RtH/4N2Uwzb4LFDW1Z1/RAp0NPfY6M++OseYzXmeA5QV1wL3ENnaxnodLJpkS71P
E2I30dK3zaGGi9DbX9WS9ji9NcJRfsXzDvWKv3fc5wchqf8ZQVE6AIilDjT9kR8v
s+rQKBvO9kJ8McV4mlcmVFajYh2C/G2rxRxsDbqVQ1FYMsxhLoWhp+91uAJgz7mr
smDcoVlirO/7fr3DAIW2r4lSdM9nqw3V8IWM5KNQNAORu6t11gQMmd/KN0P9kaMF
KFezRZdvZcXhMZrIdokjclF2XcelGEpCbLclpZMoZ15NQ6n0yx87M6GFkmoPfDlz
ujCb3KlCClsTEi6h8kGlyFAHGMms+IsEA4V5jVfsFR8ug+8TyCD2OuMFMWKA+BNk
RZvwIRa1jkHRHYJKkLRv5hdYcn94jcoJhL55gLHAn+fnp+lSpubFwLIMvae/XzCv
92RLqlP5rCuxMlyLdS8xsPJNdu4fgbKADBIM5pgbmHJKy11rsXjnHOpLXrJvIw/R
f5iwxXuKEGTuwONFDYsrAcWCdLxJUf3sxaf66T1K+LDwtQutY5AALduxS19fq+mn
QikezY2lGVYCShvClFNDA92MAQgjvxzUveoHYsesA654BqgaIou6Pe4bvguCqVFv
o0NSoyW81fE5S3p1DgkJKSxvUr2IaiwzzDBHncFBSl5v2GGEv0/uwLr0lv9zNA1Z
5GmIP/RJI6D/fRbcftBbbW7UDNRmrkUOQPzBkrRndUgIbYp0DQFfaLgokKg2+GcL
rU6DFUMEvWsyyB9aRm8vyeI7U7+/2kIbHNhLaY6RCIBGUk/H6g9+mpPViIW6sz3s
vrRz9HjZdc1ypBKRwyylX3Nng8BCHb6MUWqNf16nuk6ZfXYCzCCJykA+6LS2+tkw
FAJjd7schYr+MX+z+PClL3Ovbul6IW92AfUuNPwS6kSyjdpgKa77qSB4/SbPNbbn
W1G43/aioRVcQwDhN2cgYHS1FUlcr19NLUA+xBIv9KG0yvj0WWJsaZXmOTcejpmM
Gc0zWUYW1sbMspep3Q1JXdTXKdx4ZsHEcYph6y8g7Vt5ETlhmgRn2YErVzyIW7fe
7/Kb0gmKAtmZCmOrLJsyd5y0Fce0knG0CoBCxFev5OjF/GTBv3jNQJJIUpkA4Bzc
YL/aMRTupJXTwaLMj2aZkCUU+P2+TWcNaYQgvRxMubPViBHTWib2g5E/xsHCox0v
QuNrpJB15vpsQ0i73yEIpJ++RaxxywhXNAnOE9f8QOVguGd8b7XtE6VAWVexbx8O
S0+lS4KLLt3mIvxN+GS98NWhBykBVSM+OwH2gvh1zveSz+Oio7XZZNg8jDjq+k1g
MRV9skO3/ECOTd4o0bigKQtxNxPynvuWzuSL7aFzNx7H/CshqOWr04uarYHwjs3L
+oAA6nde4lNlEOgah3TUsFgm4r+2804JJJkYMrPIS9BN7+qJjrw5Q0YS+Ca7H/Ey
7S/9EtJXOwYtmVhEaaN2ZKqtXYRoSzGrH7cZbbp8Rj74/JHEYihfTENQtysh26bl
AsVl9FOM73dBXR/g+R2oDdHkt5+eQh5Vwd6C4I5eLFcmLAJZRh4OoxSwLFVRKRtp
jRfRQRH93dvn29gx1kaTERfCHoGwoRdWOL4YKT/IG5JbGOuzl+v89LjC7io9u5tf
w8PZhB9l0Dap8+TLYzzsExMGK6S35Z8m9ULS3alkMeMRbKlrcn0VaIGmyO6lpdQ/
C+c2LSuPNWrCadjNcKWQhu4vC9UGkEVuBR5FFAeh4/xppQYCh5bFxkW3hwiTt5ec
WFnec+sc9Sa2z/VugY57qoWfA7/AdiGDlz3WJP25n9iVLaweN0ZbmNvCti565WEc
mQmPTBW2jt/APg+ftAvU4snHI9PWRIr+PLKKl71YScfI+kLCZfKKfgndfBtpJfrq
pKOOkoHseOGpeRmGYUD2Wc6LG9xNMndk5AnIFGTBnGOLsltXqQ88ZWTNRibnDoxU
elvCIoeYAfiE7mnWLeZ8oP7Dd1giI++2a/q69X8O6l5LMrFcPx1c3hgtQHJxagLC
+i9oVo6VoKeUg8UwpyhiIk0ItqWhAvRZ+SPFtUHNW39BYSWFU8hj8u0DWqtrT7uy
NyQ6KG2EYjDBqSvlOkIaI/4l1xPWgDUeBGMVaoADqgMbkF6qPcbAINLhCUM8P6LF
eAzp+qJ8W++hJm3sZ/15MgAAvONjFpqOiKpWZchHY8D4jbLfGpkF2gdThpZHwLG2
kwXYRYQv3qXve/jdVLsaWIoM23L8uMYyoSMDhE9gmZ3uQmWBvShBWbviO5aPQDkF
4j7U6Js6ARW/nrJcVbIwdRh8espPKZFUHhja0j7TIfUg9nTnBYUpvHlFoVWxDbHf
HxUbEq7A4zp6XQTdc1RwdJnp6fYuJhMdtnBWPeFe6b7nrb5alZ3u9k3D43QgBwxc
dAZyte0I0xulwbL8neDdX8JX6P5rqkFNy+uSRr6RAzj5n2N8UwVHtyd5hKj/Ujlp
GiVgy3OhZ7zNmnSchBKe5CI7HxIXiy5k+PUsGTYblcvEzE5rCF1+OMkGj62oQnWz
7Yr+icaN8G1TsUOAkNJWvZNt3ySQnCKe2QIVybC15rA/mJ2iLAeU5ILyu+uREbAP
0ZI3e8bYFrYMR6cA0xIATBAoOcDw6STgu3s41LgRUmZ9vrFQ5qh4VM+nRgjhk6cB
Nj8G08r2CDcjWIKnQJbUCM3UOiu7ktUsk/BKgyWFzSDfX7PiSyb52iKGNff8xFIY
f9U8qDd1F5iCNNVSM0E3YTma2yvBueBLXsv2ihrj7leHQtjEKXOy9c7QXnbtKcEX
yzboGvAOlrOnirGMQW6ymvWpqF6Xa0tW6tSGZR4rqmsn7fs1h+j0bJ6i66R952BM
upRbgiAM+SFneJ+D1H9kuibPPsHn3QVc5JIYHDJneBWBVLzseGqms6MoBcpevqc0
7GZ/dPzBse2qmcLLYkM2SkrujkcjldZuhHKRtvbkpX6IT8uaCzIJpnz3KxXEhyGI
64wqGmi6u+9VVcZ+GR4QBKjZE62JfFF2iav/FINkCSIZxR4elt0pdW1HL3XQlW/V
prUUUqZb+YTIIwScvJcLubIoeq24ij4hKuKu6n/1U3strEmSuRl8+dpN5UDpRfEA
EhL4LeNcFoRFKdqBIfIF+FOctZ66W1pWYg5yBQVKISpqJMxP5+MSXzauSyZ62AyG
rEvu9wf9usTSvhzAMKTrg1hMv5879AGqHC1DhetTj5NzmBRNCM+obODkfDVftk5a
LgoTLhln48MKbe+W/7D/PovUILvZUu5ReGIB6tuWGhNeeHnbCQgCvZphesHt56m1
W7YPI2Q5M+4a6vJQeaE0MxFWV3FzCCLaJg8sQjXA092jRCuK2Fq8IJndHQuar7hb
J9Yx9HpObdKVg+KSVeWhPjXA3jtDZj+a31wRvy7w+EnYWZkWdNj8n4bXUr5PwkFE
9bB5iEaIy85JrlrxBGESI3kiOo0uVYi1leJ0wjCxMz+pscIy6Ro2Ee7ARqGzdkGo
wnlMFxVXbFeaENSLA1KhsGzjezwDn3+pNn6wDUvpa6Ne92MiGwniCMbSbfzr1XtS
VSKQG332FB/kDYCSPjjwmWv4esrNg95E3nZEd0V/usQiZ8li19vscAxnEuyteEVz
nS9ccsFLUvLNhUcYilbkKA1lrB3UcjEwY7oeeu9+PN35A89jBD5IbWmHc2d+Yz/C
4X5oFyU1y2ePzxR6gS1i/4Kz1ELUAtkMmtsg+FVbrSEAv7lxV/OdCWzPT2iE9kva
JyR7lqvON0dDWHUcHyx7LiJ7a1kJ4CsXcoY8nhncW7VI5zbee3D4KUSZpHiQze68
hqBfvBfZ3TrDI7+M+cOkT/yhBtKirDDJLn/2QsQo5Iidq09cqTq0srwpb0Mh8ira
O88kneZdLye3QKw1xWCOVUv7aoGGItU00phCfmstFitV72NjEWV5f3hsX5YWDJOi
6Fz6cJcSWP09eJ6X8gXC6TbrycX06bIFQ13AYstYp3XEc6Zzh7WJRqHHb7KqJejT
/k64FZmmh2NiaFZRYKnLPcHe40WLv1ks1ztcGfZ3JFkGk7BMTlvt0R1rbb2lZceQ
na1N003yfyCX3zfHISsJDHlEcszLk9PSFRYilrDgsaJYyt5soCOn2CDAqFxGYFlU
gsYzujT/JbqvhtigS0+n6KR981wm5Uh37lSSf5UwssUCZzQ8gJwbIfcYbVtuAQ1o
WSP3QrGI5gu5xlilw8QKIr1Izh/pK70KHyoA/W7SLz6zF4zkHlyZ/PpgIcjT+DXp
7X+o7Kt/ox4rGGBT0zd4Sobe23zegpeqguWtVZQJRGUKevW9Sq2Y4zoYf2Z8pfvp
ndxZZuPfthvq0ZgWRMZgUPitXH9TcGoLNDxOy6Jmvc8j0j74q0NntQ9Bsn5dgCsG
JzTkkcUudmhwMLtwG1iOgwNvDaar8RTwOZhU8hr8Dgt/LUh1w6+M/D8KE1qrZvbf
lYB43WP2y3rym0nHBWHeuYYxGkqogXF6rtKDnMazQwhY3PhI71OONX4V50EXw2Ti
iszln3JgMZMgohzSkQwEf6JPVudmnOqG2lUyNLEN8G36aBEgk2C0zr9cC3trMtQ4
2lxCTk2HbYW/oucmm17bd7l2BAVJEy10xpocCdnVJ8uSQd09HMOaF2yyJUHrtvqn
NfvD6uAJsCBIraat79c+pYGHxDgA5k0z+dpQAoiMl3MNJ0N8WGMQxjXYH4kpoNy0
OHpgNFu0zvfkrBebfeRAMRhe5/LnKAz1zJERD6L5UBe86rxbFYzROoiEG89YWT+Z
672BQpIcDT6XGK6OimoI4fVOX2RIm+mZsUPxuJX5/AaZmY2lDipXdsYVDyizogF2
7M38e1DvZGxk/rxndPvkfyJDU/ifhsRHyik+UNjv+c8/lpeVppm3aLDjz/wXqKA7
LnQhbgXq3VbLOroaT50oleOokTUAAsxwoz3QmZxRCPVbqOF1gWDc9jaIJpA8P/4D
rUmdfz+ZpctBYOi9CZoLk7gJm6P+32mV8Ed/ioyiZG6eEn6Z49J9Og/db3xGROT3
ooRa1iiBuQE2MOAVQW6+SRSv4zT5nnagYMfOFU/gE2ewpTEr5//LlUMMoClyNOIe
qBO60z/fHdS7fBN7GomyWrf+gIecOZh1pP+5FVfvGFF/6x3bf7tNLytQAiwVMRFg
bcXmgsgUEZxEjaxnXEoxUE7KCHw5SjOJWNheCWx7FdcrZrqZigV9kKtUM1S9RsW8
/CRc6H54AJEmiehE4U1X+NG23p/u1JB7AC64jsXMrc+Av0H3RyFrcN0vdsRDsgWa
hQaWFiIDqWKAdN/483MxrOoDrNN5L5G/hP7fnFavJPMYNfMkJpcljQl2chDJ7Ess
l70jjEz1YfuXnSd8b0orYdY/u9KkUvfGkOo2UH32hZReuakYiSIyV9kUYod34Mx1
2O1T7GWUzKo2IJ8sEq4vNgPXTIvW/gE/6EyfVG6vho1shrJXusLX1WGWUYlxElaf
/Ld4E0otJrcTF5VYHyUAXb7Z/2es5ZnVT1rP+4uaavG6z2nxbbPAz3f4wZvPYBbs
1x6Vcxy20GKy7/S6/TjI/SClW+bcBY2pEaxMat2ytMx4aLlW7DB7xguLpaDfU706
yPHNbZLz++fb4YUI+dSB3hYo/KAC6RtfolWtM7pnHvvCy8BXyPCvUzQu6QWTan2l
ZHj4fLIkDrVNQy7VDird7GGOhmtIrnIqq83kctxxHB04QYfVdZVuKIQMRKOWBIM3
A80XA3yRGU3zfuwLiZePA/2Nth3Whn25p8SisdFYTpixH5yar9kF7pdoxkAxDI8W
jtjRducMa245Hmk2Kfq80vwEOA3qeVL49uRj5oYNrBGch2/dtXcqXRqcK/mQaotz
XDB2cDHzL8q/yZM8EQoXpLU8gsWNrspLvfWzntG8tLAxFuEdZet7/SqHYuGbdzY9
MRBPOVtamZW/SpiQqoPEIxJGvsNn822LVcgQD3DOW5K7hgeraT5TY7/WRcPTOH8e
BFnlhX/t3yyElxqAqaW6MTxmw6C8pL3R61Pm/nVGG6Fjfc6YwJMiv1VKCVRwO2hm
mmukwsZAkb1xs8cLFr0351CipOxE7kckQFs6NqcDf5IaLF/DYRilsshLBMaN/atZ
z6wPSPg5DuVaj+ApwfqoArmQN1cKTRznqJwIcSL3LaDbPtq4S9zb+l1Lkyh2Zrxa
nDD8h6TFK/BQ5hQk0NsWThjggeoDf0D95w+JlfKytteOMC6aB8pgiHDhILccI3BB
GyL7qZlMvQlJblM/+ntUifMDxj1PJ3fNo0zuarJTG4yD42j+QPmO2uJ+PPLaVdOz
KHjA+jjO4x/YbDiI0RWHKfZD+dfc0vJQdO825kd7ON85Nxymv7jwpXYchychlxcw
7iPzAX7kuh5EPfX6B7Ku5IKJuDuGY0/4G3LKzVY5g4kmg5W27tzAheSDH4BeVAEa
c6VS7lcql5f+jS7nNMAXHgbcnVkqirbe47nkl7MIjXAnhjipZZkAowOJgFMNAxTa
C55hGyJzfhw1ne59g/NPQhGASZQwCnO8iY6UV7jFjXGoUWNNTDMsMgTsQmMcX99S
t6p2reK7Li3avz4iqGSwX5ODMKx1GYLFeUpDqV3ZcnaX00G+3vl7+A+2VzaNPdMM
tU2UmcNQivZ8h6uvjO+5/CD3JMpkVqNzVU2uuaXb5QJkI7R84mEcOfLCxahWNztE
JHAK10g1gLRc1lzoDk1vXa0tTkqwDRipyXrJJ3aUEkmiBGoBGcwXLkdkpPpBqhe7
lgWfkK6h18FcDPiyUSeboOHRDVaK3MFLPDinOrQnbkXOtqPhqgaB0MB+VwSxAaOd
aDonoPdwqlwxJIXrSMrwph6Jv7BMyT7YhgjKnAXPD/6mFGkcpG5Sx4XwNG0icxx/
pZRs57fuDoOTNqu+rYiF5gu7CvB5Z2cVQ3+8cpbNOQA83Xqqes+gY6Cs3totH1gL
Ixj+avsWtcqyCDezYVIbbkZUfks92z7Y6dwOZQ/L6lSJXANBJKP8VgG+V3ucW4iU
wwTiqpP+2FLBWXP87CCw1pUdvypD5Sr9hXeREGAzcsP9Fy7dKvrlkHZim5/zEm8Z
iXHVkSeS73FA6OpNUltJh//05WRmUvdOwW+dFmtdUCkgDS5eR6VnArkq4TVPUCe+
HtxKPuZghiX6L7u3nWzbGD5ynjjOdnfQltwi9089FhBKNX1z8cTrd0Zrz6/MqCoI
MejEWq4HBddXs6g5rFMZxJNfy0OYbn7h2P3xfwQl93mwiT9O/Tv9/EYCyZu1LV7o
VZBCcTrtNcWDFX59hlj298sHb/0iMeMwFx9emldTuHBcw37F/VkT+LblxXTr6fLI
I4sTwHnnv7tdQrjAYspb7qeTr4+IfXbLWgF8w7sPs+O4KT+QRmfsGumZi8HMnQ10
sMypK2AMBDXObHATzc9Ce9BTYS0CvVxcsVGRk6/wLFw7STRKI8c0QKk55nt1yYDW
ZJ4h6T6tey09x+UUwptyfdvLyau68NDLHpsWlam+6Z2RAUBT/8NBSop+hnstv/Sj
LDvDbvyUFfJa8G6qGGdNl99tqZXkY9vPdI84xbfq0z/jT/itbltJ7ZI8foBXVSYO
Ecfw6G2HB2uUPUYOwQYjUug29iBvgGKdOEE2rgqxmx08SGNmnOqCeHyGmE7HDL4P
DFlb/2foWezYmyJtPcL23mjhkzc8TQnZxp+BMzeR8dp7U/ulfJQTym7oHxMhhIYp
DpDLM27R+zTK13iA3bWKlyAIiI9MpsFclZG3aMWqodmS0q7N4xZDW8Yz5CQ/6kqy
eX8Df/HScwCuOga43NnP+YzoJpqICIG0S3ONCf4jPe1BMSHVH2+sIg/mbAYrKvIw
SSkDqDCUh7JIpTBzZRIn44mQZ4JrxVsWQnx/Jod/LWPN6xjlurJYUODhQLeRg3hd
K4fP19ZWXAcHy40uS2wvajWGyS4oAtKBVzWfbeaM24cZJdcXQmfR/d4OO1teiOmW
XN0IdA/bgOqbKezQMvlbMd5xXHWAhqb3XZdT9OQAA2o5PCuUq79sNsukgMtPlXiY
YK5FIRUbY2ZRcA0+4wOTkTgMKujFc0XSQGAa8oeVjKMh334gxy/fzd6kM0n6jXay
xYKV7ALPOEoYc8pXqLWPAB/uE3OyD/WSj3/+gKnYCPVkVdndYLtybLwNwN4l5YMb
NmElrSodnMbQNu2I5S/za6RcXqhOziS2mhd48PSOH+9CBoTwnB5SQdjVmYeQ+IAG
NXCJu/QJT5qymc5viVGvrNjZjx/SyVCrWz8YiFVdVaT4C+uIQOckvw0KeoaJSBFm
qMSZ1Pj2RPj1j2QB910kfcQddxSEGi83IKXdju28z3ferNW7wionz4NcfXUizWK4
lCUTjlXID3h0FTI85uf4JP14aTEJQPKW59nLC1AhCOIJDXWRsHq+H0bx0nELXyB4
2UjA92vxqTApLf0IGGjgOKeNbE6KP6w2Slh678MgfIh11/4mnOd4fEGtXVFHNMUm
WTpfqgRzl5j2Cbsh/6uTrCGNmjj1/23Ko2fSLlFyt61LrvA04iQMZtEp7ViWeeOg
VkDU/wtGsxeRsxTgz3DjQPJz4ZLqOUZAjQ/vOLZ/reRS3vYa5F5AAOwGzwCIl+3r
yAaHr56DPSenQDG9Kxmcds8T/JJgjzavBKgqvHErQG0oRuRw3JgWiTf/MzFu7hW2
ssB3UF/Ozux71Nf4m6KrJuBi/YluRsO89avkMED/p64E8YwpgBFwDMFwmbsn+Fel
3Auj4us6SExiOBg8P3/pjlh+XuiHN5nAJQ/531Z7TcpHXuvdBgvxY2EOf1ylbSeE
HA5TIdXMplNJ2GUcFJRyDYsFnuKvkz71AkuGLz90PPYdReE/TamyMPUYZRmC/XiT
nu8f2WXdewE87FypqDDj/ajCwlXkaUdPew56Au6ngEjYTYFFEf8JT4KnZgoJnDNK
oFnJY35fXsgrYb6t5wgDB/eVtiI6LOcFNn0TThZTrbru1hTE6IC963fEjyRO/7YF
qCdCgP4cI8wU5MHM5X5PRIeilRZ+WBWSUVGMZRup7M8wuU+vafqqvV4Wt/ICuj0Q
X3prHnQr6+6hFr37TYCD9k/RLMQoMbEwnCTP9BTUVKTd7gGCC6OnFruIJvp5ZH2/
WvJ1Zfv+xcKjB1DRrgErSH4bf9BfxegOE+9J4yW8r7cYWXhAyHVys12f/Sj/7INX
Nn7/3IhBSsziDqZUrcpG+yiB4WCDhvLVyluQBnStXQGTR6fatho8jLA2GKkHyHTQ
/DqHAYfcxrOtytY6s+CbxBp2ABnM7ahOQkHqBXt5qlJzwpYoCkO0k/1gLtvER7UV
84qBR7jB3y+95ON9cwzRpgzf1W16uNyozEcugW+QlcZ/wZ3jjvOk1NEM/A/eNlaX
kfx5iPsIa3PRCpeXdgYwUnN00fJeeNmNF+OFXHHLLiJ7s4CgX/AdN4IlLwaAIXUl
GsiM9fFBZD4X8CBDxvPF2ACaUgCvxewTT/ORT67Yjtn32vk0NEyYiGle1mOoAaNi
nVa6VYSpZO09WWXcbRd1gvxFn8uXccrRGVZBovbyjvMvgKKvxcCkV0GHrI4UGuTn
j7SC7CuAywxxhbkv7JXhuImWW+vyqLcnazG26ZEzIsR3gt1xJ8DtKT2pPli3SjmP
bUfBPVx2l1TbUk89rv1dG3MKKHn3QWYvend00lo7zC8u+vHs9IUKSfiu4tOfFFJg
ZN+w0Bt8lcCbihWmrMifHLKRqdLFqkinJRMz2vm2O4ezRjappPXT+Pzkxdb4jYtJ
dTHuXr4M3JI5abN88LrainjKhBv3jfATEweCid5DuswJP3yQ8HlehWVq1IRCfTfh
F4BMRuhoX3sszhNBxN9BiPv3wjtrqkf3ub8UBYz7rzfD+SAHorr4kX07fF4EioNL
9issf04MeiwZ4aNvP0i+meL8A0F5zO2RzvVLq75rF6mgFhJDlo8pVHyj7s3WNBy+
t8z4ACKeNefpeYInjL0GOiRZlWdpXNus8O0Sz83mEZ2RdhaMRE/RSuwPrkNyeReq
ADawE5jWDSp3atw8I0YIYwoxXDA448RKPGTXfk81aza8pgGBaR1ALSE48Sk8v1Dj
2YSCZzMn/Vt6otC+8TmwPrTrKTcAycMQakNJ7phPP/C52XAKOq2pFMKkpywKkEv2
r7IM6R8pmkZK3a8O+OGSOQF1WWPp9WUoFIBy1nqGrpzND8JlUSx6VbwoOJ//Bct1
dShJDjLpn6cF2BigaAX6lgCOjSKYT6eW8ezCQ/1M7U2QvPMEJSK/J4Ok7mjk0cxi
SqFrlNMc/9sPN4u+J1xw4nHY912WdwCJ82Qzd0JKIAZVcw0/lYNWeoqO6h+lLlYh
s5CHRlJni4dDwMNWhms3lIKSFw4fEQ1Vubl1NBFiXt/Z+81Kzr7xc7HnTkaD1YZI
3iaMd0+VolBtopHGKOfF3Mtty7tDzIUxPrQcHizr2L0h+CKMe5J8tlYj20eycrdf
Arb1PQqMNvfOmpZ+eLq09dhGVlvpxTgq5mi0IK/7l7m9CwY8mmDtnnXIox7+YkNp
Dr1RzrQc1JDaV1AK6ga44jhtg0+FZPuG6LmViE0vNu8Vf4uSvSTK7vUAL6Nvm0wX
o7AErXYsxpFDjWuQHSLnH/USB8lP+s+UrFc8n7NiB7Hb5VvKf1rRw0S7ALKW1/E6
JU7Wv88tc3/YQsOqowy4l6/mZgKLOqAM/bxUCNp7l7ijI36W1EqpWQGFw/0PqNpF
cYDi1qdAI4yEvXw3KV0VjYZ9gmMibeR+6l/VpC6iPPnU5O9Q9p4wm/pa0Fodleu8
Ry06iXaA8LKVeuSU2+sR9r3kSZC8fuQjmaPJFaARsxEgTz16AHUCI7gR+fYJW+Dm
3MJaud3RRgTOoywj+3DjaovAnJ+O+DjWkK/PyCZJp5wxYflJL18Sy462qs1ub98a
9n3W2XL/3cxnrwFCUeM6+t7haQtEmwBYpGuuAV/OCvB0Xes4Kqo+38ok7g1lKmzK
hRCI1lGxZkoR4pSXXGqzixIrgLO1PaS++kRj/EmjhAjsCq8jljA4F53a4/Sz5DDE
9J1UZRm8GXemc2t/VLJ6hsjyUsYv3p7kqvsrqPFWbQZIlk0xGrBQtU4fS4ucE6zS
JcWPjaG1tivD+WWnjfBri9O2itEmcw0pB6q/od7Vz756iSVIQdeTrvxV44GQNgP1
sq8Ts8o/pOklB1+fuGmc6kuZY5Sengd8cjXjL4qPqQtuM5ElBxnr02/jyv7MfcT9
C5wajYcKvJaXmpNqQg+yvXKXSvrsbhTRzcpRlAjAkNgq4UU4zlxX3V9DEUN2Bmta
zqEBUl8jNV3+CL+gaxT7OMYDWVvf94hLo9QCMdU5Wx+pFxOqya74gfHvXz3SY5wQ
joOWVK5TEAH/swi0ZPdYBcsin9z4Fitbb22RC7VwMEvPo3gEYnc6YLI2c2N/IDal
hJ8lvNW6NfWBBuJrIqovcrJBI+APKN77M4VphHcPWQGXYGC1WtAZI8OMDiuljoc8
g/GKXpiqk0+HF4hmNMxKkkhCpDFAsKh33QO7wauP4NencLRJjwBCEj94PqjjrojC
0zkJhlZ1zpfXjSuSGpI/06rIVAc5m7AoaPpWTYwPaiJiQxDgkxvMTWdV94iOfk7G
zSMiY2nvRUkYBQXgxfVKJY0nB44dk7a4ZhgRkUBN24ytxW/+JwZOIYkLoEy4bASR
74/doKzbMoou4baxkSzLAQembpc6CuDrae3aMYrYbxRhD5k2E6pr8t5suuqmQGN8
FVozWurNejpm+zFjBhv60m21Ln0f3pjQI6fqnwbUHhyXTDsFU9KIhrM7u6PdXI6n
MDOmCmoirdfU0l/Y9dYWxTBMajLIxhG5f8IYCXQCJdLVzOWUDJEZh1UHeudCEBAD
a+OgY/Go/IabFniu1vwx1zFaTqQPgMPoPqbXlyt1Xr2FhBDPnr3pC9+kBRBPYY5j
hXvsBXV7wbN0kO+9zutsiE2Y4CTnSdwoCPv3u0Ce0qAla2+PO4JFo65KLv53spy5
fSOOz07rZBlAn2jKX5S52RdVWvk1Q9ccBLB5hmTg1oWq2CqjbMLKaxb3QZetjF2d
AQc+/1JJ5nuWSLnSzUSMAhEa7OvqNO/9vJbCtfcxBqqWHM1eWXLbCuDh5xIIMlYc
cttQSzBPG7fHcVqaKwD+dP6XuvXbStQSXgzlC7ITwZWuiS0A/1qQM8NuQHbuYxTN
OYxS0wpTUUsl3pOk1ufaL5JY/XMy0JkM6uKTmWgdNFLWKLu1BG8cha7jtzVxAjrc
yEyZCMPoOm6+Yynw7L76UrLvlzFL1LaYPw/vh5p1/sInpYPqq1ohGazRdxDaq392
Mg1ADoiBP3JPHa8Ri7Ikcp7zsMfiHvpbJQqwRJiYZo3sNlZqd4fIdPoQZ9d4aNx8
S8Pt8KSqwiJsL4JI1NdvrnuzJFyODZ6Fy9VXy6dGKaTpT2ktVn2of07vvt8Mheg/
MKXu6NeTh8mUqhMjtrBI8jmdYPkop/LCYH69MFDp4DPY72ielGSya+o8Ds0Upi64
KJzFFNvUvcGRb445lFaWaNnYP1Pye1qyS883Cgw0uSe7FHXDcTAZvqQ5rBXKJq1y
kkg3kIcVRUPryoo6AUs2hfUH9hlrvkAS3WzcQ6LU/eCaOQ6lx4JbqpmT2tI4RJdR
z82k726fRWRwEm5rMo9yo75dyO1AsY41XJYu+FheeRcGd2r/arPEzbrJhlQKWKjH
2dfx90Tua33hLRxagFhnftUtuBt/uAk3Zx37xNvFgt73LsMP/RVtL1p2rbTytVA0
9kAKU7eJji18os2CSguCi5KRVETUc4TNPiw3hY1ccztn7QX2+67vC5M6YVGHivpv
NcZP2WnYPHEV9ozvTKgQ5bNiB1ogGzFT7XDodDz2IcqKl6h4SgKrerEOu42NqdNe
sRNztmSnle7wB6y7pWWaA6MDb+YgUrdkMG+62VfqBfALN5YHcjg1rdsuB/kz1BK2
XAJ05OBYVGGuy8m1bikxwIisYIg2NUrCIhynKU7bsxztQWpHWgw6zjVTNwE/+99+
uLfBzrU/tQ8demAHBMhoOoDUmZoUf0MjJ6dikMgZsri8IIEVxKXW9dOBSqik0NEf
v7PWi84ohjYwjx5ID0Tg3l/97Oh4mq437KJvOFg4I5FvU8DhT99+DshlsNxlDuGh
UkKqekVxnsQAZhx4FIDUFHEYmrWSgEYJguHlCGBh9G1ibvCWDFj7yqGmU4RE2sSn
myQZD1hbaevhc97CeFZvWGow7FZZSDbe8+EUmH15+688wkEAsPEouzFk4as5dzfj
DY1+fUJkk6mgYNGsu7EMRopulLG4GzrHxUG2odpUdxRd1OEMmgyF+WQHWhs02nSH
XyZxMmfXMesL7AvAZM00JZ9gD09+EYm2nPZSHicU/RgO0U3l4TVgP8tEWW8YesAI
+T2/1gzSssKM1U/HdNm1PDTpPFdAswhIA1eN6r1NfkbwdNaPg+YhInB9nqFE9ZGK
cY6QajjP/3NvWxHEFg3s7aLRs1i07LbqxKe9CPp5E0W2gI1v5XckVeHw8JjfcahR
cUl2Y6KGuqcxxcgr8Tnsh1FmsrVLguXdUdKFS096i0j+O0sRiIdhLa1ZyJ8CR16Z
Tlgoku4WvmxVZhsKuPLDF2u3Sp9qVXIETDTJC0xMyomYrEcB46ZO83T87QbtJs6e
QlinQJiOl+RNOLyjui28fOn6XLkLhzOfLnsdkndaWb8iz1v5lG4XTmPdTLC3Pa+3
dUVIi78QvxNA/apP9YSSfsGXWH98qENlUwwsCESMf7ZCKMdAwJaG/cW2BphN74eb
R60S1ig/CuTfxUilUcuEmPuAspY28+3oDZn9IVGR39qD8bgrpyBJc1GcUCmVXVFx
hWAPr9kxGmS5Y/rXhiRb7BV8D4XXnmz1j43idw3cLK22q1IfQjvH0M5FRYHOLVSP
lO+WpGXQKUtcKPJILVattIJnXXRPB7ksQZjGLaFxlB2MkN3IqpnppDPqGtRazuq5
K929ikkEAlufTsfqSEJpOzYVHMhCuwut7/CR2lxIDUWav/yC1fuEC8QWIvbu1pBb
e1uvJ2GQbotISkFDhZW6FGM1sV1x8eS9tUpTO072Rq4yzzlCiFyo6UzygCknNKek
5oqYrmav9OvL2mRpkznC1BE9M9zX0h9qld4K+RNv+j0POvNQQIBV3WbRLz054I9L
MGRRyGixJ4Vqfbwf5p4Y0I0BAQjMAgAX5YSxuxx091zUdxhHckFTNaZVCb0dcGtu
0Tme2OIHd4fFAwdL5mzNSfo9IXj2TRC9ikLNPIX1uRy6zQb09oycsU/gNH6YvlbO
U17JaE6C5XsaB6vjSm8zFb2pu5U0aVvwmWbTHOpehEiVxOgg5cIJSgy1sVc2VHdO
14Kz+iguKK7SPHZ6LylkYD4+AmQanWvAzKVtiI/lVwJ/Vg43ewpeP7jEvQ2Ra+wB
NeTbQ5s99MyhTftd8f8mP7zPK5ljyPyM74cqLgLzDGdzy5njtvI6kTw1Wi62yxuo
7+Tb0f5neVLxxJdIe1crUewJ4QAAGw4A6p3ziQVvaJ/g7liX4Eh8H2ZcJpfd6kUn
pegvVKuYBRGrEiLWqO4jBTSZ4INPhhnECWAeRgqnSWyJiqp+drLLiP5M6nmwaaML
9y28ijCLQfCWIrCsHRuBEo+fFF2KtW3KZrOGbyenVxeB6Qy4Gf7ebbzcj36pLEto
m0+pp+ftM0EoXXNGrCE24aV1KJZmjujWcx/OkMvDPYzkIoExjb96LECncc4UIamC
5jL5EGEIagB8dK6gJk3QKg1t0v42H2+OX8Cvrw5kUBUFwlOxKeAvEfosL0VBExYJ
8UPrw/1PpGdRU/k/pLrWp4VdCCdJ43RwuBEqdlv8eNkj5dy1ODzFNVXitQ4WOWbu
haj03gxxFlkrGhnlr4f4DC4yzo7qlAT31y0u1VvguFXWwlfXIr24QMJ1NsiViw8m
BvQJc6CbqnhX+IiVnBiI8jxNkMV7BnthTkHufVdgB6X4RcKoD6N7ta4siMFXPVPF
7KC1v3UyHeLa9xj92CngJuQDpAkkAEh3mn+ScUHM6Qu4FXtQSOdpXT5ud7u+RmC2
vx5Ay+TTq36zS3yx6hhOVG9UIaoETZzeFllU0wa0l51aW8a2XHHO+y7ze+KVY0PP
2+9HumOpooEVVg5f+TJxO8/dLSBW7dx/9cjQdJ4EXfiTwA1s8KcaIQsvhs8dEDbN
hNFh7ymUQCCRIzv8klILlrSDIKYHBphkeupaObyYXTSGdiUE+tkQAjtCpjVHJ/Bv
tpnfc+gJ3i9eC536zzWF0rj6Mm9p06h0f8A8q74bFznXGNlDiqluMETsU2xJkZU/
6fSXNhOxuCN5dCFIMizKgSXawaWCgfPXitX7rdHPu7M6yv9qFIh3oaom6eJFGIAu
3PgS7HDs7smXQniehpxscWrg44zR+GgHx799VDuaFBg7vlmfsD8NxqX/1XAbjI7Z
r58pS/6AYffT+wKdkAdbs0rotldlnqtHT7W17dEHB1UMW6flwTROINOTxXo6tMvs
R8jeAWq2mdjFnZ2pzoKESjP9TFoo9i+cXPZ5f6xHMioBQHx+lB1o88qw9WzUTA02
Q+G3Eokvs6v/bhkwvirS45LWOwuAcp8mpydul1+8K4bC+qrfUALqEoT8m+I//qxk
61rNsBP9wQfU0Xa6kKf0gFre/lE822PsWVDfoZGRFFKKA0zdE1sqSRBr0v2+3iUM
altbBUgtJ8czGo+aAZsDoMV2Sfl+EmwnZea35o1lBHSLiwieoSqwIQQ7UGgEA64C
/XJzwKpHMwYH5J680zaNQdrPF0ZVDHrpIik4yrcqyOkM5dK85Ju+MFVVIOaYo26O
UeJpRITwdIEqKx3TyRjvkmXWNok52ApCjcMK2UFYf0qKIXrQfxrODrX/NxTed4oL
0ICmwCcFqSotGHQa70kEtANcQ9sYNzS/RNXHhZbTnqgs/QNrQ2TIyQontTMro9hH
p4ASs67WxutJ5TS5/LyBIgwfVmTqrG53i1JqghJPAdPBdslhBgwIQ9ul79DhmU7O
2tLMhMPtcZN15yzBh04w4W1BxeleZKBn5oH30jsUn1CHigvuc08N2tyyBFWhhWP0
QdPsjQf+AIbMzPbr69FzGvoTEvHSkbUGLjPcx7qUrsg=
`pragma protect end_protected
